magic
tech sky130A
magscale 1 2
timestamp 1607837775
<< locali >>
rect 318809 650675 318843 650777
rect 144929 650471 144963 650573
rect 154497 650403 154531 650573
rect 183569 650539 183603 650641
rect 176853 650403 176887 650505
rect 193137 650471 193171 650641
rect 202889 650539 202923 650641
rect 212457 650471 212491 650641
rect 222209 650539 222243 650641
rect 231777 650471 231811 650641
rect 241529 650539 241563 650641
rect 251097 650471 251131 650641
rect 328377 650607 328411 650777
rect 338129 650675 338163 650777
rect 347697 650607 347731 650777
rect 357449 650675 357483 650777
rect 367017 650607 367051 650777
rect 454049 650675 454083 650777
rect 463617 650607 463651 650777
rect 473369 650675 473403 650777
rect 482937 650607 482971 650777
rect 492689 650675 492723 650777
rect 502257 650607 502291 650777
rect 311851 650573 311909 650607
rect 331171 650573 331229 650607
rect 350491 650573 350549 650607
rect 369903 650573 369961 650607
rect 447091 650573 447149 650607
rect 466411 650573 466469 650607
rect 485731 650573 485789 650607
rect 505143 650573 505201 650607
rect 195931 650437 195989 650471
rect 215251 650437 215309 650471
rect 234571 650437 234629 650471
rect 253891 650437 254075 650471
rect 157291 650369 157349 650403
rect 164249 650199 164283 650301
rect 173817 650199 173851 650369
rect 254041 650335 254075 650437
rect 260849 650403 260883 650505
rect 270509 650267 270543 650369
rect 280077 650199 280111 650369
rect 289829 650335 289863 650437
rect 299397 650335 299431 650505
rect 386429 650267 386463 650437
rect 389649 650267 389683 650505
rect 396089 650335 396123 650505
rect 405749 650199 405783 650301
rect 415317 650199 415351 650369
rect 425069 650335 425103 650437
rect 434637 650335 434671 650505
rect 86417 557923 86451 558433
rect 97549 558399 97583 558637
rect 86509 557651 86543 558365
rect 96905 557583 96939 558365
rect 101413 557855 101447 558705
rect 101505 558535 101539 558705
rect 129657 557855 129691 558705
rect 220737 558671 220771 558841
rect 222209 558671 222243 558841
rect 230765 558399 230799 558773
rect 231903 558229 232053 558263
rect 222209 557991 222243 558093
rect 231777 557991 231811 558161
rect 96997 557583 97031 557753
rect 122757 557651 122791 557821
rect 125149 557651 125183 557821
rect 129507 557549 129841 557583
rect 292497 557515 292531 558569
rect 302065 558535 302099 558977
rect 302157 558671 302191 558909
rect 302249 558671 302283 558909
rect 302341 558535 302375 558977
rect 302249 558467 302283 558501
rect 302433 558467 302467 558909
rect 311817 558603 311851 558909
rect 334173 558671 334207 558841
rect 345857 558671 345891 558705
rect 345581 558637 345891 558671
rect 302249 558433 302467 558467
rect 320833 558263 320867 558501
rect 345581 558467 345615 558637
rect 345673 558467 345707 558569
rect 344661 558263 344695 558433
rect 422953 558195 422987 558569
rect 432613 558195 432647 558569
rect 432797 558127 432831 558637
rect 418169 558093 418353 558127
rect 418169 557787 418203 558093
rect 418261 558025 418445 558059
rect 418261 557719 418295 558025
rect 418445 557583 418479 557753
rect 432521 557719 432555 558025
rect 432705 557787 432739 558093
rect 441629 557787 441663 558569
rect 418295 557549 418479 557583
rect 432613 557583 432647 557753
rect 441721 557719 441755 558637
rect 443561 557991 443595 558705
rect 451841 558535 451875 558773
rect 451933 558603 451967 558773
rect 480269 558671 480303 558773
rect 447149 557651 447183 558501
rect 452209 557991 452243 558637
rect 449081 557583 449115 557889
rect 452301 557855 452335 558501
rect 453313 557651 453347 558569
rect 456717 557583 456751 558433
rect 458189 557855 458223 557889
rect 458189 557821 458373 557855
rect 462513 557583 462547 558637
rect 475393 558467 475427 558569
rect 468861 557991 468895 558433
rect 475301 557991 475335 558433
rect 468711 557957 468895 557991
rect 475209 557583 475243 557957
rect 145481 542487 145515 543677
rect 152381 542419 152415 543541
rect 152473 542555 152507 543677
rect 282009 410567 282043 412233
rect 60289 318087 60323 318801
rect 61025 318563 61059 318801
rect 142813 318665 142997 318699
rect 142813 318631 142847 318665
rect 60783 318461 60875 318495
rect 60841 318291 60875 318461
rect 60749 318189 60933 318223
rect 60749 318087 60783 318189
rect 60691 318053 60783 318087
rect 115949 317679 115983 317781
rect 66821 299523 66855 309077
rect 74457 299523 74491 309077
rect 75009 299523 75043 302345
rect 77585 299523 77619 309077
rect 72249 289867 72283 292621
rect 74457 280211 74491 298061
rect 74917 289867 74951 299353
rect 80253 296735 80287 301529
rect 85957 298163 85991 307717
rect 95433 299523 95467 309077
rect 124413 307887 124447 318257
rect 138029 317883 138063 317985
rect 143641 317951 143675 318597
rect 125609 317611 125643 317713
rect 126989 317475 127023 317645
rect 135453 317339 135487 317577
rect 138121 317543 138155 317849
rect 137845 317407 137879 317509
rect 138581 317475 138615 317713
rect 140697 317645 140881 317679
rect 140697 317543 140731 317645
rect 143549 317543 143583 317917
rect 145665 317679 145699 318665
rect 147539 317985 147631 318019
rect 146677 317679 146711 317917
rect 146677 317645 147539 317679
rect 147505 317611 147539 317645
rect 147413 317407 147447 317577
rect 147597 317475 147631 317985
rect 147781 317747 147815 317985
rect 149805 317951 149839 318665
rect 152473 318631 152507 318801
rect 151461 317815 151495 317985
rect 152197 317883 152231 317985
rect 152381 317951 152415 318597
rect 147723 317713 147815 317747
rect 147873 317407 147907 317645
rect 147965 317577 148425 317611
rect 147965 317543 147999 317577
rect 151369 317543 151403 317781
rect 152473 317747 152507 318121
rect 152657 317679 152691 318053
rect 152749 317883 152783 318053
rect 155325 317543 155359 317781
rect 155417 317543 155451 318597
rect 135085 309179 135119 311933
rect 160753 309179 160787 318461
rect 169769 318155 169803 318325
rect 219265 318019 219299 318733
rect 162133 317679 162167 317917
rect 189917 317611 189951 317781
rect 229017 317611 229051 317917
rect 248613 317747 248647 318121
rect 268393 317883 268427 318053
rect 271521 317883 271555 318461
rect 277317 318087 277351 318461
rect 248521 317611 248555 317713
rect 124229 298231 124263 307717
rect 134993 299523 135027 302209
rect 124413 292451 124447 298061
rect 74917 280211 74951 289697
rect 66545 270555 66579 280109
rect 72249 270555 72283 280109
rect 77585 270555 77619 282897
rect 81725 278783 81759 283577
rect 134901 280211 134935 289765
rect 95617 270555 95651 280109
rect 124413 273955 124447 280109
rect 66545 251243 66579 260797
rect 72249 251243 72283 260797
rect 75009 251243 75043 260797
rect 77585 251243 77619 260797
rect 95617 251243 95651 260797
rect 124321 259471 124355 263585
rect 134901 260899 134935 270453
rect 134901 241519 134935 251141
rect 124321 222207 124355 224961
rect 134901 222207 134935 224961
rect 124321 202895 124355 205649
rect 134901 202895 134935 205649
rect 124321 183583 124355 186337
rect 124321 164271 124355 167025
rect 74457 153255 74491 162809
rect 78873 153255 78907 162809
rect 135085 154615 135119 157437
rect 140881 157335 140915 164169
rect 150265 157335 150299 164169
rect 135085 144959 135119 147645
rect 74457 133943 74491 143497
rect 75009 133943 75043 143497
rect 140881 137955 140915 144857
rect 150265 137955 150299 144857
rect 72249 113203 72283 122757
rect 75009 117283 75043 122757
rect 134993 114563 135027 124117
rect 140881 118643 140915 125545
rect 150265 118643 150299 125545
rect 77585 104907 77619 114461
rect 72249 92531 72283 102085
rect 74457 95251 74491 104805
rect 78781 95251 78815 104805
rect 85957 95251 85991 104805
rect 66361 77299 66395 86921
rect 75009 84303 75043 93789
rect 134993 89675 135027 104805
rect 140881 99331 140915 106233
rect 150265 99331 150299 106233
rect 66361 70295 66395 77129
rect 75009 74579 75043 84133
rect 85865 77299 85899 86921
rect 95433 77299 95467 86921
rect 140881 77299 140915 86921
rect 150265 77299 150299 86921
rect 160753 77299 160787 86853
rect 74825 66283 74859 71077
rect 81633 70295 81667 77197
rect 95433 70295 95467 77129
rect 140881 67643 140915 77129
rect 66545 48331 66579 57885
rect 72433 56559 72467 64821
rect 74457 56627 74491 66181
rect 74825 55267 74859 64821
rect 72341 45679 72375 55165
rect 77493 48399 77527 66181
rect 95617 48331 95651 57885
rect 124413 46971 124447 56525
rect 140881 51051 140915 57885
rect 150265 48331 150299 57885
rect 66545 29019 66579 38573
rect 72341 31739 72375 45509
rect 74457 37315 74491 46869
rect 75009 37247 75043 45509
rect 78873 29019 78907 38573
rect 95617 29019 95651 38573
rect 140881 31739 140915 38573
rect 150265 29019 150299 38573
rect 66637 9707 66671 19261
rect 74273 9707 74307 27557
rect 74917 9707 74951 27557
rect 95709 9707 95743 19261
rect 134901 18003 134935 27557
rect 66269 4199 66303 5185
rect 30389 3383 30423 4029
rect 35909 3111 35943 4029
rect 40693 3179 40727 4097
rect 55229 4063 55263 4165
rect 60933 4131 60967 4165
rect 60783 4097 60967 4131
rect 66637 4131 66671 4233
rect 45477 3111 45511 4029
rect 64705 3689 65165 3723
rect 64705 3587 64739 3689
rect 65717 3315 65751 3349
rect 65567 3281 65751 3315
rect 69213 3315 69247 3961
rect 54125 2907 54159 3145
rect 70409 3043 70443 4097
rect 75377 4063 75411 4165
rect 74215 3893 74399 3927
rect 74365 3859 74399 3893
rect 75101 3723 75135 4029
rect 75285 3791 75319 3893
rect 70593 3247 70627 3349
rect 74917 3213 75009 3247
rect 70501 3043 70535 3213
rect 74917 3111 74951 3213
rect 75009 2839 75043 3077
rect 75101 2839 75135 3417
rect 79425 3383 79459 3961
rect 80069 3859 80103 4029
rect 79517 3111 79551 3757
rect 81265 3383 81299 3893
rect 81357 3723 81391 3893
rect 86969 3451 87003 4777
rect 120825 3723 120859 3893
rect 122021 3791 122055 4165
rect 133153 3791 133187 3893
rect 120733 3383 120767 3689
rect 123309 3655 123343 3757
rect 133061 3723 133095 3757
rect 133245 3723 133279 3893
rect 131347 3689 131589 3723
rect 133061 3689 133279 3723
rect 123309 3621 123493 3655
rect 112453 3349 112637 3383
rect 112453 3315 112487 3349
rect 126713 2839 126747 3689
rect 127909 3383 127943 3621
rect 133153 3111 133187 3417
rect 133889 2839 133923 3689
rect 137477 3587 137511 3893
rect 137569 2839 137603 3893
rect 140881 595 140915 9605
rect 148275 4097 148367 4131
rect 141801 3111 141835 3553
rect 141893 3451 141927 3553
rect 141985 2907 142019 3417
rect 142813 3043 142847 3281
rect 143457 3179 143491 4029
rect 148333 3723 148367 4097
rect 161857 4097 162041 4131
rect 161857 4063 161891 4097
rect 161983 4029 162133 4063
rect 175933 3961 176577 3995
rect 148241 3383 148275 3689
rect 156521 3247 156555 3689
rect 147689 3111 147723 3213
rect 152473 3179 152507 3213
rect 152473 3145 152841 3179
rect 157993 2975 158027 3145
rect 159373 2907 159407 3825
rect 169861 3791 169895 3893
rect 162041 3757 162259 3791
rect 169861 3757 170045 3791
rect 162041 3723 162075 3757
rect 162133 3383 162167 3689
rect 162225 3383 162259 3757
rect 171701 3723 171735 3757
rect 175933 3723 175967 3961
rect 176669 3859 176703 3961
rect 176669 3825 176887 3859
rect 171701 3689 171885 3723
rect 160511 3009 160661 3043
rect 162041 2975 162075 3077
rect 162041 2941 162225 2975
rect 165997 2907 166031 3349
rect 173173 2771 173207 3145
rect 176853 3043 176887 3825
rect 181361 3043 181395 3213
rect 181453 3179 181487 3757
rect 181545 3043 181579 6069
rect 202797 4199 202831 6885
rect 182649 3383 182683 3961
rect 185501 3247 185535 3757
rect 186237 3383 186271 3961
rect 186789 3723 186823 3961
rect 187065 3791 187099 4097
rect 187157 3723 187191 3757
rect 186789 3689 187191 3723
rect 187249 3655 187283 4029
rect 190837 3961 190929 3995
rect 193171 3961 193413 3995
rect 186329 3621 187283 3655
rect 186329 3587 186363 3621
rect 189365 3587 189399 3893
rect 190377 3655 190411 3757
rect 190837 3723 190871 3961
rect 190929 3723 190963 3825
rect 190929 3689 191113 3723
rect 185501 3213 186145 3247
rect 277961 3043 277995 3349
rect 278053 3111 278087 3349
rect 282561 3111 282595 3281
rect 278145 3043 278179 3077
rect 277961 3009 278179 3043
<< viali >>
rect 318809 650777 318843 650811
rect 183569 650641 183603 650675
rect 144929 650573 144963 650607
rect 144929 650437 144963 650471
rect 154497 650573 154531 650607
rect 176853 650505 176887 650539
rect 183569 650505 183603 650539
rect 193137 650641 193171 650675
rect 202889 650641 202923 650675
rect 202889 650505 202923 650539
rect 212457 650641 212491 650675
rect 222209 650641 222243 650675
rect 222209 650505 222243 650539
rect 231777 650641 231811 650675
rect 241529 650641 241563 650675
rect 241529 650505 241563 650539
rect 251097 650641 251131 650675
rect 318809 650641 318843 650675
rect 328377 650777 328411 650811
rect 338129 650777 338163 650811
rect 338129 650641 338163 650675
rect 347697 650777 347731 650811
rect 357449 650777 357483 650811
rect 357449 650641 357483 650675
rect 367017 650777 367051 650811
rect 454049 650777 454083 650811
rect 454049 650641 454083 650675
rect 463617 650777 463651 650811
rect 473369 650777 473403 650811
rect 473369 650641 473403 650675
rect 482937 650777 482971 650811
rect 492689 650777 492723 650811
rect 492689 650641 492723 650675
rect 502257 650777 502291 650811
rect 311817 650573 311851 650607
rect 311909 650573 311943 650607
rect 328377 650573 328411 650607
rect 331137 650573 331171 650607
rect 331229 650573 331263 650607
rect 347697 650573 347731 650607
rect 350457 650573 350491 650607
rect 350549 650573 350583 650607
rect 367017 650573 367051 650607
rect 369869 650573 369903 650607
rect 369961 650573 369995 650607
rect 447057 650573 447091 650607
rect 447149 650573 447183 650607
rect 463617 650573 463651 650607
rect 466377 650573 466411 650607
rect 466469 650573 466503 650607
rect 482937 650573 482971 650607
rect 485697 650573 485731 650607
rect 485789 650573 485823 650607
rect 502257 650573 502291 650607
rect 505109 650573 505143 650607
rect 505201 650573 505235 650607
rect 260849 650505 260883 650539
rect 193137 650437 193171 650471
rect 195897 650437 195931 650471
rect 195989 650437 196023 650471
rect 212457 650437 212491 650471
rect 215217 650437 215251 650471
rect 215309 650437 215343 650471
rect 231777 650437 231811 650471
rect 234537 650437 234571 650471
rect 234629 650437 234663 650471
rect 251097 650437 251131 650471
rect 253857 650437 253891 650471
rect 154497 650369 154531 650403
rect 157257 650369 157291 650403
rect 157349 650369 157383 650403
rect 173817 650369 173851 650403
rect 176853 650369 176887 650403
rect 164249 650301 164283 650335
rect 164249 650165 164283 650199
rect 299397 650505 299431 650539
rect 289829 650437 289863 650471
rect 260849 650369 260883 650403
rect 270509 650369 270543 650403
rect 254041 650301 254075 650335
rect 270509 650233 270543 650267
rect 280077 650369 280111 650403
rect 173817 650165 173851 650199
rect 289829 650301 289863 650335
rect 389649 650505 389683 650539
rect 299397 650301 299431 650335
rect 386429 650437 386463 650471
rect 386429 650233 386463 650267
rect 396089 650505 396123 650539
rect 434637 650505 434671 650539
rect 425069 650437 425103 650471
rect 415317 650369 415351 650403
rect 396089 650301 396123 650335
rect 405749 650301 405783 650335
rect 389649 650233 389683 650267
rect 280077 650165 280111 650199
rect 405749 650165 405783 650199
rect 425069 650301 425103 650335
rect 434637 650301 434671 650335
rect 415317 650165 415351 650199
rect 302065 558977 302099 559011
rect 220737 558841 220771 558875
rect 101413 558705 101447 558739
rect 97549 558637 97583 558671
rect 86417 558433 86451 558467
rect 86417 557889 86451 557923
rect 86509 558365 86543 558399
rect 86509 557617 86543 557651
rect 96905 558365 96939 558399
rect 97549 558365 97583 558399
rect 101505 558705 101539 558739
rect 101505 558501 101539 558535
rect 129657 558705 129691 558739
rect 220737 558637 220771 558671
rect 222209 558841 222243 558875
rect 222209 558637 222243 558671
rect 230765 558773 230799 558807
rect 230765 558365 230799 558399
rect 292497 558569 292531 558603
rect 231869 558229 231903 558263
rect 232053 558229 232087 558263
rect 231777 558161 231811 558195
rect 222209 558093 222243 558127
rect 222209 557957 222243 557991
rect 231777 557957 231811 557991
rect 101413 557821 101447 557855
rect 122757 557821 122791 557855
rect 96905 557549 96939 557583
rect 96997 557753 97031 557787
rect 122757 557617 122791 557651
rect 125149 557821 125183 557855
rect 129657 557821 129691 557855
rect 125149 557617 125183 557651
rect 96997 557549 97031 557583
rect 129473 557549 129507 557583
rect 129841 557549 129875 557583
rect 302341 558977 302375 559011
rect 302157 558909 302191 558943
rect 302157 558637 302191 558671
rect 302249 558909 302283 558943
rect 302249 558637 302283 558671
rect 302065 558501 302099 558535
rect 302249 558501 302283 558535
rect 302341 558501 302375 558535
rect 302433 558909 302467 558943
rect 311817 558909 311851 558943
rect 334173 558841 334207 558875
rect 451841 558773 451875 558807
rect 345857 558705 345891 558739
rect 443561 558705 443595 558739
rect 334173 558637 334207 558671
rect 432797 558637 432831 558671
rect 311817 558569 311851 558603
rect 320833 558501 320867 558535
rect 320833 558229 320867 558263
rect 344661 558433 344695 558467
rect 345581 558433 345615 558467
rect 345673 558569 345707 558603
rect 345673 558433 345707 558467
rect 422953 558569 422987 558603
rect 344661 558229 344695 558263
rect 422953 558161 422987 558195
rect 432613 558569 432647 558603
rect 432613 558161 432647 558195
rect 441721 558637 441755 558671
rect 418353 558093 418387 558127
rect 432705 558093 432739 558127
rect 432797 558093 432831 558127
rect 441629 558569 441663 558603
rect 418169 557753 418203 557787
rect 418445 558025 418479 558059
rect 432521 558025 432555 558059
rect 418261 557685 418295 557719
rect 418445 557753 418479 557787
rect 432521 557685 432555 557719
rect 432613 557753 432647 557787
rect 432705 557753 432739 557787
rect 441629 557753 441663 557787
rect 418261 557549 418295 557583
rect 451933 558773 451967 558807
rect 480269 558773 480303 558807
rect 451933 558569 451967 558603
rect 452209 558637 452243 558671
rect 443561 557957 443595 557991
rect 447149 558501 447183 558535
rect 451841 558501 451875 558535
rect 441721 557685 441755 557719
rect 462513 558637 462547 558671
rect 480269 558637 480303 558671
rect 453313 558569 453347 558603
rect 452209 557957 452243 557991
rect 452301 558501 452335 558535
rect 447149 557617 447183 557651
rect 449081 557889 449115 557923
rect 432613 557549 432647 557583
rect 452301 557821 452335 557855
rect 453313 557617 453347 557651
rect 456717 558433 456751 558467
rect 449081 557549 449115 557583
rect 458189 557889 458223 557923
rect 458373 557821 458407 557855
rect 456717 557549 456751 557583
rect 475393 558569 475427 558603
rect 468861 558433 468895 558467
rect 475301 558433 475335 558467
rect 475393 558433 475427 558467
rect 468677 557957 468711 557991
rect 475209 557957 475243 557991
rect 475301 557957 475335 557991
rect 462513 557549 462547 557583
rect 475209 557549 475243 557583
rect 292497 557481 292531 557515
rect 145481 543677 145515 543711
rect 152473 543677 152507 543711
rect 145481 542453 145515 542487
rect 152381 543541 152415 543575
rect 152473 542521 152507 542555
rect 152381 542385 152415 542419
rect 282009 412233 282043 412267
rect 282009 410533 282043 410567
rect 60289 318801 60323 318835
rect 61025 318801 61059 318835
rect 152473 318801 152507 318835
rect 142997 318665 143031 318699
rect 145665 318665 145699 318699
rect 142813 318597 142847 318631
rect 143641 318597 143675 318631
rect 61025 318529 61059 318563
rect 60749 318461 60783 318495
rect 60841 318257 60875 318291
rect 124413 318257 124447 318291
rect 60933 318189 60967 318223
rect 60289 318053 60323 318087
rect 60657 318053 60691 318087
rect 115949 317781 115983 317815
rect 115949 317645 115983 317679
rect 66821 309077 66855 309111
rect 66821 299489 66855 299523
rect 74457 309077 74491 309111
rect 77585 309077 77619 309111
rect 74457 299489 74491 299523
rect 75009 302345 75043 302379
rect 75009 299489 75043 299523
rect 95433 309077 95467 309111
rect 85957 307717 85991 307751
rect 77585 299489 77619 299523
rect 80253 301529 80287 301563
rect 74917 299353 74951 299387
rect 74457 298061 74491 298095
rect 72249 292621 72283 292655
rect 72249 289833 72283 289867
rect 138029 317985 138063 318019
rect 143549 317917 143583 317951
rect 143641 317917 143675 317951
rect 138029 317849 138063 317883
rect 138121 317849 138155 317883
rect 125609 317713 125643 317747
rect 125609 317577 125643 317611
rect 126989 317645 127023 317679
rect 126989 317441 127023 317475
rect 135453 317577 135487 317611
rect 137845 317509 137879 317543
rect 138121 317509 138155 317543
rect 138581 317713 138615 317747
rect 140881 317645 140915 317679
rect 140697 317509 140731 317543
rect 149805 318665 149839 318699
rect 147505 317985 147539 318019
rect 145665 317645 145699 317679
rect 146677 317917 146711 317951
rect 143549 317509 143583 317543
rect 147413 317577 147447 317611
rect 147505 317577 147539 317611
rect 138581 317441 138615 317475
rect 137845 317373 137879 317407
rect 147781 317985 147815 318019
rect 219265 318733 219299 318767
rect 152381 318597 152415 318631
rect 152473 318597 152507 318631
rect 155417 318597 155451 318631
rect 149805 317917 149839 317951
rect 151461 317985 151495 318019
rect 152197 317985 152231 318019
rect 152381 317917 152415 317951
rect 152473 318121 152507 318155
rect 152197 317849 152231 317883
rect 147689 317713 147723 317747
rect 151369 317781 151403 317815
rect 151461 317781 151495 317815
rect 147597 317441 147631 317475
rect 147873 317645 147907 317679
rect 147413 317373 147447 317407
rect 148425 317577 148459 317611
rect 147965 317509 147999 317543
rect 152473 317713 152507 317747
rect 152657 318053 152691 318087
rect 152749 318053 152783 318087
rect 152749 317849 152783 317883
rect 152657 317645 152691 317679
rect 155325 317781 155359 317815
rect 151369 317509 151403 317543
rect 155325 317509 155359 317543
rect 155417 317509 155451 317543
rect 160753 318461 160787 318495
rect 147873 317373 147907 317407
rect 135453 317305 135487 317339
rect 135085 311933 135119 311967
rect 135085 309145 135119 309179
rect 169769 318325 169803 318359
rect 169769 318121 169803 318155
rect 271521 318461 271555 318495
rect 219265 317985 219299 318019
rect 248613 318121 248647 318155
rect 162133 317917 162167 317951
rect 229017 317917 229051 317951
rect 162133 317645 162167 317679
rect 189917 317781 189951 317815
rect 189917 317577 189951 317611
rect 268393 318053 268427 318087
rect 268393 317849 268427 317883
rect 277317 318461 277351 318495
rect 277317 318053 277351 318087
rect 271521 317849 271555 317883
rect 229017 317577 229051 317611
rect 248521 317713 248555 317747
rect 248613 317713 248647 317747
rect 248521 317577 248555 317611
rect 160753 309145 160787 309179
rect 124413 307853 124447 307887
rect 95433 299489 95467 299523
rect 124229 307717 124263 307751
rect 134993 302209 135027 302243
rect 134993 299489 135027 299523
rect 124229 298197 124263 298231
rect 85957 298129 85991 298163
rect 80253 296701 80287 296735
rect 124413 298061 124447 298095
rect 124413 292417 124447 292451
rect 74917 289833 74951 289867
rect 134901 289765 134935 289799
rect 74457 280177 74491 280211
rect 74917 289697 74951 289731
rect 81725 283577 81759 283611
rect 74917 280177 74951 280211
rect 77585 282897 77619 282931
rect 66545 280109 66579 280143
rect 66545 270521 66579 270555
rect 72249 280109 72283 280143
rect 72249 270521 72283 270555
rect 134901 280177 134935 280211
rect 81725 278749 81759 278783
rect 95617 280109 95651 280143
rect 77585 270521 77619 270555
rect 124413 280109 124447 280143
rect 124413 273921 124447 273955
rect 95617 270521 95651 270555
rect 134901 270453 134935 270487
rect 124321 263585 124355 263619
rect 66545 260797 66579 260831
rect 66545 251209 66579 251243
rect 72249 260797 72283 260831
rect 72249 251209 72283 251243
rect 75009 260797 75043 260831
rect 75009 251209 75043 251243
rect 77585 260797 77619 260831
rect 77585 251209 77619 251243
rect 95617 260797 95651 260831
rect 134901 260865 134935 260899
rect 124321 259437 124355 259471
rect 95617 251209 95651 251243
rect 134901 251141 134935 251175
rect 134901 241485 134935 241519
rect 124321 224961 124355 224995
rect 124321 222173 124355 222207
rect 134901 224961 134935 224995
rect 134901 222173 134935 222207
rect 124321 205649 124355 205683
rect 124321 202861 124355 202895
rect 134901 205649 134935 205683
rect 134901 202861 134935 202895
rect 124321 186337 124355 186371
rect 124321 183549 124355 183583
rect 124321 167025 124355 167059
rect 124321 164237 124355 164271
rect 140881 164169 140915 164203
rect 74457 162809 74491 162843
rect 74457 153221 74491 153255
rect 78873 162809 78907 162843
rect 135085 157437 135119 157471
rect 140881 157301 140915 157335
rect 150265 164169 150299 164203
rect 150265 157301 150299 157335
rect 135085 154581 135119 154615
rect 78873 153221 78907 153255
rect 135085 147645 135119 147679
rect 135085 144925 135119 144959
rect 140881 144857 140915 144891
rect 74457 143497 74491 143531
rect 74457 133909 74491 133943
rect 75009 143497 75043 143531
rect 140881 137921 140915 137955
rect 150265 144857 150299 144891
rect 150265 137921 150299 137955
rect 75009 133909 75043 133943
rect 140881 125545 140915 125579
rect 134993 124117 135027 124151
rect 72249 122757 72283 122791
rect 75009 122757 75043 122791
rect 75009 117249 75043 117283
rect 140881 118609 140915 118643
rect 150265 125545 150299 125579
rect 150265 118609 150299 118643
rect 134993 114529 135027 114563
rect 72249 113169 72283 113203
rect 77585 114461 77619 114495
rect 77585 104873 77619 104907
rect 140881 106233 140915 106267
rect 74457 104805 74491 104839
rect 72249 102085 72283 102119
rect 74457 95217 74491 95251
rect 78781 104805 78815 104839
rect 78781 95217 78815 95251
rect 85957 104805 85991 104839
rect 85957 95217 85991 95251
rect 134993 104805 135027 104839
rect 72249 92497 72283 92531
rect 75009 93789 75043 93823
rect 66361 86921 66395 86955
rect 140881 99297 140915 99331
rect 150265 106233 150299 106267
rect 150265 99297 150299 99331
rect 134993 89641 135027 89675
rect 75009 84269 75043 84303
rect 85865 86921 85899 86955
rect 66361 77265 66395 77299
rect 75009 84133 75043 84167
rect 66361 77129 66395 77163
rect 85865 77265 85899 77299
rect 95433 86921 95467 86955
rect 95433 77265 95467 77299
rect 140881 86921 140915 86955
rect 140881 77265 140915 77299
rect 150265 86921 150299 86955
rect 150265 77265 150299 77299
rect 160753 86853 160787 86887
rect 160753 77265 160787 77299
rect 75009 74545 75043 74579
rect 81633 77197 81667 77231
rect 66361 70261 66395 70295
rect 74825 71077 74859 71111
rect 81633 70261 81667 70295
rect 95433 77129 95467 77163
rect 95433 70261 95467 70295
rect 140881 77129 140915 77163
rect 140881 67609 140915 67643
rect 74825 66249 74859 66283
rect 74457 66181 74491 66215
rect 72433 64821 72467 64855
rect 66545 57885 66579 57919
rect 77493 66181 77527 66215
rect 74457 56593 74491 56627
rect 74825 64821 74859 64855
rect 72433 56525 72467 56559
rect 74825 55233 74859 55267
rect 66545 48297 66579 48331
rect 72341 55165 72375 55199
rect 77493 48365 77527 48399
rect 95617 57885 95651 57919
rect 140881 57885 140915 57919
rect 95617 48297 95651 48331
rect 124413 56525 124447 56559
rect 140881 51017 140915 51051
rect 150265 57885 150299 57919
rect 150265 48297 150299 48331
rect 124413 46937 124447 46971
rect 72341 45645 72375 45679
rect 74457 46869 74491 46903
rect 72341 45509 72375 45543
rect 66545 38573 66579 38607
rect 74457 37281 74491 37315
rect 75009 45509 75043 45543
rect 75009 37213 75043 37247
rect 78873 38573 78907 38607
rect 72341 31705 72375 31739
rect 66545 28985 66579 29019
rect 78873 28985 78907 29019
rect 95617 38573 95651 38607
rect 140881 38573 140915 38607
rect 140881 31705 140915 31739
rect 150265 38573 150299 38607
rect 95617 28985 95651 29019
rect 150265 28985 150299 29019
rect 74273 27557 74307 27591
rect 66637 19261 66671 19295
rect 66637 9673 66671 9707
rect 74273 9673 74307 9707
rect 74917 27557 74951 27591
rect 134901 27557 134935 27591
rect 74917 9673 74951 9707
rect 95709 19261 95743 19295
rect 134901 17969 134935 18003
rect 95709 9673 95743 9707
rect 140881 9605 140915 9639
rect 66269 5185 66303 5219
rect 86969 4777 87003 4811
rect 55229 4165 55263 4199
rect 40693 4097 40727 4131
rect 30389 4029 30423 4063
rect 30389 3349 30423 3383
rect 35909 4029 35943 4063
rect 60933 4165 60967 4199
rect 66269 4165 66303 4199
rect 66637 4233 66671 4267
rect 60749 4097 60783 4131
rect 75377 4165 75411 4199
rect 66637 4097 66671 4131
rect 70409 4097 70443 4131
rect 40693 3145 40727 3179
rect 45477 4029 45511 4063
rect 55229 4029 55263 4063
rect 35909 3077 35943 3111
rect 69213 3961 69247 3995
rect 65165 3689 65199 3723
rect 64705 3553 64739 3587
rect 65717 3349 65751 3383
rect 65533 3281 65567 3315
rect 69213 3281 69247 3315
rect 45477 3077 45511 3111
rect 54125 3145 54159 3179
rect 75101 4029 75135 4063
rect 75377 4029 75411 4063
rect 80069 4029 80103 4063
rect 74181 3893 74215 3927
rect 74365 3825 74399 3859
rect 79425 3961 79459 3995
rect 75285 3893 75319 3927
rect 75285 3757 75319 3791
rect 75101 3689 75135 3723
rect 75101 3417 75135 3451
rect 70593 3349 70627 3383
rect 70409 3009 70443 3043
rect 70501 3213 70535 3247
rect 70593 3213 70627 3247
rect 75009 3213 75043 3247
rect 74917 3077 74951 3111
rect 75009 3077 75043 3111
rect 70501 3009 70535 3043
rect 54125 2873 54159 2907
rect 75009 2805 75043 2839
rect 80069 3825 80103 3859
rect 81265 3893 81299 3927
rect 79425 3349 79459 3383
rect 79517 3757 79551 3791
rect 81357 3893 81391 3927
rect 81357 3689 81391 3723
rect 122021 4165 122055 4199
rect 120825 3893 120859 3927
rect 133153 3893 133187 3927
rect 122021 3757 122055 3791
rect 123309 3757 123343 3791
rect 86969 3417 87003 3451
rect 120733 3689 120767 3723
rect 120825 3689 120859 3723
rect 133061 3757 133095 3791
rect 133153 3757 133187 3791
rect 133245 3893 133279 3927
rect 137477 3893 137511 3927
rect 126713 3689 126747 3723
rect 131313 3689 131347 3723
rect 131589 3689 131623 3723
rect 133889 3689 133923 3723
rect 123493 3621 123527 3655
rect 81265 3349 81299 3383
rect 112637 3349 112671 3383
rect 120733 3349 120767 3383
rect 112453 3281 112487 3315
rect 79517 3077 79551 3111
rect 75101 2805 75135 2839
rect 127909 3621 127943 3655
rect 127909 3349 127943 3383
rect 133153 3417 133187 3451
rect 133153 3077 133187 3111
rect 126713 2805 126747 2839
rect 137477 3553 137511 3587
rect 137569 3893 137603 3927
rect 133889 2805 133923 2839
rect 137569 2805 137603 2839
rect 202797 6885 202831 6919
rect 181545 6069 181579 6103
rect 148241 4097 148275 4131
rect 143457 4029 143491 4063
rect 141801 3553 141835 3587
rect 141893 3553 141927 3587
rect 141893 3417 141927 3451
rect 141985 3417 142019 3451
rect 141801 3077 141835 3111
rect 142813 3281 142847 3315
rect 162041 4097 162075 4131
rect 161857 4029 161891 4063
rect 161949 4029 161983 4063
rect 162133 4029 162167 4063
rect 176577 3961 176611 3995
rect 176669 3961 176703 3995
rect 169861 3893 169895 3927
rect 159373 3825 159407 3859
rect 148241 3689 148275 3723
rect 148333 3689 148367 3723
rect 156521 3689 156555 3723
rect 148241 3349 148275 3383
rect 143457 3145 143491 3179
rect 147689 3213 147723 3247
rect 152473 3213 152507 3247
rect 156521 3213 156555 3247
rect 152841 3145 152875 3179
rect 157993 3145 158027 3179
rect 147689 3077 147723 3111
rect 142813 3009 142847 3043
rect 157993 2941 158027 2975
rect 141985 2873 142019 2907
rect 170045 3757 170079 3791
rect 171701 3757 171735 3791
rect 162041 3689 162075 3723
rect 162133 3689 162167 3723
rect 162133 3349 162167 3383
rect 171885 3689 171919 3723
rect 175933 3689 175967 3723
rect 162225 3349 162259 3383
rect 165997 3349 166031 3383
rect 162041 3077 162075 3111
rect 160477 3009 160511 3043
rect 160661 3009 160695 3043
rect 162225 2941 162259 2975
rect 159373 2873 159407 2907
rect 165997 2873 166031 2907
rect 173173 3145 173207 3179
rect 181453 3757 181487 3791
rect 176853 3009 176887 3043
rect 181361 3213 181395 3247
rect 181453 3145 181487 3179
rect 181361 3009 181395 3043
rect 202797 4165 202831 4199
rect 187065 4097 187099 4131
rect 182649 3961 182683 3995
rect 186237 3961 186271 3995
rect 182649 3349 182683 3383
rect 185501 3757 185535 3791
rect 186789 3961 186823 3995
rect 187249 4029 187283 4063
rect 187065 3757 187099 3791
rect 187157 3757 187191 3791
rect 190929 3961 190963 3995
rect 193137 3961 193171 3995
rect 193413 3961 193447 3995
rect 189365 3893 189399 3927
rect 186329 3553 186363 3587
rect 190377 3757 190411 3791
rect 190837 3689 190871 3723
rect 190929 3825 190963 3859
rect 191113 3689 191147 3723
rect 190377 3621 190411 3655
rect 189365 3553 189399 3587
rect 186237 3349 186271 3383
rect 277961 3349 277995 3383
rect 186145 3213 186179 3247
rect 181545 3009 181579 3043
rect 278053 3349 278087 3383
rect 282561 3281 282595 3315
rect 278053 3077 278087 3111
rect 278145 3077 278179 3111
rect 282561 3077 282595 3111
rect 173173 2737 173207 2771
rect 140881 561 140915 595
<< metal1 >>
rect 264882 653352 264888 653404
rect 264940 653392 264946 653404
rect 378134 653392 378140 653404
rect 264940 653364 378140 653392
rect 264940 653352 264946 653364
rect 378134 653352 378140 653364
rect 378192 653352 378198 653404
rect 383562 653352 383568 653404
rect 383620 653392 383626 653404
rect 508406 653392 508412 653404
rect 383620 653364 508412 653392
rect 383620 653352 383626 653364
rect 508406 653352 508412 653364
rect 508464 653352 508470 653404
rect 259178 652876 259184 652928
rect 259236 652916 259242 652928
rect 263594 652916 263600 652928
rect 259236 652888 263600 652916
rect 259236 652876 259242 652888
rect 263594 652876 263600 652888
rect 263652 652916 263658 652928
rect 264882 652916 264888 652928
rect 263652 652888 264888 652916
rect 263652 652876 263658 652888
rect 264882 652876 264888 652888
rect 264940 652876 264946 652928
rect 378134 652876 378140 652928
rect 378192 652916 378198 652928
rect 383562 652916 383568 652928
rect 378192 652888 383568 652916
rect 378192 652876 378198 652888
rect 383562 652876 383568 652888
rect 383620 652876 383626 652928
rect 508406 652808 508412 652860
rect 508464 652848 508470 652860
rect 513374 652848 513380 652860
rect 508464 652820 513380 652848
rect 508464 652808 508470 652820
rect 513374 652808 513380 652820
rect 513432 652808 513438 652860
rect 129274 652740 129280 652792
rect 129332 652780 129338 652792
rect 133690 652780 133696 652792
rect 129332 652752 133696 652780
rect 129332 652740 129338 652752
rect 133690 652740 133696 652752
rect 133748 652780 133754 652792
rect 139394 652780 139400 652792
rect 133748 652752 139400 652780
rect 133748 652740 133754 652752
rect 139394 652740 139400 652752
rect 139452 652740 139458 652792
rect 513392 652780 513420 652808
rect 518894 652780 518900 652792
rect 513392 652752 518900 652780
rect 518894 652740 518900 652752
rect 518952 652740 518958 652792
rect 318797 650811 318855 650817
rect 318797 650777 318809 650811
rect 318843 650808 318855 650811
rect 328365 650811 328423 650817
rect 328365 650808 328377 650811
rect 318843 650780 328377 650808
rect 318843 650777 318855 650780
rect 318797 650771 318855 650777
rect 328365 650777 328377 650780
rect 328411 650777 328423 650811
rect 328365 650771 328423 650777
rect 338117 650811 338175 650817
rect 338117 650777 338129 650811
rect 338163 650808 338175 650811
rect 347685 650811 347743 650817
rect 347685 650808 347697 650811
rect 338163 650780 347697 650808
rect 338163 650777 338175 650780
rect 338117 650771 338175 650777
rect 347685 650777 347697 650780
rect 347731 650777 347743 650811
rect 347685 650771 347743 650777
rect 357437 650811 357495 650817
rect 357437 650777 357449 650811
rect 357483 650808 357495 650811
rect 367005 650811 367063 650817
rect 367005 650808 367017 650811
rect 357483 650780 367017 650808
rect 357483 650777 357495 650780
rect 357437 650771 357495 650777
rect 367005 650777 367017 650780
rect 367051 650777 367063 650811
rect 367005 650771 367063 650777
rect 454037 650811 454095 650817
rect 454037 650777 454049 650811
rect 454083 650808 454095 650811
rect 463605 650811 463663 650817
rect 463605 650808 463617 650811
rect 454083 650780 463617 650808
rect 454083 650777 454095 650780
rect 454037 650771 454095 650777
rect 463605 650777 463617 650780
rect 463651 650777 463663 650811
rect 463605 650771 463663 650777
rect 473357 650811 473415 650817
rect 473357 650777 473369 650811
rect 473403 650808 473415 650811
rect 482925 650811 482983 650817
rect 482925 650808 482937 650811
rect 473403 650780 482937 650808
rect 473403 650777 473415 650780
rect 473357 650771 473415 650777
rect 482925 650777 482937 650780
rect 482971 650777 482983 650811
rect 482925 650771 482983 650777
rect 492677 650811 492735 650817
rect 492677 650777 492689 650811
rect 492723 650808 492735 650811
rect 502245 650811 502303 650817
rect 502245 650808 502257 650811
rect 492723 650780 502257 650808
rect 492723 650777 492735 650780
rect 492677 650771 492735 650777
rect 502245 650777 502257 650780
rect 502291 650777 502303 650811
rect 502245 650771 502303 650777
rect 183557 650675 183615 650681
rect 183557 650641 183569 650675
rect 183603 650672 183615 650675
rect 193125 650675 193183 650681
rect 193125 650672 193137 650675
rect 183603 650644 193137 650672
rect 183603 650641 183615 650644
rect 183557 650635 183615 650641
rect 193125 650641 193137 650644
rect 193171 650641 193183 650675
rect 193125 650635 193183 650641
rect 202877 650675 202935 650681
rect 202877 650641 202889 650675
rect 202923 650672 202935 650675
rect 212445 650675 212503 650681
rect 212445 650672 212457 650675
rect 202923 650644 212457 650672
rect 202923 650641 202935 650644
rect 202877 650635 202935 650641
rect 212445 650641 212457 650644
rect 212491 650641 212503 650675
rect 212445 650635 212503 650641
rect 222197 650675 222255 650681
rect 222197 650641 222209 650675
rect 222243 650672 222255 650675
rect 231765 650675 231823 650681
rect 231765 650672 231777 650675
rect 222243 650644 231777 650672
rect 222243 650641 222255 650644
rect 222197 650635 222255 650641
rect 231765 650641 231777 650644
rect 231811 650641 231823 650675
rect 231765 650635 231823 650641
rect 241517 650675 241575 650681
rect 241517 650641 241529 650675
rect 241563 650672 241575 650675
rect 251085 650675 251143 650681
rect 251085 650672 251097 650675
rect 241563 650644 251097 650672
rect 241563 650641 241575 650644
rect 241517 650635 241575 650641
rect 251085 650641 251097 650644
rect 251131 650641 251143 650675
rect 318797 650675 318855 650681
rect 318797 650672 318809 650675
rect 251085 650635 251143 650641
rect 313108 650644 318809 650672
rect 144917 650607 144975 650613
rect 144917 650573 144929 650607
rect 144963 650604 144975 650607
rect 154485 650607 154543 650613
rect 154485 650604 154497 650607
rect 144963 650576 154497 650604
rect 144963 650573 144975 650576
rect 144917 650567 144975 650573
rect 154485 650573 154497 650576
rect 154531 650573 154543 650607
rect 311805 650607 311863 650613
rect 311805 650604 311817 650607
rect 154485 650567 154543 650573
rect 302160 650576 311817 650604
rect 176841 650539 176899 650545
rect 176841 650505 176853 650539
rect 176887 650536 176899 650539
rect 183557 650539 183615 650545
rect 183557 650536 183569 650539
rect 176887 650508 183569 650536
rect 176887 650505 176899 650508
rect 176841 650499 176899 650505
rect 183557 650505 183569 650508
rect 183603 650505 183615 650539
rect 202877 650539 202935 650545
rect 202877 650536 202889 650539
rect 183557 650499 183615 650505
rect 197188 650508 202889 650536
rect 137646 650428 137652 650480
rect 137704 650468 137710 650480
rect 144917 650471 144975 650477
rect 144917 650468 144929 650471
rect 137704 650440 144929 650468
rect 137704 650428 137710 650440
rect 144917 650437 144929 650440
rect 144963 650437 144975 650471
rect 144917 650431 144975 650437
rect 193125 650471 193183 650477
rect 193125 650437 193137 650471
rect 193171 650468 193183 650471
rect 195885 650471 195943 650477
rect 195885 650468 195897 650471
rect 193171 650440 195897 650468
rect 193171 650437 193183 650440
rect 193125 650431 193183 650437
rect 195885 650437 195897 650440
rect 195931 650437 195943 650471
rect 195885 650431 195943 650437
rect 195977 650471 196035 650477
rect 195977 650437 195989 650471
rect 196023 650468 196035 650471
rect 197188 650468 197216 650508
rect 202877 650505 202889 650508
rect 202923 650505 202935 650539
rect 222197 650539 222255 650545
rect 222197 650536 222209 650539
rect 202877 650499 202935 650505
rect 216508 650508 222209 650536
rect 196023 650440 197216 650468
rect 212445 650471 212503 650477
rect 196023 650437 196035 650440
rect 195977 650431 196035 650437
rect 212445 650437 212457 650471
rect 212491 650468 212503 650471
rect 215205 650471 215263 650477
rect 215205 650468 215217 650471
rect 212491 650440 215217 650468
rect 212491 650437 212503 650440
rect 212445 650431 212503 650437
rect 215205 650437 215217 650440
rect 215251 650437 215263 650471
rect 215205 650431 215263 650437
rect 215297 650471 215355 650477
rect 215297 650437 215309 650471
rect 215343 650468 215355 650471
rect 216508 650468 216536 650508
rect 222197 650505 222209 650508
rect 222243 650505 222255 650539
rect 241517 650539 241575 650545
rect 241517 650536 241529 650539
rect 222197 650499 222255 650505
rect 235828 650508 241529 650536
rect 215343 650440 216536 650468
rect 231765 650471 231823 650477
rect 215343 650437 215355 650440
rect 215297 650431 215355 650437
rect 231765 650437 231777 650471
rect 231811 650468 231823 650471
rect 234525 650471 234583 650477
rect 234525 650468 234537 650471
rect 231811 650440 234537 650468
rect 231811 650437 231823 650440
rect 231765 650431 231823 650437
rect 234525 650437 234537 650440
rect 234571 650437 234583 650471
rect 234525 650431 234583 650437
rect 234617 650471 234675 650477
rect 234617 650437 234629 650471
rect 234663 650468 234675 650471
rect 235828 650468 235856 650508
rect 241517 650505 241529 650508
rect 241563 650505 241575 650539
rect 241517 650499 241575 650505
rect 260837 650539 260895 650545
rect 260837 650505 260849 650539
rect 260883 650536 260895 650539
rect 266446 650536 266452 650548
rect 260883 650508 266452 650536
rect 260883 650505 260895 650508
rect 260837 650499 260895 650505
rect 266446 650496 266452 650508
rect 266504 650496 266510 650548
rect 299385 650539 299443 650545
rect 299385 650505 299397 650539
rect 299431 650536 299443 650539
rect 302160 650536 302188 650576
rect 311805 650573 311817 650576
rect 311851 650573 311863 650607
rect 311805 650567 311863 650573
rect 311897 650607 311955 650613
rect 311897 650573 311909 650607
rect 311943 650604 311955 650607
rect 313108 650604 313136 650644
rect 318797 650641 318809 650644
rect 318843 650641 318855 650675
rect 338117 650675 338175 650681
rect 338117 650672 338129 650675
rect 318797 650635 318855 650641
rect 332428 650644 338129 650672
rect 311943 650576 313136 650604
rect 328365 650607 328423 650613
rect 311943 650573 311955 650576
rect 311897 650567 311955 650573
rect 328365 650573 328377 650607
rect 328411 650604 328423 650607
rect 331125 650607 331183 650613
rect 331125 650604 331137 650607
rect 328411 650576 331137 650604
rect 328411 650573 328423 650576
rect 328365 650567 328423 650573
rect 331125 650573 331137 650576
rect 331171 650573 331183 650607
rect 331125 650567 331183 650573
rect 331217 650607 331275 650613
rect 331217 650573 331229 650607
rect 331263 650604 331275 650607
rect 332428 650604 332456 650644
rect 338117 650641 338129 650644
rect 338163 650641 338175 650675
rect 357437 650675 357495 650681
rect 357437 650672 357449 650675
rect 338117 650635 338175 650641
rect 351748 650644 357449 650672
rect 331263 650576 332456 650604
rect 347685 650607 347743 650613
rect 331263 650573 331275 650576
rect 331217 650567 331275 650573
rect 347685 650573 347697 650607
rect 347731 650604 347743 650607
rect 350445 650607 350503 650613
rect 350445 650604 350457 650607
rect 347731 650576 350457 650604
rect 347731 650573 347743 650576
rect 347685 650567 347743 650573
rect 350445 650573 350457 650576
rect 350491 650573 350503 650607
rect 350445 650567 350503 650573
rect 350537 650607 350595 650613
rect 350537 650573 350549 650607
rect 350583 650604 350595 650607
rect 351748 650604 351776 650644
rect 357437 650641 357449 650644
rect 357483 650641 357495 650675
rect 454037 650675 454095 650681
rect 454037 650672 454049 650675
rect 357437 650635 357495 650641
rect 448348 650644 454049 650672
rect 350583 650576 351776 650604
rect 367005 650607 367063 650613
rect 350583 650573 350595 650576
rect 350537 650567 350595 650573
rect 367005 650573 367017 650607
rect 367051 650604 367063 650607
rect 369857 650607 369915 650613
rect 369857 650604 369869 650607
rect 367051 650576 369869 650604
rect 367051 650573 367063 650576
rect 367005 650567 367063 650573
rect 369857 650573 369869 650576
rect 369903 650573 369915 650607
rect 369857 650567 369915 650573
rect 369949 650607 370007 650613
rect 369949 650573 369961 650607
rect 369995 650604 370007 650607
rect 447045 650607 447103 650613
rect 447045 650604 447057 650607
rect 369995 650576 376708 650604
rect 369995 650573 370007 650576
rect 369949 650567 370007 650573
rect 299431 650508 302188 650536
rect 376680 650536 376708 650576
rect 437400 650576 447057 650604
rect 389637 650539 389695 650545
rect 376680 650508 379468 650536
rect 299431 650505 299443 650508
rect 299385 650499 299443 650505
rect 234663 650440 235856 650468
rect 251085 650471 251143 650477
rect 234663 650437 234675 650440
rect 234617 650431 234675 650437
rect 251085 650437 251097 650471
rect 251131 650468 251143 650471
rect 253845 650471 253903 650477
rect 253845 650468 253857 650471
rect 251131 650440 253857 650468
rect 251131 650437 251143 650440
rect 251085 650431 251143 650437
rect 253845 650437 253857 650440
rect 253891 650437 253903 650471
rect 253845 650431 253903 650437
rect 282822 650428 282828 650480
rect 282880 650468 282886 650480
rect 289817 650471 289875 650477
rect 289817 650468 289829 650471
rect 282880 650440 289829 650468
rect 282880 650428 282886 650440
rect 289817 650437 289829 650440
rect 289863 650437 289875 650471
rect 379440 650468 379468 650508
rect 389637 650505 389649 650539
rect 389683 650536 389695 650539
rect 396077 650539 396135 650545
rect 396077 650536 396089 650539
rect 389683 650508 396089 650536
rect 389683 650505 389695 650508
rect 389637 650499 389695 650505
rect 396077 650505 396089 650508
rect 396123 650505 396135 650539
rect 396077 650499 396135 650505
rect 434625 650539 434683 650545
rect 434625 650505 434637 650539
rect 434671 650536 434683 650539
rect 437400 650536 437428 650576
rect 447045 650573 447057 650576
rect 447091 650573 447103 650607
rect 447045 650567 447103 650573
rect 447137 650607 447195 650613
rect 447137 650573 447149 650607
rect 447183 650604 447195 650607
rect 448348 650604 448376 650644
rect 454037 650641 454049 650644
rect 454083 650641 454095 650675
rect 473357 650675 473415 650681
rect 473357 650672 473369 650675
rect 454037 650635 454095 650641
rect 467668 650644 473369 650672
rect 447183 650576 448376 650604
rect 463605 650607 463663 650613
rect 447183 650573 447195 650576
rect 447137 650567 447195 650573
rect 463605 650573 463617 650607
rect 463651 650604 463663 650607
rect 466365 650607 466423 650613
rect 466365 650604 466377 650607
rect 463651 650576 466377 650604
rect 463651 650573 463663 650576
rect 463605 650567 463663 650573
rect 466365 650573 466377 650576
rect 466411 650573 466423 650607
rect 466365 650567 466423 650573
rect 466457 650607 466515 650613
rect 466457 650573 466469 650607
rect 466503 650604 466515 650607
rect 467668 650604 467696 650644
rect 473357 650641 473369 650644
rect 473403 650641 473415 650675
rect 492677 650675 492735 650681
rect 492677 650672 492689 650675
rect 473357 650635 473415 650641
rect 486988 650644 492689 650672
rect 466503 650576 467696 650604
rect 482925 650607 482983 650613
rect 466503 650573 466515 650576
rect 466457 650567 466515 650573
rect 482925 650573 482937 650607
rect 482971 650604 482983 650607
rect 485685 650607 485743 650613
rect 485685 650604 485697 650607
rect 482971 650576 485697 650604
rect 482971 650573 482983 650576
rect 482925 650567 482983 650573
rect 485685 650573 485697 650576
rect 485731 650573 485743 650607
rect 485685 650567 485743 650573
rect 485777 650607 485835 650613
rect 485777 650573 485789 650607
rect 485823 650604 485835 650607
rect 486988 650604 487016 650644
rect 492677 650641 492689 650644
rect 492723 650641 492735 650675
rect 492677 650635 492735 650641
rect 485823 650576 487016 650604
rect 502245 650607 502303 650613
rect 485823 650573 485835 650576
rect 485777 650567 485835 650573
rect 502245 650573 502257 650607
rect 502291 650604 502303 650607
rect 505097 650607 505155 650613
rect 505097 650604 505109 650607
rect 502291 650576 505109 650604
rect 502291 650573 502303 650576
rect 502245 650567 502303 650573
rect 505097 650573 505109 650576
rect 505143 650573 505155 650607
rect 505097 650567 505155 650573
rect 505189 650607 505247 650613
rect 505189 650573 505201 650607
rect 505235 650604 505247 650607
rect 505235 650576 511948 650604
rect 505235 650573 505247 650576
rect 505189 650567 505247 650573
rect 434671 650508 437428 650536
rect 511920 650536 511948 650576
rect 511920 650508 514708 650536
rect 434671 650505 434683 650508
rect 434625 650499 434683 650505
rect 386417 650471 386475 650477
rect 386417 650468 386429 650471
rect 379440 650440 386429 650468
rect 289817 650431 289875 650437
rect 386417 650437 386429 650440
rect 386463 650437 386475 650471
rect 425057 650471 425115 650477
rect 425057 650468 425069 650471
rect 386417 650431 386475 650437
rect 418080 650440 425069 650468
rect 154485 650403 154543 650409
rect 154485 650369 154497 650403
rect 154531 650400 154543 650403
rect 157245 650403 157303 650409
rect 157245 650400 157257 650403
rect 154531 650372 157257 650400
rect 154531 650369 154543 650372
rect 154485 650363 154543 650369
rect 157245 650369 157257 650372
rect 157291 650369 157303 650403
rect 157245 650363 157303 650369
rect 157337 650403 157395 650409
rect 157337 650369 157349 650403
rect 157383 650400 157395 650403
rect 173805 650403 173863 650409
rect 157383 650372 158576 650400
rect 157383 650369 157395 650372
rect 157337 650363 157395 650369
rect 158548 650332 158576 650372
rect 173805 650369 173817 650403
rect 173851 650400 173863 650403
rect 176841 650403 176899 650409
rect 176841 650400 176853 650403
rect 173851 650372 176853 650400
rect 173851 650369 173863 650372
rect 173805 650363 173863 650369
rect 176841 650369 176853 650372
rect 176887 650369 176899 650403
rect 176841 650363 176899 650369
rect 260837 650403 260895 650409
rect 260837 650369 260849 650403
rect 260883 650369 260895 650403
rect 260837 650363 260895 650369
rect 270497 650403 270555 650409
rect 270497 650369 270509 650403
rect 270543 650400 270555 650403
rect 280065 650403 280123 650409
rect 280065 650400 280077 650403
rect 270543 650372 280077 650400
rect 270543 650369 270555 650372
rect 270497 650363 270555 650369
rect 280065 650369 280077 650372
rect 280111 650369 280123 650403
rect 280065 650363 280123 650369
rect 415305 650403 415363 650409
rect 415305 650369 415317 650403
rect 415351 650400 415363 650403
rect 418080 650400 418108 650440
rect 425057 650437 425069 650440
rect 425103 650437 425115 650471
rect 514680 650468 514708 650508
rect 516410 650468 516416 650480
rect 514680 650440 516416 650468
rect 425057 650431 425115 650437
rect 516410 650428 516416 650440
rect 516468 650428 516474 650480
rect 415351 650372 418108 650400
rect 415351 650369 415363 650372
rect 415305 650363 415363 650369
rect 164237 650335 164295 650341
rect 164237 650332 164249 650335
rect 158548 650304 164249 650332
rect 164237 650301 164249 650304
rect 164283 650301 164295 650335
rect 164237 650295 164295 650301
rect 254029 650335 254087 650341
rect 254029 650301 254041 650335
rect 254075 650332 254087 650335
rect 260852 650332 260880 650363
rect 254075 650304 260880 650332
rect 289817 650335 289875 650341
rect 254075 650301 254087 650304
rect 254029 650295 254087 650301
rect 289817 650301 289829 650335
rect 289863 650332 289875 650335
rect 299385 650335 299443 650341
rect 299385 650332 299397 650335
rect 289863 650304 299397 650332
rect 289863 650301 289875 650304
rect 289817 650295 289875 650301
rect 299385 650301 299397 650304
rect 299431 650301 299443 650335
rect 299385 650295 299443 650301
rect 396077 650335 396135 650341
rect 396077 650301 396089 650335
rect 396123 650332 396135 650335
rect 405737 650335 405795 650341
rect 405737 650332 405749 650335
rect 396123 650304 405749 650332
rect 396123 650301 396135 650304
rect 396077 650295 396135 650301
rect 405737 650301 405749 650304
rect 405783 650301 405795 650335
rect 405737 650295 405795 650301
rect 425057 650335 425115 650341
rect 425057 650301 425069 650335
rect 425103 650332 425115 650335
rect 434625 650335 434683 650341
rect 434625 650332 434637 650335
rect 425103 650304 434637 650332
rect 425103 650301 425115 650304
rect 425057 650295 425115 650301
rect 434625 650301 434637 650304
rect 434671 650301 434683 650335
rect 434625 650295 434683 650301
rect 266446 650224 266452 650276
rect 266504 650264 266510 650276
rect 270497 650267 270555 650273
rect 270497 650264 270509 650267
rect 266504 650236 270509 650264
rect 266504 650224 266510 650236
rect 270497 650233 270509 650236
rect 270543 650233 270555 650267
rect 270497 650227 270555 650233
rect 386417 650267 386475 650273
rect 386417 650233 386429 650267
rect 386463 650264 386475 650267
rect 387150 650264 387156 650276
rect 386463 650236 387156 650264
rect 386463 650233 386475 650236
rect 386417 650227 386475 650233
rect 387150 650224 387156 650236
rect 387208 650264 387214 650276
rect 389637 650267 389695 650273
rect 389637 650264 389649 650267
rect 387208 650236 389649 650264
rect 387208 650224 387214 650236
rect 389637 650233 389649 650236
rect 389683 650233 389695 650267
rect 389637 650227 389695 650233
rect 164237 650199 164295 650205
rect 164237 650165 164249 650199
rect 164283 650196 164295 650199
rect 173805 650199 173863 650205
rect 173805 650196 173817 650199
rect 164283 650168 173817 650196
rect 164283 650165 164295 650168
rect 164237 650159 164295 650165
rect 173805 650165 173817 650168
rect 173851 650165 173863 650199
rect 173805 650159 173863 650165
rect 280065 650199 280123 650205
rect 280065 650165 280077 650199
rect 280111 650196 280123 650199
rect 282270 650196 282276 650208
rect 280111 650168 282276 650196
rect 280111 650165 280123 650168
rect 280065 650159 280123 650165
rect 282270 650156 282276 650168
rect 282328 650196 282334 650208
rect 282822 650196 282828 650208
rect 282328 650168 282828 650196
rect 282328 650156 282334 650168
rect 282822 650156 282828 650168
rect 282880 650156 282886 650208
rect 405737 650199 405795 650205
rect 405737 650165 405749 650199
rect 405783 650196 405795 650199
rect 415305 650199 415363 650205
rect 415305 650196 415317 650199
rect 405783 650168 415317 650196
rect 405783 650165 405795 650168
rect 405737 650159 405795 650165
rect 415305 650165 415317 650168
rect 415351 650165 415363 650199
rect 415305 650159 415363 650165
rect 294690 645872 294696 645924
rect 294748 645912 294754 645924
rect 307386 645912 307392 645924
rect 294748 645884 307392 645912
rect 294748 645872 294754 645884
rect 307386 645872 307392 645884
rect 307444 645872 307450 645924
rect 291838 644444 291844 644496
rect 291896 644484 291902 644496
rect 307110 644484 307116 644496
rect 291896 644456 307116 644484
rect 291896 644444 291902 644456
rect 307110 644444 307116 644456
rect 307168 644444 307174 644496
rect 290458 643084 290464 643136
rect 290516 643124 290522 643136
rect 307110 643124 307116 643136
rect 290516 643096 307116 643124
rect 290516 643084 290522 643096
rect 307110 643084 307116 643096
rect 307168 643084 307174 643136
rect 287698 641724 287704 641776
rect 287756 641764 287762 641776
rect 307662 641764 307668 641776
rect 287756 641736 307668 641764
rect 287756 641724 287762 641736
rect 307662 641724 307668 641736
rect 307720 641724 307726 641776
rect 286318 640296 286324 640348
rect 286376 640336 286382 640348
rect 307662 640336 307668 640348
rect 286376 640308 307668 640336
rect 286376 640296 286382 640308
rect 307662 640296 307668 640308
rect 307720 640296 307726 640348
rect 284938 638936 284944 638988
rect 284996 638976 285002 638988
rect 306650 638976 306656 638988
rect 284996 638948 306656 638976
rect 284996 638936 285002 638948
rect 306650 638936 306656 638948
rect 306708 638936 306714 638988
rect 294598 637576 294604 637628
rect 294656 637616 294662 637628
rect 306834 637616 306840 637628
rect 294656 637588 306840 637616
rect 294656 637576 294662 637588
rect 306834 637576 306840 637588
rect 306892 637576 306898 637628
rect 389174 580252 389180 580304
rect 389232 580292 389238 580304
rect 437842 580292 437848 580304
rect 389232 580264 437848 580292
rect 389232 580252 389238 580264
rect 437842 580252 437848 580264
rect 437900 580252 437906 580304
rect 302878 579640 302884 579692
rect 302936 579680 302942 579692
rect 306926 579680 306932 579692
rect 302936 579652 306932 579680
rect 302936 579640 302942 579652
rect 306926 579640 306932 579652
rect 306984 579640 306990 579692
rect 139394 579572 139400 579624
rect 139452 579612 139458 579624
rect 187694 579612 187700 579624
rect 139452 579584 187700 579612
rect 139452 579572 139458 579584
rect 187694 579572 187700 579584
rect 187752 579572 187758 579624
rect 282178 578892 282184 578944
rect 282236 578932 282242 578944
rect 307662 578932 307668 578944
rect 282236 578904 307668 578932
rect 282236 578892 282242 578904
rect 307662 578892 307668 578904
rect 307720 578892 307726 578944
rect 302053 559011 302111 559017
rect 302053 558977 302065 559011
rect 302099 559008 302111 559011
rect 302329 559011 302387 559017
rect 302329 559008 302341 559011
rect 302099 558980 302341 559008
rect 302099 558977 302111 558980
rect 302053 558971 302111 558977
rect 302329 558977 302341 558980
rect 302375 558977 302387 559011
rect 302329 558971 302387 558977
rect 302145 558943 302203 558949
rect 302145 558909 302157 558943
rect 302191 558940 302203 558943
rect 302237 558943 302295 558949
rect 302237 558940 302249 558943
rect 302191 558912 302249 558940
rect 302191 558909 302203 558912
rect 302145 558903 302203 558909
rect 302237 558909 302249 558912
rect 302283 558909 302295 558943
rect 302237 558903 302295 558909
rect 302421 558943 302479 558949
rect 302421 558909 302433 558943
rect 302467 558940 302479 558943
rect 311805 558943 311863 558949
rect 311805 558940 311817 558943
rect 302467 558912 311817 558940
rect 302467 558909 302479 558912
rect 302421 558903 302479 558909
rect 311805 558909 311817 558912
rect 311851 558909 311863 558943
rect 311805 558903 311863 558909
rect 66162 558832 66168 558884
rect 66220 558872 66226 558884
rect 200206 558872 200212 558884
rect 66220 558844 200212 558872
rect 66220 558832 66226 558844
rect 200206 558832 200212 558844
rect 200264 558832 200270 558884
rect 220725 558875 220783 558881
rect 220725 558841 220737 558875
rect 220771 558872 220783 558875
rect 222197 558875 222255 558881
rect 222197 558872 222209 558875
rect 220771 558844 222209 558872
rect 220771 558841 220783 558844
rect 220725 558835 220783 558841
rect 222197 558841 222209 558844
rect 222243 558841 222255 558875
rect 222197 558835 222255 558841
rect 282086 558832 282092 558884
rect 282144 558872 282150 558884
rect 282144 558844 283880 558872
rect 282144 558832 282150 558844
rect 67450 558764 67456 558816
rect 67508 558804 67514 558816
rect 201494 558804 201500 558816
rect 67508 558776 201500 558804
rect 67508 558764 67514 558776
rect 201494 558764 201500 558776
rect 201552 558764 201558 558816
rect 220078 558764 220084 558816
rect 220136 558804 220142 558816
rect 229370 558804 229376 558816
rect 220136 558776 229376 558804
rect 220136 558764 220142 558776
rect 229370 558764 229376 558776
rect 229428 558804 229434 558816
rect 230753 558807 230811 558813
rect 230753 558804 230765 558807
rect 229428 558776 230765 558804
rect 229428 558764 229434 558776
rect 230753 558773 230765 558776
rect 230799 558773 230811 558807
rect 230753 558767 230811 558773
rect 79502 558696 79508 558748
rect 79560 558736 79566 558748
rect 88886 558736 88892 558748
rect 79560 558708 88892 558736
rect 79560 558696 79566 558708
rect 88886 558696 88892 558708
rect 88944 558736 88950 558748
rect 98546 558736 98552 558748
rect 88944 558708 98552 558736
rect 88944 558696 88950 558708
rect 98546 558696 98552 558708
rect 98604 558736 98610 558748
rect 101401 558739 101459 558745
rect 101401 558736 101413 558739
rect 98604 558708 101413 558736
rect 98604 558696 98610 558708
rect 101401 558705 101413 558708
rect 101447 558705 101459 558739
rect 101401 558699 101459 558705
rect 101493 558739 101551 558745
rect 101493 558705 101505 558739
rect 101539 558736 101551 558739
rect 104894 558736 104900 558748
rect 101539 558708 104900 558736
rect 101539 558705 101551 558708
rect 101493 558699 101551 558705
rect 104894 558696 104900 558708
rect 104952 558696 104958 558748
rect 125502 558696 125508 558748
rect 125560 558736 125566 558748
rect 129645 558739 129703 558745
rect 129645 558736 129657 558739
rect 125560 558708 129657 558736
rect 125560 558696 125566 558708
rect 129645 558705 129657 558708
rect 129691 558705 129703 558739
rect 129645 558699 129703 558705
rect 208486 558696 208492 558748
rect 208544 558736 208550 558748
rect 211154 558736 211160 558748
rect 208544 558708 211160 558736
rect 208544 558696 208550 558708
rect 211154 558696 211160 558708
rect 211212 558696 211218 558748
rect 217962 558696 217968 558748
rect 218020 558736 218026 558748
rect 225966 558736 225972 558748
rect 218020 558708 225972 558736
rect 218020 558696 218026 558708
rect 225966 558696 225972 558708
rect 226024 558736 226030 558748
rect 234614 558736 234620 558748
rect 226024 558708 234620 558736
rect 226024 558696 226030 558708
rect 234614 558696 234620 558708
rect 234672 558696 234678 558748
rect 78490 558628 78496 558680
rect 78548 558668 78554 558680
rect 87874 558668 87880 558680
rect 78548 558640 87880 558668
rect 78548 558628 78554 558640
rect 87874 558628 87880 558640
rect 87932 558668 87938 558680
rect 97074 558668 97080 558680
rect 87932 558640 97080 558668
rect 87932 558628 87938 558640
rect 97074 558628 97080 558640
rect 97132 558628 97138 558680
rect 97537 558671 97595 558677
rect 97537 558637 97549 558671
rect 97583 558668 97595 558671
rect 97583 558640 101720 558668
rect 97583 558637 97595 558640
rect 97537 558631 97595 558637
rect 77386 558560 77392 558612
rect 77444 558600 77450 558612
rect 86678 558600 86684 558612
rect 77444 558572 86684 558600
rect 77444 558560 77450 558572
rect 86678 558560 86684 558572
rect 86736 558560 86742 558612
rect 94866 558600 94872 558612
rect 87800 558572 94872 558600
rect 75914 558492 75920 558544
rect 75972 558532 75978 558544
rect 85390 558532 85396 558544
rect 75972 558504 85396 558532
rect 75972 558492 75978 558504
rect 85390 558492 85396 558504
rect 85448 558532 85454 558544
rect 87800 558532 87828 558572
rect 94866 558560 94872 558572
rect 94924 558600 94930 558612
rect 101692 558600 101720 558640
rect 102042 558628 102048 558680
rect 102100 558668 102106 558680
rect 140038 558668 140044 558680
rect 102100 558640 140044 558668
rect 102100 558628 102106 558640
rect 140038 558628 140044 558640
rect 140096 558628 140102 558680
rect 220722 558668 220728 558680
rect 220683 558640 220728 558668
rect 220722 558628 220728 558640
rect 220780 558628 220786 558680
rect 222197 558671 222255 558677
rect 222197 558637 222209 558671
rect 222243 558668 222255 558671
rect 227254 558668 227260 558680
rect 222243 558640 227260 558668
rect 222243 558637 222255 558640
rect 222197 558631 222255 558637
rect 227254 558628 227260 558640
rect 227312 558668 227318 558680
rect 235994 558668 236000 558680
rect 227312 558640 236000 558668
rect 227312 558628 227318 558640
rect 235994 558628 236000 558640
rect 236052 558628 236058 558680
rect 283852 558668 283880 558844
rect 283926 558832 283932 558884
rect 283984 558872 283990 558884
rect 317414 558872 317420 558884
rect 283984 558844 317420 558872
rect 283984 558832 283990 558844
rect 317414 558832 317420 558844
rect 317472 558832 317478 558884
rect 326338 558832 326344 558884
rect 326396 558872 326402 558884
rect 334161 558875 334219 558881
rect 334161 558872 334173 558875
rect 326396 558844 334173 558872
rect 326396 558832 326402 558844
rect 334161 558841 334173 558844
rect 334207 558841 334219 558875
rect 334161 558835 334219 558841
rect 334250 558832 334256 558884
rect 334308 558872 334314 558884
rect 343634 558872 343640 558884
rect 334308 558844 343640 558872
rect 334308 558832 334314 558844
rect 343634 558832 343640 558844
rect 343692 558872 343698 558884
rect 344738 558872 344744 558884
rect 343692 558844 344744 558872
rect 343692 558832 343698 558844
rect 344738 558832 344744 558844
rect 344796 558832 344802 558884
rect 344830 558832 344836 558884
rect 344888 558872 344894 558884
rect 353294 558872 353300 558884
rect 344888 558844 353300 558872
rect 344888 558832 344894 558844
rect 353294 558832 353300 558844
rect 353352 558832 353358 558884
rect 446398 558832 446404 558884
rect 446456 558872 446462 558884
rect 480530 558872 480536 558884
rect 446456 558844 480536 558872
rect 446456 558832 446462 558844
rect 480530 558832 480536 558844
rect 480588 558832 480594 558884
rect 284202 558764 284208 558816
rect 284260 558804 284266 558816
rect 320266 558804 320272 558816
rect 284260 558776 320272 558804
rect 284260 558764 284266 558776
rect 320266 558764 320272 558776
rect 320324 558764 320330 558816
rect 332502 558764 332508 558816
rect 332560 558804 332566 558816
rect 341242 558804 341248 558816
rect 332560 558776 341248 558804
rect 332560 558764 332566 558776
rect 341242 558764 341248 558776
rect 341300 558804 341306 558816
rect 350534 558804 350540 558816
rect 341300 558776 350540 558804
rect 341300 558764 341306 558776
rect 350534 558764 350540 558776
rect 350592 558764 350598 558816
rect 441614 558764 441620 558816
rect 441672 558804 441678 558816
rect 451829 558807 451887 558813
rect 451829 558804 451841 558807
rect 441672 558776 451841 558804
rect 441672 558764 441678 558776
rect 451829 558773 451841 558776
rect 451875 558773 451887 558807
rect 451829 558767 451887 558773
rect 451921 558807 451979 558813
rect 451921 558773 451933 558807
rect 451967 558804 451979 558807
rect 457346 558804 457352 558816
rect 451967 558776 457352 558804
rect 451967 558773 451979 558776
rect 451921 558767 451979 558773
rect 457346 558764 457352 558776
rect 457404 558804 457410 558816
rect 466546 558804 466552 558816
rect 457404 558776 466552 558804
rect 457404 558764 457410 558776
rect 466546 558764 466552 558776
rect 466604 558804 466610 558816
rect 475470 558804 475476 558816
rect 466604 558776 475476 558804
rect 466604 558764 466610 558776
rect 475470 558764 475476 558776
rect 475528 558764 475534 558816
rect 480257 558807 480315 558813
rect 480257 558773 480269 558807
rect 480303 558804 480315 558807
rect 483014 558804 483020 558816
rect 480303 558776 483020 558804
rect 480303 558773 480315 558776
rect 480257 558767 480315 558773
rect 483014 558764 483020 558776
rect 483072 558764 483078 558816
rect 284110 558696 284116 558748
rect 284168 558736 284174 558748
rect 320174 558736 320180 558748
rect 284168 558708 320180 558736
rect 284168 558696 284174 558708
rect 320174 558696 320180 558708
rect 320232 558696 320238 558748
rect 324958 558696 324964 558748
rect 325016 558736 325022 558748
rect 334250 558736 334256 558748
rect 325016 558708 334256 558736
rect 325016 558696 325022 558708
rect 334250 558696 334256 558708
rect 334308 558696 334314 558748
rect 336274 558696 336280 558748
rect 336332 558736 336338 558748
rect 345750 558736 345756 558748
rect 336332 558708 345756 558736
rect 336332 558696 336338 558708
rect 345750 558696 345756 558708
rect 345808 558696 345814 558748
rect 345845 558739 345903 558745
rect 345845 558705 345857 558739
rect 345891 558736 345903 558739
rect 349338 558736 349344 558748
rect 345891 558708 349344 558736
rect 345891 558705 345903 558708
rect 345845 558699 345903 558705
rect 349338 558696 349344 558708
rect 349396 558696 349402 558748
rect 443549 558739 443607 558745
rect 443549 558705 443561 558739
rect 443595 558736 443607 558739
rect 453666 558736 453672 558748
rect 443595 558708 453672 558736
rect 443595 558705 443607 558708
rect 443549 558699 443607 558705
rect 453666 558696 453672 558708
rect 453724 558736 453730 558748
rect 462590 558736 462596 558748
rect 453724 558708 462596 558736
rect 453724 558696 453730 558708
rect 462590 558696 462596 558708
rect 462648 558736 462654 558748
rect 472158 558736 472164 558748
rect 462648 558708 472164 558736
rect 462648 558696 462654 558708
rect 472158 558696 472164 558708
rect 472216 558736 472222 558748
rect 481634 558736 481640 558748
rect 472216 558708 481640 558736
rect 472216 558696 472222 558708
rect 481634 558696 481640 558708
rect 481692 558696 481698 558748
rect 302145 558671 302203 558677
rect 302145 558668 302157 558671
rect 283852 558640 302157 558668
rect 302145 558637 302157 558640
rect 302191 558637 302203 558671
rect 302145 558631 302203 558637
rect 302237 558671 302295 558677
rect 302237 558637 302249 558671
rect 302283 558668 302295 558671
rect 322842 558668 322848 558680
rect 302283 558640 322848 558668
rect 302283 558637 302295 558640
rect 302237 558631 302295 558637
rect 322842 558628 322848 558640
rect 322900 558628 322906 558680
rect 327718 558628 327724 558680
rect 327776 558668 327782 558680
rect 334161 558671 334219 558677
rect 327776 558640 334112 558668
rect 327776 558628 327782 558640
rect 102778 558600 102784 558612
rect 94924 558572 101628 558600
rect 101692 558572 102784 558600
rect 94924 558560 94930 558572
rect 95694 558532 95700 558544
rect 85448 558504 87828 558532
rect 87892 558504 95700 558532
rect 85448 558492 85454 558504
rect 80790 558424 80796 558476
rect 80848 558464 80854 558476
rect 86405 558467 86463 558473
rect 86405 558464 86417 558467
rect 80848 558436 86417 558464
rect 80848 558424 80854 558436
rect 86405 558433 86417 558436
rect 86451 558433 86463 558467
rect 86405 558427 86463 558433
rect 86678 558424 86684 558476
rect 86736 558464 86742 558476
rect 87892 558464 87920 558504
rect 95694 558492 95700 558504
rect 95752 558532 95758 558544
rect 101493 558535 101551 558541
rect 101493 558532 101505 558535
rect 95752 558504 101505 558532
rect 95752 558492 95758 558504
rect 101493 558501 101505 558504
rect 101539 558501 101551 558535
rect 101600 558532 101628 558572
rect 102778 558560 102784 558572
rect 102836 558560 102842 558612
rect 104802 558560 104808 558612
rect 104860 558600 104866 558612
rect 144178 558600 144184 558612
rect 104860 558572 144184 558600
rect 104860 558560 104866 558572
rect 144178 558560 144184 558572
rect 144236 558560 144242 558612
rect 212534 558560 212540 558612
rect 212592 558600 212598 558612
rect 213086 558600 213092 558612
rect 212592 558572 213092 558600
rect 212592 558560 212598 558572
rect 213086 558560 213092 558572
rect 213144 558600 213150 558612
rect 222286 558600 222292 558612
rect 213144 558572 222292 558600
rect 213144 558560 213150 558572
rect 222286 558560 222292 558572
rect 222344 558600 222350 558612
rect 231854 558600 231860 558612
rect 222344 558572 231860 558600
rect 222344 558560 222350 558572
rect 231854 558560 231860 558572
rect 231912 558560 231918 558612
rect 292485 558603 292543 558609
rect 292485 558569 292497 558603
rect 292531 558600 292543 558603
rect 292574 558600 292580 558612
rect 292531 558572 292580 558600
rect 292531 558569 292543 558572
rect 292485 558563 292543 558569
rect 292574 558560 292580 558572
rect 292632 558560 292638 558612
rect 311805 558603 311863 558609
rect 311805 558569 311817 558603
rect 311851 558600 311863 558603
rect 323486 558600 323492 558612
rect 311851 558572 323492 558600
rect 311851 558569 311863 558572
rect 311805 558563 311863 558569
rect 323486 558560 323492 558572
rect 323544 558600 323550 558612
rect 333146 558600 333152 558612
rect 323544 558572 333152 558600
rect 323544 558560 323550 558572
rect 333146 558560 333152 558572
rect 333204 558600 333210 558612
rect 333882 558600 333888 558612
rect 333204 558572 333888 558600
rect 333204 558560 333210 558572
rect 333882 558560 333888 558572
rect 333940 558560 333946 558612
rect 334084 558600 334112 558640
rect 334161 558637 334173 558671
rect 334207 558668 334219 558671
rect 335906 558668 335912 558680
rect 334207 558640 335912 558668
rect 334207 558637 334219 558640
rect 334161 558631 334219 558637
rect 335906 558628 335912 558640
rect 335964 558668 335970 558680
rect 344830 558668 344836 558680
rect 335964 558640 344836 558668
rect 335964 558628 335970 558640
rect 344830 558628 344836 558640
rect 344888 558628 344894 558680
rect 336274 558600 336280 558612
rect 334084 558572 336280 558600
rect 336274 558560 336280 558572
rect 336332 558560 336338 558612
rect 336734 558560 336740 558612
rect 336792 558600 336798 558612
rect 337746 558600 337752 558612
rect 336792 558572 337752 558600
rect 336792 558560 336798 558572
rect 337746 558560 337752 558572
rect 337804 558600 337810 558612
rect 345661 558603 345719 558609
rect 345661 558600 345673 558603
rect 337804 558572 345673 558600
rect 337804 558560 337810 558572
rect 345661 558569 345673 558572
rect 345707 558569 345719 558603
rect 345768 558600 345796 558696
rect 346486 558628 346492 558680
rect 346544 558668 346550 558680
rect 356054 558668 356060 558680
rect 346544 558640 356060 558668
rect 346544 558628 346550 558640
rect 356054 558628 356060 558640
rect 356112 558628 356118 558680
rect 418246 558628 418252 558680
rect 418304 558668 418310 558680
rect 432785 558671 432843 558677
rect 432785 558668 432797 558671
rect 418304 558640 432797 558668
rect 418304 558628 418310 558640
rect 432785 558637 432797 558640
rect 432831 558637 432843 558671
rect 432785 558631 432843 558637
rect 441709 558671 441767 558677
rect 441709 558637 441721 558671
rect 441755 558668 441767 558671
rect 452197 558671 452255 558677
rect 452197 558668 452209 558671
rect 441755 558640 452209 558668
rect 441755 558637 441767 558640
rect 441709 558631 441767 558637
rect 452197 558637 452209 558640
rect 452243 558637 452255 558671
rect 452197 558631 452255 558637
rect 454034 558628 454040 558680
rect 454092 558668 454098 558680
rect 454678 558668 454684 558680
rect 454092 558640 454684 558668
rect 454092 558628 454098 558640
rect 454678 558628 454684 558640
rect 454736 558668 454742 558680
rect 462501 558671 462559 558677
rect 462501 558668 462513 558671
rect 454736 558640 462513 558668
rect 454736 558628 454742 558640
rect 462501 558637 462513 558640
rect 462547 558637 462559 558671
rect 465258 558668 465264 558680
rect 462501 558631 462559 558637
rect 462884 558640 465264 558668
rect 354674 558600 354680 558612
rect 345768 558572 354680 558600
rect 345661 558563 345719 558569
rect 354674 558560 354680 558572
rect 354732 558560 354738 558612
rect 422941 558603 422999 558609
rect 422941 558569 422953 558603
rect 422987 558600 422999 558603
rect 432601 558603 432659 558609
rect 432601 558600 432613 558603
rect 422987 558572 432613 558600
rect 422987 558569 422999 558572
rect 422941 558563 422999 558569
rect 432601 558569 432613 558572
rect 432647 558569 432659 558603
rect 432601 558563 432659 558569
rect 441617 558603 441675 558609
rect 441617 558569 441629 558603
rect 441663 558600 441675 558603
rect 451921 558603 451979 558609
rect 451921 558600 451933 558603
rect 441663 558572 451933 558600
rect 441663 558569 441675 558572
rect 441617 558563 441675 558569
rect 451921 558569 451933 558572
rect 451967 558569 451979 558603
rect 451921 558563 451979 558569
rect 453301 558603 453359 558609
rect 453301 558569 453313 558603
rect 453347 558600 453359 558603
rect 455966 558600 455972 558612
rect 453347 558572 455972 558600
rect 453347 558569 453359 558572
rect 453301 558563 453359 558569
rect 455966 558560 455972 558572
rect 456024 558600 456030 558612
rect 462884 558600 462912 558640
rect 465258 558628 465264 558640
rect 465316 558668 465322 558680
rect 474826 558668 474832 558680
rect 465316 558640 474832 558668
rect 465316 558628 465322 558640
rect 474826 558628 474832 558640
rect 474884 558668 474890 558680
rect 480257 558671 480315 558677
rect 480257 558668 480269 558671
rect 474884 558640 480269 558668
rect 474884 558628 474890 558640
rect 480257 558637 480269 558640
rect 480303 558637 480315 558671
rect 480257 558631 480315 558637
rect 456024 558572 462912 558600
rect 456024 558560 456030 558572
rect 462958 558560 462964 558612
rect 463016 558600 463022 558612
rect 468662 558600 468668 558612
rect 463016 558572 468668 558600
rect 463016 558560 463022 558572
rect 468662 558560 468668 558572
rect 468720 558600 468726 558612
rect 475381 558603 475439 558609
rect 475381 558600 475393 558603
rect 468720 558572 475393 558600
rect 468720 558560 468726 558572
rect 475381 558569 475393 558572
rect 475427 558569 475439 558603
rect 475381 558563 475439 558569
rect 475470 558560 475476 558612
rect 475528 558600 475534 558612
rect 484394 558600 484400 558612
rect 475528 558572 484400 558600
rect 475528 558560 475534 558572
rect 484394 558560 484400 558572
rect 484452 558560 484458 558612
rect 104158 558532 104164 558544
rect 101600 558504 104164 558532
rect 101493 558495 101551 558501
rect 104158 558492 104164 558504
rect 104216 558492 104222 558544
rect 108482 558492 108488 558544
rect 108540 558532 108546 558544
rect 148318 558532 148324 558544
rect 108540 558504 148324 558532
rect 108540 558492 108546 558504
rect 148318 558492 148324 558504
rect 148376 558492 148382 558544
rect 218790 558492 218796 558544
rect 218848 558532 218854 558544
rect 228082 558532 228088 558544
rect 218848 558504 228088 558532
rect 218848 558492 218854 558504
rect 228082 558492 228088 558504
rect 228140 558532 228146 558544
rect 237374 558532 237380 558544
rect 228140 558504 237380 558532
rect 228140 558492 228146 558504
rect 237374 558492 237380 558504
rect 237432 558492 237438 558544
rect 284018 558492 284024 558544
rect 284076 558532 284082 558544
rect 302053 558535 302111 558541
rect 302053 558532 302065 558535
rect 284076 558504 302065 558532
rect 284076 558492 284082 558504
rect 302053 558501 302065 558504
rect 302099 558501 302111 558535
rect 302053 558495 302111 558501
rect 302142 558492 302148 558544
rect 302200 558532 302206 558544
rect 302237 558535 302295 558541
rect 302237 558532 302249 558535
rect 302200 558504 302249 558532
rect 302200 558492 302206 558504
rect 302237 558501 302249 558504
rect 302283 558501 302295 558535
rect 302237 558495 302295 558501
rect 302329 558535 302387 558541
rect 302329 558501 302341 558535
rect 302375 558532 302387 558535
rect 318794 558532 318800 558544
rect 302375 558504 318800 558532
rect 302375 558501 302387 558504
rect 302329 558495 302387 558501
rect 318794 558492 318800 558504
rect 318852 558492 318858 558544
rect 320821 558535 320879 558541
rect 320821 558501 320833 558535
rect 320867 558532 320879 558535
rect 383562 558532 383568 558544
rect 320867 558504 383568 558532
rect 320867 558501 320879 558504
rect 320821 558495 320879 558501
rect 383562 558492 383568 558504
rect 383620 558532 383626 558544
rect 443086 558532 443092 558544
rect 383620 558504 443092 558532
rect 383620 558492 383626 558504
rect 443086 558492 443092 558504
rect 443144 558492 443150 558544
rect 447137 558535 447195 558541
rect 447137 558501 447149 558535
rect 447183 558532 447195 558535
rect 451734 558532 451740 558544
rect 447183 558504 451740 558532
rect 447183 558501 447195 558504
rect 447137 558495 447195 558501
rect 451734 558492 451740 558504
rect 451792 558492 451798 558544
rect 451829 558535 451887 558541
rect 451829 558501 451841 558535
rect 451875 558532 451887 558535
rect 452289 558535 452347 558541
rect 452289 558532 452301 558535
rect 451875 558504 452301 558532
rect 451875 558501 451887 558504
rect 451829 558495 451887 558501
rect 452289 558501 452301 558504
rect 452335 558501 452347 558535
rect 452289 558495 452347 558501
rect 452378 558492 452384 558544
rect 452436 558532 452442 558544
rect 452436 558504 452792 558532
rect 452436 558492 452442 558504
rect 86736 558436 87920 558464
rect 86736 558424 86742 558436
rect 89806 558424 89812 558476
rect 89864 558464 89870 558476
rect 99374 558464 99380 558476
rect 89864 558436 99380 558464
rect 89864 558424 89870 558436
rect 99374 558424 99380 558436
rect 99432 558464 99438 558476
rect 100110 558464 100116 558476
rect 99432 558436 100116 558464
rect 99432 558424 99438 558436
rect 100110 558424 100116 558436
rect 100168 558424 100174 558476
rect 100570 558424 100576 558476
rect 100628 558464 100634 558476
rect 140130 558464 140136 558476
rect 100628 558436 140136 558464
rect 100628 558424 100634 558436
rect 140130 558424 140136 558436
rect 140188 558424 140194 558476
rect 281902 558424 281908 558476
rect 281960 558464 281966 558476
rect 329558 558464 329564 558476
rect 281960 558436 329564 558464
rect 281960 558424 281966 558436
rect 329558 558424 329564 558436
rect 329616 558464 329622 558476
rect 339034 558464 339040 558476
rect 329616 558436 339040 558464
rect 329616 558424 329622 558436
rect 339034 558424 339040 558436
rect 339092 558464 339098 558476
rect 344649 558467 344707 558473
rect 339092 558436 344600 558464
rect 339092 558424 339098 558436
rect 73706 558356 73712 558408
rect 73764 558396 73770 558408
rect 82906 558396 82912 558408
rect 73764 558368 82912 558396
rect 73764 558356 73770 558368
rect 82906 558356 82912 558368
rect 82964 558396 82970 558408
rect 86497 558399 86555 558405
rect 86497 558396 86509 558399
rect 82964 558368 86509 558396
rect 82964 558356 82970 558368
rect 86497 558365 86509 558368
rect 86543 558365 86555 558399
rect 86497 558359 86555 558365
rect 96893 558399 96951 558405
rect 96893 558365 96905 558399
rect 96939 558396 96951 558399
rect 97537 558399 97595 558405
rect 97537 558396 97549 558399
rect 96939 558368 97549 558396
rect 96939 558365 96951 558368
rect 96893 558359 96951 558365
rect 97537 558365 97549 558368
rect 97583 558365 97595 558399
rect 97537 558359 97595 558365
rect 97626 558356 97632 558408
rect 97684 558396 97690 558408
rect 138658 558396 138664 558408
rect 97684 558368 138664 558396
rect 97684 558356 97690 558368
rect 138658 558356 138664 558368
rect 138716 558356 138722 558408
rect 211154 558356 211160 558408
rect 211212 558396 211218 558408
rect 211890 558396 211896 558408
rect 211212 558368 211896 558396
rect 211212 558356 211218 558368
rect 211890 558356 211896 558368
rect 211948 558396 211954 558408
rect 221090 558396 221096 558408
rect 211948 558368 221096 558396
rect 211948 558356 211954 558368
rect 221090 558356 221096 558368
rect 221148 558396 221154 558408
rect 230474 558396 230480 558408
rect 221148 558368 230480 558396
rect 221148 558356 221154 558368
rect 230474 558356 230480 558368
rect 230532 558356 230538 558408
rect 230753 558399 230811 558405
rect 230753 558365 230765 558399
rect 230799 558396 230811 558399
rect 230799 558368 233372 558396
rect 230799 558365 230811 558368
rect 230753 558359 230811 558365
rect 81434 558288 81440 558340
rect 81492 558328 81498 558340
rect 81986 558328 81992 558340
rect 81492 558300 81992 558328
rect 81492 558288 81498 558300
rect 81986 558288 81992 558300
rect 82044 558328 82050 558340
rect 91094 558328 91100 558340
rect 82044 558300 91100 558328
rect 82044 558288 82050 558300
rect 91094 558288 91100 558300
rect 91152 558288 91158 558340
rect 92290 558288 92296 558340
rect 92348 558328 92354 558340
rect 137462 558328 137468 558340
rect 92348 558300 137468 558328
rect 92348 558288 92354 558300
rect 137462 558288 137468 558300
rect 137520 558288 137526 558340
rect 206370 558288 206376 558340
rect 206428 558328 206434 558340
rect 215294 558328 215300 558340
rect 206428 558300 215300 558328
rect 206428 558288 206434 558300
rect 215294 558288 215300 558300
rect 215352 558328 215358 558340
rect 223942 558328 223948 558340
rect 215352 558300 223948 558328
rect 215352 558288 215358 558300
rect 223942 558288 223948 558300
rect 224000 558328 224006 558340
rect 233234 558328 233240 558340
rect 224000 558300 233240 558328
rect 224000 558288 224006 558300
rect 233234 558288 233240 558300
rect 233292 558288 233298 558340
rect 233344 558328 233372 558368
rect 281994 558356 282000 558408
rect 282052 558396 282058 558408
rect 328546 558396 328552 558408
rect 282052 558368 328552 558396
rect 282052 558356 282058 558368
rect 328546 558356 328552 558368
rect 328604 558396 328610 558408
rect 336734 558396 336740 558408
rect 328604 558368 336740 558396
rect 328604 558356 328610 558368
rect 336734 558356 336740 558368
rect 336792 558356 336798 558408
rect 344572 558396 344600 558436
rect 344649 558433 344661 558467
rect 344695 558464 344707 558467
rect 345569 558467 345627 558473
rect 345569 558464 345581 558467
rect 344695 558436 345581 558464
rect 344695 558433 344707 558436
rect 344649 558427 344707 558433
rect 345569 558433 345581 558436
rect 345615 558433 345627 558467
rect 345569 558427 345627 558433
rect 345661 558467 345719 558473
rect 345661 558433 345673 558467
rect 345707 558464 345719 558467
rect 346486 558464 346492 558476
rect 345707 558436 346492 558464
rect 345707 558433 345719 558436
rect 345661 558427 345719 558433
rect 346486 558424 346492 558436
rect 346544 558424 346550 558476
rect 348234 558464 348240 558476
rect 346596 558436 348240 558464
rect 346596 558396 346624 558436
rect 348234 558424 348240 558436
rect 348292 558464 348298 558476
rect 357434 558464 357440 558476
rect 348292 558436 357440 558464
rect 348292 558424 348298 558436
rect 357434 558424 357440 558436
rect 357492 558424 357498 558476
rect 358078 558424 358084 558476
rect 358136 558464 358142 558476
rect 452654 558464 452660 558476
rect 358136 558436 452660 558464
rect 358136 558424 358142 558436
rect 452654 558424 452660 558436
rect 452712 558424 452718 558476
rect 452764 558464 452792 558504
rect 453942 558492 453948 558544
rect 454000 558532 454006 558544
rect 461670 558532 461676 558544
rect 454000 558504 461676 558532
rect 454000 558492 454006 558504
rect 461670 558492 461676 558504
rect 461728 558532 461734 558544
rect 471330 558532 471336 558544
rect 461728 558504 471336 558532
rect 461728 558492 461734 558504
rect 471330 558492 471336 558504
rect 471388 558532 471394 558544
rect 480346 558532 480352 558544
rect 471388 558504 480352 558532
rect 471388 558492 471394 558504
rect 480346 558492 480352 558504
rect 480404 558492 480410 558544
rect 456705 558467 456763 558473
rect 456705 558464 456717 558467
rect 452764 558436 456717 558464
rect 456705 558433 456717 558436
rect 456751 558433 456763 558467
rect 456705 558427 456763 558433
rect 459462 558424 459468 558476
rect 459520 558464 459526 558476
rect 468018 558464 468024 558476
rect 459520 558436 468024 558464
rect 459520 558424 459526 558436
rect 468018 558424 468024 558436
rect 468076 558464 468082 558476
rect 468754 558464 468760 558476
rect 468076 558436 468760 558464
rect 468076 558424 468082 558436
rect 468754 558424 468760 558436
rect 468812 558424 468818 558476
rect 468849 558467 468907 558473
rect 468849 558433 468861 558467
rect 468895 558464 468907 558467
rect 470042 558464 470048 558476
rect 468895 558436 470048 558464
rect 468895 558433 468907 558436
rect 468849 558427 468907 558433
rect 470042 558424 470048 558436
rect 470100 558464 470106 558476
rect 475289 558467 475347 558473
rect 475289 558464 475301 558467
rect 470100 558436 475301 558464
rect 470100 558424 470106 558436
rect 475289 558433 475301 558436
rect 475335 558433 475347 558467
rect 475289 558427 475347 558433
rect 475381 558467 475439 558473
rect 475381 558433 475393 558467
rect 475427 558464 475439 558467
rect 477586 558464 477592 558476
rect 475427 558436 477592 558464
rect 475427 558433 475439 558436
rect 475381 558427 475439 558433
rect 477586 558424 477592 558436
rect 477644 558424 477650 558476
rect 348418 558396 348424 558408
rect 344572 558368 346624 558396
rect 346688 558368 348424 558396
rect 238754 558328 238760 558340
rect 233344 558300 238760 558328
rect 238754 558288 238760 558300
rect 238812 558288 238818 558340
rect 281810 558288 281816 558340
rect 281868 558328 281874 558340
rect 330478 558328 330484 558340
rect 281868 558300 330484 558328
rect 281868 558288 281874 558300
rect 330478 558288 330484 558300
rect 330536 558328 330542 558340
rect 330536 558300 333836 558328
rect 330536 558288 330542 558300
rect 74258 558220 74264 558272
rect 74316 558260 74322 558272
rect 137370 558260 137376 558272
rect 74316 558232 137376 558260
rect 74316 558220 74322 558232
rect 137370 558220 137376 558232
rect 137428 558220 137434 558272
rect 194410 558220 194416 558272
rect 194468 558260 194474 558272
rect 231857 558263 231915 558269
rect 231857 558260 231869 558263
rect 194468 558232 231869 558260
rect 194468 558220 194474 558232
rect 231857 558229 231869 558232
rect 231903 558229 231915 558263
rect 231857 558223 231915 558229
rect 232041 558263 232099 558269
rect 232041 558229 232053 558263
rect 232087 558260 232099 558263
rect 313734 558260 313740 558272
rect 232087 558232 313740 558260
rect 232087 558229 232099 558232
rect 232041 558223 232099 558229
rect 313734 558220 313740 558232
rect 313792 558260 313798 558272
rect 320821 558263 320879 558269
rect 320821 558260 320833 558263
rect 313792 558232 320833 558260
rect 313792 558220 313798 558232
rect 320821 558229 320833 558232
rect 320867 558229 320879 558263
rect 320821 558223 320879 558229
rect 322842 558220 322848 558272
rect 322900 558260 322906 558272
rect 332502 558260 332508 558272
rect 322900 558232 332508 558260
rect 322900 558220 322906 558232
rect 332502 558220 332508 558232
rect 332560 558220 332566 558272
rect 333808 558260 333836 558300
rect 333882 558288 333888 558340
rect 333940 558328 333946 558340
rect 342530 558328 342536 558340
rect 333940 558300 342536 558328
rect 333940 558288 333946 558300
rect 342530 558288 342536 558300
rect 342588 558328 342594 558340
rect 346688 558328 346716 558368
rect 348418 558356 348424 558368
rect 348476 558356 348482 558408
rect 359458 558356 359464 558408
rect 359516 558396 359522 558408
rect 476114 558396 476120 558408
rect 359516 558368 476120 558396
rect 359516 558356 359522 558368
rect 476114 558356 476120 558368
rect 476172 558356 476178 558408
rect 476298 558356 476304 558408
rect 476356 558396 476362 558408
rect 477126 558396 477132 558408
rect 476356 558368 477132 558396
rect 476356 558356 476362 558368
rect 477126 558356 477132 558368
rect 477184 558396 477190 558408
rect 485774 558396 485780 558408
rect 477184 558368 485780 558396
rect 477184 558356 477190 558368
rect 485774 558356 485780 558368
rect 485832 558356 485838 558408
rect 342588 558300 346716 558328
rect 342588 558288 342594 558300
rect 349338 558288 349344 558340
rect 349396 558328 349402 558340
rect 357710 558328 357716 558340
rect 349396 558300 357716 558328
rect 349396 558288 349402 558300
rect 357710 558288 357716 558300
rect 357768 558288 357774 558340
rect 359550 558288 359556 558340
rect 359608 558328 359614 558340
rect 477494 558328 477500 558340
rect 359608 558300 477500 558328
rect 359608 558288 359614 558300
rect 477494 558288 477500 558300
rect 477552 558288 477558 558340
rect 339862 558260 339868 558272
rect 333808 558232 339868 558260
rect 339862 558220 339868 558232
rect 339920 558260 339926 558272
rect 344649 558263 344707 558269
rect 344649 558260 344661 558263
rect 339920 558232 344661 558260
rect 339920 558220 339926 558232
rect 344649 558229 344661 558232
rect 344695 558229 344707 558263
rect 344649 558223 344707 558229
rect 344738 558220 344744 558272
rect 344796 558260 344802 558272
rect 352006 558260 352012 558272
rect 344796 558232 352012 558260
rect 344796 558220 344802 558232
rect 352006 558220 352012 558232
rect 352064 558220 352070 558272
rect 358170 558220 358176 558272
rect 358228 558260 358234 558272
rect 476206 558260 476212 558272
rect 358228 558232 476212 558260
rect 358228 558220 358234 558232
rect 476206 558220 476212 558232
rect 476264 558220 476270 558272
rect 477586 558220 477592 558272
rect 477644 558260 477650 558272
rect 478230 558260 478236 558272
rect 477644 558232 478236 558260
rect 477644 558220 477650 558232
rect 478230 558220 478236 558232
rect 478288 558260 478294 558272
rect 487154 558260 487160 558272
rect 478288 558232 487160 558260
rect 478288 558220 478294 558232
rect 487154 558220 487160 558232
rect 487212 558220 487218 558272
rect 72510 558152 72516 558204
rect 72568 558192 72574 558204
rect 81434 558192 81440 558204
rect 72568 558164 81440 558192
rect 72568 558152 72574 558164
rect 81434 558152 81440 558164
rect 81492 558152 81498 558204
rect 83826 558152 83832 558204
rect 83884 558192 83890 558204
rect 149698 558192 149704 558204
rect 83884 558164 149704 558192
rect 83884 558152 83890 558164
rect 149698 558152 149704 558164
rect 149756 558152 149762 558204
rect 203794 558152 203800 558204
rect 203852 558192 203858 558204
rect 212534 558192 212540 558204
rect 203852 558164 212540 558192
rect 203852 558152 203858 558164
rect 212534 558152 212540 558164
rect 212592 558152 212598 558204
rect 231765 558195 231823 558201
rect 231765 558161 231777 558195
rect 231811 558192 231823 558195
rect 231946 558192 231952 558204
rect 231811 558164 231952 558192
rect 231811 558161 231823 558164
rect 231765 558155 231823 558161
rect 231946 558152 231952 558164
rect 232004 558152 232010 558204
rect 283558 558152 283564 558204
rect 283616 558192 283622 558204
rect 422941 558195 422999 558201
rect 422941 558192 422953 558195
rect 283616 558164 422953 558192
rect 283616 558152 283622 558164
rect 422941 558161 422953 558164
rect 422987 558161 422999 558195
rect 422941 558155 422999 558161
rect 432601 558195 432659 558201
rect 432601 558161 432613 558195
rect 432647 558192 432659 558195
rect 447594 558192 447600 558204
rect 432647 558164 447600 558192
rect 432647 558161 432659 558164
rect 432601 558155 432659 558161
rect 447594 558152 447600 558164
rect 447652 558152 447658 558204
rect 478874 558192 478880 558204
rect 451936 558164 478880 558192
rect 76834 558084 76840 558136
rect 76892 558124 76898 558136
rect 145558 558124 145564 558136
rect 76892 558096 145564 558124
rect 76892 558084 76898 558096
rect 145558 558084 145564 558096
rect 145616 558084 145622 558136
rect 213914 558084 213920 558136
rect 213972 558124 213978 558136
rect 222197 558127 222255 558133
rect 222197 558124 222209 558127
rect 213972 558096 222209 558124
rect 213972 558084 213978 558096
rect 222197 558093 222209 558096
rect 222243 558093 222255 558127
rect 222197 558087 222255 558093
rect 283742 558084 283748 558136
rect 283800 558124 283806 558136
rect 418246 558124 418252 558136
rect 283800 558096 418252 558124
rect 283800 558084 283806 558096
rect 418246 558084 418252 558096
rect 418304 558084 418310 558136
rect 418341 558127 418399 558133
rect 418341 558093 418353 558127
rect 418387 558124 418399 558127
rect 432693 558127 432751 558133
rect 432693 558124 432705 558127
rect 418387 558096 432705 558124
rect 418387 558093 418399 558096
rect 418341 558087 418399 558093
rect 432693 558093 432705 558096
rect 432739 558093 432751 558127
rect 432693 558087 432751 558093
rect 432785 558127 432843 558133
rect 432785 558093 432797 558127
rect 432831 558124 432843 558127
rect 449894 558124 449900 558136
rect 432831 558096 449900 558124
rect 432831 558093 432843 558096
rect 432785 558087 432843 558093
rect 449894 558084 449900 558096
rect 449952 558084 449958 558136
rect 81250 558016 81256 558068
rect 81308 558056 81314 558068
rect 152550 558056 152556 558068
rect 81308 558028 152556 558056
rect 81308 558016 81314 558028
rect 152550 558016 152556 558028
rect 152608 558016 152614 558068
rect 283834 558016 283840 558068
rect 283892 558056 283898 558068
rect 418154 558056 418160 558068
rect 283892 558028 418160 558056
rect 283892 558016 283898 558028
rect 418154 558016 418160 558028
rect 418212 558016 418218 558068
rect 418433 558059 418491 558065
rect 418433 558025 418445 558059
rect 418479 558056 418491 558059
rect 432509 558059 432567 558065
rect 432509 558056 432521 558059
rect 418479 558028 432521 558056
rect 418479 558025 418491 558028
rect 418433 558019 418491 558025
rect 432509 558025 432521 558028
rect 432555 558025 432567 558059
rect 432509 558019 432567 558025
rect 432598 558016 432604 558068
rect 432656 558056 432662 558068
rect 451274 558056 451280 558068
rect 432656 558028 451280 558056
rect 432656 558016 432662 558028
rect 451274 558016 451280 558028
rect 451332 558016 451338 558068
rect 79318 557948 79324 558000
rect 79376 557988 79382 558000
rect 152458 557988 152464 558000
rect 79376 557960 152464 557988
rect 79376 557948 79382 557960
rect 152458 557948 152464 557960
rect 152516 557948 152522 558000
rect 222197 557991 222255 557997
rect 222197 557957 222209 557991
rect 222243 557988 222255 557991
rect 223574 557988 223580 558000
rect 222243 557960 223580 557988
rect 222243 557957 222255 557960
rect 222197 557951 222255 557957
rect 223574 557948 223580 557960
rect 223632 557988 223638 558000
rect 231765 557991 231823 557997
rect 231765 557988 231777 557991
rect 223632 557960 231777 557988
rect 223632 557948 223638 557960
rect 231765 557957 231777 557960
rect 231811 557957 231823 557991
rect 231765 557951 231823 557957
rect 282270 557948 282276 558000
rect 282328 557988 282334 558000
rect 443549 557991 443607 557997
rect 443549 557988 443561 557991
rect 282328 557960 443561 557988
rect 282328 557948 282334 557960
rect 443549 557957 443561 557960
rect 443595 557957 443607 557991
rect 443549 557951 443607 557957
rect 443638 557948 443644 558000
rect 443696 557988 443702 558000
rect 451936 557988 451964 558164
rect 478874 558152 478880 558164
rect 478932 558152 478938 558204
rect 478966 558152 478972 558204
rect 479024 558192 479030 558204
rect 488534 558192 488540 558204
rect 479024 558164 488540 558192
rect 479024 558152 479030 558164
rect 488534 558152 488540 558164
rect 488592 558152 488598 558204
rect 483014 558124 483020 558136
rect 443696 557960 451964 557988
rect 452028 558096 483020 558124
rect 443696 557948 443702 557960
rect 74994 557880 75000 557932
rect 75052 557920 75058 557932
rect 84194 557920 84200 557932
rect 75052 557892 84200 557920
rect 75052 557880 75058 557892
rect 84194 557880 84200 557892
rect 84252 557880 84258 557932
rect 86405 557923 86463 557929
rect 86405 557889 86417 557923
rect 86451 557920 86463 557923
rect 89806 557920 89812 557932
rect 86451 557892 89812 557920
rect 86451 557889 86463 557892
rect 86405 557883 86463 557889
rect 89806 557880 89812 557892
rect 89864 557880 89870 557932
rect 93762 557880 93768 557932
rect 93820 557920 93826 557932
rect 137278 557920 137284 557932
rect 93820 557892 137284 557920
rect 93820 557880 93826 557892
rect 137278 557880 137284 557892
rect 137336 557880 137342 557932
rect 202138 557880 202144 557932
rect 202196 557920 202202 557932
rect 211154 557920 211160 557932
rect 202196 557892 211160 557920
rect 202196 557880 202202 557892
rect 211154 557880 211160 557892
rect 211212 557880 211218 557932
rect 282362 557880 282368 557932
rect 282420 557920 282426 557932
rect 449069 557923 449127 557929
rect 449069 557920 449081 557923
rect 282420 557892 449081 557920
rect 282420 557880 282426 557892
rect 449069 557889 449081 557892
rect 449115 557889 449127 557923
rect 449069 557883 449127 557889
rect 449158 557880 449164 557932
rect 449216 557920 449222 557932
rect 452028 557920 452056 558096
rect 483014 558084 483020 558096
rect 483072 558084 483078 558136
rect 481634 558056 481640 558068
rect 449216 557892 452056 557920
rect 452120 558028 481640 558056
rect 449216 557880 449222 557892
rect 101401 557855 101459 557861
rect 101401 557821 101413 557855
rect 101447 557852 101459 557855
rect 107654 557852 107660 557864
rect 101447 557824 107660 557852
rect 101447 557821 101459 557824
rect 101401 557815 101459 557821
rect 107654 557812 107660 557824
rect 107712 557812 107718 557864
rect 122745 557855 122803 557861
rect 122745 557821 122757 557855
rect 122791 557852 122803 557855
rect 125137 557855 125195 557861
rect 125137 557852 125149 557855
rect 122791 557824 125149 557852
rect 122791 557821 122803 557824
rect 122745 557815 122803 557821
rect 125137 557821 125149 557824
rect 125183 557821 125195 557855
rect 125137 557815 125195 557821
rect 129645 557855 129703 557861
rect 129645 557821 129657 557855
rect 129691 557852 129703 557855
rect 208486 557852 208492 557864
rect 129691 557824 208492 557852
rect 129691 557821 129703 557824
rect 129645 557815 129703 557821
rect 208486 557812 208492 557824
rect 208544 557812 208550 557864
rect 282454 557812 282460 557864
rect 282512 557852 282518 557864
rect 282512 557824 447640 557852
rect 282512 557812 282518 557824
rect 89346 557744 89352 557796
rect 89404 557784 89410 557796
rect 96985 557787 97043 557793
rect 96985 557784 96997 557787
rect 89404 557756 96997 557784
rect 89404 557744 89410 557756
rect 96985 557753 96997 557756
rect 97031 557753 97043 557787
rect 96985 557747 97043 557753
rect 97074 557744 97080 557796
rect 97132 557784 97138 557796
rect 106274 557784 106280 557796
rect 97132 557756 106280 557784
rect 97132 557744 97138 557756
rect 106274 557744 106280 557756
rect 106332 557744 106338 557796
rect 121362 557744 121368 557796
rect 121420 557784 121426 557796
rect 206370 557784 206376 557796
rect 121420 557756 206376 557784
rect 121420 557744 121426 557756
rect 206370 557744 206376 557756
rect 206428 557744 206434 557796
rect 207658 557744 207664 557796
rect 207716 557784 207722 557796
rect 217962 557784 217968 557796
rect 207716 557756 217968 557784
rect 207716 557744 207722 557756
rect 217962 557744 217968 557756
rect 218020 557744 218026 557796
rect 282546 557744 282552 557796
rect 282604 557784 282610 557796
rect 418157 557787 418215 557793
rect 418157 557784 418169 557787
rect 282604 557756 418169 557784
rect 282604 557744 282610 557756
rect 418157 557753 418169 557756
rect 418203 557753 418215 557787
rect 418157 557747 418215 557753
rect 418433 557787 418491 557793
rect 418433 557753 418445 557787
rect 418479 557784 418491 557787
rect 432601 557787 432659 557793
rect 432601 557784 432613 557787
rect 418479 557756 432613 557784
rect 418479 557753 418491 557756
rect 418433 557747 418491 557753
rect 432601 557753 432613 557756
rect 432647 557753 432659 557787
rect 432601 557747 432659 557753
rect 432693 557787 432751 557793
rect 432693 557753 432705 557787
rect 432739 557784 432751 557787
rect 441617 557787 441675 557793
rect 441617 557784 441629 557787
rect 432739 557756 441629 557784
rect 432739 557753 432751 557756
rect 432693 557747 432751 557753
rect 441617 557753 441629 557756
rect 441663 557753 441675 557787
rect 441617 557747 441675 557753
rect 91094 557676 91100 557728
rect 91152 557716 91158 557728
rect 100018 557716 100024 557728
rect 91152 557688 100024 557716
rect 91152 557676 91158 557688
rect 100018 557676 100024 557688
rect 100076 557676 100082 557728
rect 100110 557676 100116 557728
rect 100168 557716 100174 557728
rect 108298 557716 108304 557728
rect 100168 557688 108304 557716
rect 100168 557676 100174 557688
rect 108298 557676 108304 557688
rect 108356 557676 108362 557728
rect 117222 557676 117228 557728
rect 117280 557716 117286 557728
rect 203794 557716 203800 557728
rect 117280 557688 203800 557716
rect 117280 557676 117286 557688
rect 203794 557676 203800 557688
rect 203852 557676 203858 557728
rect 204898 557676 204904 557728
rect 204956 557716 204962 557728
rect 213914 557716 213920 557728
rect 204956 557688 213920 557716
rect 204956 557676 204962 557688
rect 213914 557676 213920 557688
rect 213972 557676 213978 557728
rect 282638 557676 282644 557728
rect 282696 557716 282702 557728
rect 418249 557719 418307 557725
rect 418249 557716 418261 557719
rect 282696 557688 418261 557716
rect 282696 557676 282702 557688
rect 418249 557685 418261 557688
rect 418295 557685 418307 557719
rect 418249 557679 418307 557685
rect 432509 557719 432567 557725
rect 432509 557685 432521 557719
rect 432555 557716 432567 557719
rect 441709 557719 441767 557725
rect 441709 557716 441721 557719
rect 432555 557688 441721 557716
rect 432555 557685 432567 557688
rect 432509 557679 432567 557685
rect 441709 557685 441721 557688
rect 441755 557685 441767 557719
rect 441709 557679 441767 557685
rect 86497 557651 86555 557657
rect 86497 557617 86509 557651
rect 86543 557648 86555 557651
rect 92474 557648 92480 557660
rect 86543 557620 92480 557648
rect 86543 557617 86555 557620
rect 86497 557611 86555 557617
rect 92474 557608 92480 557620
rect 92532 557648 92538 557660
rect 100846 557648 100852 557660
rect 92532 557620 100852 557648
rect 92532 557608 92538 557620
rect 100846 557608 100852 557620
rect 100904 557608 100910 557660
rect 122745 557651 122803 557657
rect 122745 557648 122757 557651
rect 102612 557620 122757 557648
rect 84194 557540 84200 557592
rect 84252 557580 84258 557592
rect 93578 557580 93584 557592
rect 84252 557552 93584 557580
rect 84252 557540 84258 557552
rect 93578 557540 93584 557552
rect 93636 557580 93642 557592
rect 96893 557583 96951 557589
rect 96893 557580 96905 557583
rect 93636 557552 96905 557580
rect 93636 557540 93642 557552
rect 96893 557549 96905 557552
rect 96939 557549 96951 557583
rect 96893 557543 96951 557549
rect 96985 557583 97043 557589
rect 96985 557549 96997 557583
rect 97031 557580 97043 557583
rect 102612 557580 102640 557620
rect 122745 557617 122757 557620
rect 122791 557617 122803 557651
rect 122745 557611 122803 557617
rect 125137 557651 125195 557657
rect 125137 557617 125149 557651
rect 125183 557648 125195 557651
rect 125183 557620 129596 557648
rect 125183 557617 125195 557620
rect 125137 557611 125195 557617
rect 97031 557552 102640 557580
rect 97031 557549 97043 557552
rect 96985 557543 97043 557549
rect 107470 557540 107476 557592
rect 107528 557580 107534 557592
rect 129461 557583 129519 557589
rect 129461 557580 129473 557583
rect 107528 557552 129473 557580
rect 107528 557540 107534 557552
rect 129461 557549 129473 557552
rect 129507 557549 129519 557583
rect 129461 557543 129519 557549
rect 129568 557512 129596 557620
rect 129734 557608 129740 557660
rect 129792 557648 129798 557660
rect 210510 557648 210516 557660
rect 129792 557620 210516 557648
rect 129792 557608 129798 557620
rect 210510 557608 210516 557620
rect 210568 557648 210574 557660
rect 220078 557648 220084 557660
rect 210568 557620 220084 557648
rect 210568 557608 210574 557620
rect 220078 557608 220084 557620
rect 220136 557608 220142 557660
rect 282730 557608 282736 557660
rect 282788 557648 282794 557660
rect 447137 557651 447195 557657
rect 447137 557648 447149 557651
rect 282788 557620 447149 557648
rect 282788 557608 282794 557620
rect 447137 557617 447149 557620
rect 447183 557617 447195 557651
rect 447612 557648 447640 557824
rect 447778 557812 447784 557864
rect 447836 557852 447842 557864
rect 452120 557852 452148 558028
rect 481634 558016 481640 558028
rect 481692 558016 481698 558068
rect 452197 557991 452255 557997
rect 452197 557957 452209 557991
rect 452243 557988 452255 557991
rect 458266 557988 458272 558000
rect 452243 557960 458272 557988
rect 452243 557957 452255 557960
rect 452197 557951 452255 557957
rect 458266 557948 458272 557960
rect 458324 557988 458330 558000
rect 459462 557988 459468 558000
rect 458324 557960 459468 557988
rect 458324 557948 458330 557960
rect 459462 557948 459468 557960
rect 459520 557948 459526 558000
rect 460842 557948 460848 558000
rect 460900 557988 460906 558000
rect 468665 557991 468723 557997
rect 468665 557988 468677 557991
rect 460900 557960 468677 557988
rect 460900 557948 460906 557960
rect 468665 557957 468677 557960
rect 468711 557957 468723 557991
rect 468665 557951 468723 557957
rect 468754 557948 468760 558000
rect 468812 557988 468818 558000
rect 475197 557991 475255 557997
rect 475197 557988 475209 557991
rect 468812 557960 475209 557988
rect 468812 557948 468818 557960
rect 475197 557957 475209 557960
rect 475243 557957 475255 557991
rect 475197 557951 475255 557957
rect 475289 557991 475347 557997
rect 475289 557957 475301 557991
rect 475335 557988 475347 557991
rect 478966 557988 478972 558000
rect 475335 557960 478972 557988
rect 475335 557957 475347 557960
rect 475289 557951 475347 557957
rect 478966 557948 478972 557960
rect 479024 557948 479030 558000
rect 454678 557880 454684 557932
rect 454736 557920 454742 557932
rect 458177 557923 458235 557929
rect 458177 557920 458189 557923
rect 454736 557892 458189 557920
rect 454736 557880 454742 557892
rect 458177 557889 458189 557892
rect 458223 557889 458235 557923
rect 460860 557920 460888 557948
rect 458177 557883 458235 557889
rect 458284 557892 460888 557920
rect 447836 557824 452148 557852
rect 452289 557855 452347 557861
rect 447836 557812 447842 557824
rect 452289 557821 452301 557855
rect 452335 557852 452347 557855
rect 458284 557852 458312 557892
rect 464338 557880 464344 557932
rect 464396 557920 464402 557932
rect 488534 557920 488540 557932
rect 464396 557892 488540 557920
rect 464396 557880 464402 557892
rect 488534 557880 488540 557892
rect 488592 557880 488598 557932
rect 452335 557824 458312 557852
rect 458361 557855 458419 557861
rect 452335 557821 452347 557824
rect 452289 557815 452347 557821
rect 458361 557821 458373 557855
rect 458407 557852 458419 557855
rect 487154 557852 487160 557864
rect 458407 557824 487160 557852
rect 458407 557821 458419 557824
rect 458361 557815 458419 557821
rect 487154 557812 487160 557824
rect 487212 557812 487218 557864
rect 451918 557744 451924 557796
rect 451976 557784 451982 557796
rect 484394 557784 484400 557796
rect 451976 557756 484400 557784
rect 451976 557744 451982 557756
rect 484394 557744 484400 557756
rect 484452 557744 484458 557796
rect 450538 557676 450544 557728
rect 450596 557716 450602 557728
rect 483106 557716 483112 557728
rect 450596 557688 483112 557716
rect 450596 557676 450602 557688
rect 483106 557676 483112 557688
rect 483164 557676 483170 557728
rect 453301 557651 453359 557657
rect 453301 557648 453313 557651
rect 447612 557620 453313 557648
rect 447137 557611 447195 557617
rect 453301 557617 453313 557620
rect 453347 557617 453359 557651
rect 453301 557611 453359 557617
rect 453482 557608 453488 557660
rect 453540 557648 453546 557660
rect 485774 557648 485780 557660
rect 453540 557620 485780 557648
rect 453540 557608 453546 557620
rect 485774 557608 485780 557620
rect 485832 557608 485838 557660
rect 129829 557583 129887 557589
rect 129829 557549 129841 557583
rect 129875 557580 129887 557583
rect 141418 557580 141424 557592
rect 129875 557552 141424 557580
rect 129875 557549 129887 557552
rect 129829 557543 129887 557549
rect 141418 557540 141424 557552
rect 141476 557540 141482 557592
rect 209038 557540 209044 557592
rect 209096 557580 209102 557592
rect 218790 557580 218796 557592
rect 209096 557552 218796 557580
rect 209096 557540 209102 557552
rect 218790 557540 218796 557552
rect 218848 557540 218854 557592
rect 282822 557540 282828 557592
rect 282880 557580 282886 557592
rect 418249 557583 418307 557589
rect 418249 557580 418261 557583
rect 282880 557552 418261 557580
rect 282880 557540 282886 557552
rect 418249 557549 418261 557552
rect 418295 557549 418307 557583
rect 418249 557543 418307 557549
rect 418338 557540 418344 557592
rect 418396 557580 418402 557592
rect 432506 557580 432512 557592
rect 418396 557552 432512 557580
rect 418396 557540 418402 557552
rect 432506 557540 432512 557552
rect 432564 557540 432570 557592
rect 432601 557583 432659 557589
rect 432601 557549 432613 557583
rect 432647 557580 432659 557583
rect 441614 557580 441620 557592
rect 432647 557552 441620 557580
rect 432647 557549 432659 557552
rect 432601 557543 432659 557549
rect 441614 557540 441620 557552
rect 441672 557540 441678 557592
rect 449069 557583 449127 557589
rect 449069 557549 449081 557583
rect 449115 557580 449127 557583
rect 454034 557580 454040 557592
rect 449115 557552 454040 557580
rect 449115 557549 449127 557552
rect 449069 557543 449127 557549
rect 454034 557540 454040 557552
rect 454092 557540 454098 557592
rect 456705 557583 456763 557589
rect 456705 557549 456717 557583
rect 456751 557580 456763 557583
rect 459646 557580 459652 557592
rect 456751 557552 459652 557580
rect 456751 557549 456763 557552
rect 456705 557543 456763 557549
rect 459646 557540 459652 557552
rect 459704 557540 459710 557592
rect 462501 557583 462559 557589
rect 462501 557549 462513 557583
rect 462547 557580 462559 557583
rect 464246 557580 464252 557592
rect 462547 557552 464252 557580
rect 462547 557549 462559 557552
rect 462501 557543 462559 557549
rect 464246 557540 464252 557552
rect 464304 557580 464310 557592
rect 473446 557580 473452 557592
rect 464304 557552 473452 557580
rect 464304 557540 464310 557552
rect 473446 557540 473452 557552
rect 473504 557580 473510 557592
rect 474642 557580 474648 557592
rect 473504 557552 474648 557580
rect 473504 557540 473510 557552
rect 474642 557540 474648 557552
rect 474700 557540 474706 557592
rect 475197 557583 475255 557589
rect 475197 557549 475209 557583
rect 475243 557580 475255 557583
rect 476298 557580 476304 557592
rect 475243 557552 476304 557580
rect 475243 557549 475255 557552
rect 475197 557543 475255 557549
rect 476298 557540 476304 557552
rect 476356 557540 476362 557592
rect 476390 557540 476396 557592
rect 476448 557580 476454 557592
rect 483014 557580 483020 557592
rect 476448 557552 483020 557580
rect 476448 557540 476454 557552
rect 483014 557540 483020 557552
rect 483072 557540 483078 557592
rect 131758 557512 131764 557524
rect 129568 557484 131764 557512
rect 131758 557472 131764 557484
rect 131816 557472 131822 557524
rect 283466 557472 283472 557524
rect 283524 557512 283530 557524
rect 292485 557515 292543 557521
rect 292485 557512 292497 557515
rect 283524 557484 292497 557512
rect 283524 557472 283530 557484
rect 292485 557481 292497 557484
rect 292531 557481 292543 557515
rect 292485 557475 292543 557481
rect 96522 545028 96528 545080
rect 96580 545068 96586 545080
rect 189626 545068 189632 545080
rect 96580 545040 189632 545068
rect 96580 545028 96586 545040
rect 189626 545028 189632 545040
rect 189684 545028 189690 545080
rect 94130 544960 94136 545012
rect 94188 545000 94194 545012
rect 188430 545000 188436 545012
rect 94188 544972 188436 545000
rect 94188 544960 94194 544972
rect 188430 544960 188436 544972
rect 188488 544960 188494 545012
rect 102042 544892 102048 544944
rect 102100 544932 102106 544944
rect 197906 544932 197912 544944
rect 102100 544904 197912 544932
rect 102100 544892 102106 544904
rect 197906 544892 197912 544904
rect 197964 544892 197970 544944
rect 92106 544824 92112 544876
rect 92164 544864 92170 544876
rect 188522 544864 188528 544876
rect 92164 544836 188528 544864
rect 92164 544824 92170 544836
rect 188522 544824 188528 544836
rect 188580 544824 188586 544876
rect 89990 544756 89996 544808
rect 90048 544796 90054 544808
rect 188614 544796 188620 544808
rect 90048 544768 188620 544796
rect 90048 544756 90054 544768
rect 188614 544756 188620 544768
rect 188672 544756 188678 544808
rect 106182 544688 106188 544740
rect 106240 544728 106246 544740
rect 206186 544728 206192 544740
rect 106240 544700 206192 544728
rect 106240 544688 106246 544700
rect 206186 544688 206192 544700
rect 206244 544688 206250 544740
rect 87966 544620 87972 544672
rect 88024 544660 88030 544672
rect 188706 544660 188712 544672
rect 88024 544632 188712 544660
rect 88024 544620 88030 544632
rect 188706 544620 188712 544632
rect 188764 544620 188770 544672
rect 110322 544552 110328 544604
rect 110380 544592 110386 544604
rect 212442 544592 212448 544604
rect 110380 544564 212448 544592
rect 110380 544552 110386 544564
rect 212442 544552 212448 544564
rect 212500 544552 212506 544604
rect 85850 544484 85856 544536
rect 85908 544524 85914 544536
rect 188798 544524 188804 544536
rect 85908 544496 188804 544524
rect 85908 544484 85914 544496
rect 188798 544484 188804 544496
rect 188856 544484 188862 544536
rect 83826 544416 83832 544468
rect 83884 544456 83890 544468
rect 188890 544456 188896 544468
rect 83884 544428 188896 544456
rect 83884 544416 83890 544428
rect 188890 544416 188896 544428
rect 188948 544416 188954 544468
rect 81710 544348 81716 544400
rect 81768 544388 81774 544400
rect 195974 544388 195980 544400
rect 81768 544360 195980 544388
rect 81768 544348 81774 544360
rect 195974 544348 195980 544360
rect 196032 544348 196038 544400
rect 86770 544280 86776 544332
rect 86828 544320 86834 544332
rect 173066 544320 173072 544332
rect 86828 544292 173072 544320
rect 86828 544280 86834 544292
rect 173066 544280 173072 544292
rect 173124 544280 173130 544332
rect 88242 544212 88248 544264
rect 88300 544252 88306 544264
rect 175090 544252 175096 544264
rect 88300 544224 175096 544252
rect 88300 544212 88306 544224
rect 175090 544212 175096 544224
rect 175148 544212 175154 544264
rect 86862 544144 86868 544196
rect 86920 544184 86926 544196
rect 170950 544184 170956 544196
rect 86920 544156 170956 544184
rect 86920 544144 86926 544156
rect 170950 544144 170956 544156
rect 171008 544144 171014 544196
rect 85482 544076 85488 544128
rect 85540 544116 85546 544128
rect 168834 544116 168840 544128
rect 85540 544088 168840 544116
rect 85540 544076 85546 544088
rect 168834 544076 168840 544088
rect 168892 544076 168898 544128
rect 82722 544008 82728 544060
rect 82780 544048 82786 544060
rect 164694 544048 164700 544060
rect 82780 544020 164700 544048
rect 82780 544008 82786 544020
rect 164694 544008 164700 544020
rect 164752 544008 164758 544060
rect 73062 543940 73068 543992
rect 73120 543980 73126 543992
rect 148134 543980 148140 543992
rect 73120 543952 148140 543980
rect 73120 543940 73126 543952
rect 148134 543940 148140 543952
rect 148192 543940 148198 543992
rect 57882 543872 57888 543924
rect 57940 543912 57946 543924
rect 112806 543912 112812 543924
rect 57940 543884 112812 543912
rect 57940 543872 57946 543884
rect 112806 543872 112812 543884
rect 112864 543872 112870 543924
rect 57790 543804 57796 543856
rect 57848 543844 57854 543856
rect 110782 543844 110788 543856
rect 57848 543816 110788 543844
rect 57848 543804 57854 543816
rect 110782 543804 110788 543816
rect 110840 543804 110846 543856
rect 220722 543736 220728 543788
rect 220780 543736 220786 543788
rect 71682 543668 71688 543720
rect 71740 543708 71746 543720
rect 75454 543708 75460 543720
rect 71740 543680 75460 543708
rect 71740 543668 71746 543680
rect 75454 543668 75460 543680
rect 75512 543668 75518 543720
rect 75822 543668 75828 543720
rect 75880 543708 75886 543720
rect 145469 543711 145527 543717
rect 145469 543708 145481 543711
rect 75880 543680 145481 543708
rect 75880 543668 75886 543680
rect 145469 543677 145481 543680
rect 145515 543677 145527 543711
rect 145469 543671 145527 543677
rect 145558 543668 145564 543720
rect 145616 543708 145622 543720
rect 152461 543711 152519 543717
rect 152461 543708 152473 543711
rect 145616 543680 152473 543708
rect 145616 543668 145622 543680
rect 152461 543677 152473 543680
rect 152507 543677 152519 543711
rect 152461 543671 152519 543677
rect 152550 543668 152556 543720
rect 152608 543708 152614 543720
rect 162670 543708 162676 543720
rect 152608 543680 162676 543708
rect 152608 543668 152614 543680
rect 162670 543668 162676 543680
rect 162728 543668 162734 543720
rect 205542 543668 205548 543720
rect 205600 543708 205606 543720
rect 218698 543708 218704 543720
rect 205600 543680 218704 543708
rect 205600 543668 205606 543680
rect 218698 543668 218704 543680
rect 218756 543668 218762 543720
rect 220538 543668 220544 543720
rect 220596 543708 220602 543720
rect 220740 543708 220768 543736
rect 220596 543680 220768 543708
rect 220596 543668 220602 543680
rect 227622 543668 227628 543720
rect 227680 543708 227686 543720
rect 258074 543708 258080 543720
rect 227680 543680 258080 543708
rect 227680 543668 227686 543680
rect 258074 543668 258080 543680
rect 258132 543668 258138 543720
rect 78582 543600 78588 543652
rect 78640 543640 78646 543652
rect 156414 543640 156420 543652
rect 78640 543612 156420 543640
rect 78640 543600 78646 543612
rect 156414 543600 156420 543612
rect 156472 543600 156478 543652
rect 206922 543600 206928 543652
rect 206980 543640 206986 543652
rect 220722 543640 220728 543652
rect 206980 543612 220728 543640
rect 206980 543600 206986 543612
rect 220722 543600 220728 543612
rect 220780 543600 220786 543652
rect 229002 543600 229008 543652
rect 229060 543640 229066 543652
rect 260190 543640 260196 543652
rect 229060 543612 260196 543640
rect 229060 543600 229066 543612
rect 260190 543600 260196 543612
rect 260248 543600 260254 543652
rect 61010 543532 61016 543584
rect 61068 543572 61074 543584
rect 62022 543572 62028 543584
rect 61068 543544 62028 543572
rect 61068 543532 61074 543544
rect 62022 543532 62028 543544
rect 62080 543532 62086 543584
rect 65150 543532 65156 543584
rect 65208 543572 65214 543584
rect 66162 543572 66168 543584
rect 65208 543544 66168 543572
rect 65208 543532 65214 543544
rect 66162 543532 66168 543544
rect 66220 543532 66226 543584
rect 70302 543532 70308 543584
rect 70360 543572 70366 543584
rect 71314 543572 71320 543584
rect 70360 543544 71320 543572
rect 70360 543532 70366 543544
rect 71314 543532 71320 543544
rect 71372 543532 71378 543584
rect 79962 543532 79968 543584
rect 80020 543572 80026 543584
rect 152369 543575 152427 543581
rect 152369 543572 152381 543575
rect 80020 543544 152381 543572
rect 80020 543532 80026 543544
rect 152369 543541 152381 543544
rect 152415 543541 152427 543575
rect 152369 543535 152427 543541
rect 152458 543532 152464 543584
rect 152516 543572 152522 543584
rect 158530 543572 158536 543584
rect 152516 543544 158536 543572
rect 152516 543532 152522 543544
rect 158530 543532 158536 543544
rect 158588 543532 158594 543584
rect 208302 543532 208308 543584
rect 208360 543572 208366 543584
rect 222838 543572 222844 543584
rect 208360 543544 222844 543572
rect 208360 543532 208366 543544
rect 222838 543532 222844 543544
rect 222896 543532 222902 543584
rect 230382 543532 230388 543584
rect 230440 543572 230446 543584
rect 262214 543572 262220 543584
rect 230440 543544 262220 543572
rect 230440 543532 230446 543544
rect 262214 543532 262220 543544
rect 262272 543532 262278 543584
rect 57422 543464 57428 543516
rect 57480 543504 57486 543516
rect 102502 543504 102508 543516
rect 57480 543476 102508 543504
rect 57480 543464 57486 543476
rect 102502 543464 102508 543476
rect 102560 543464 102566 543516
rect 127342 543464 127348 543516
rect 127400 543504 127406 543516
rect 209038 543504 209044 543516
rect 127400 543476 209044 543504
rect 127400 543464 127406 543476
rect 209038 543464 209044 543476
rect 209096 543464 209102 543516
rect 209682 543464 209688 543516
rect 209740 543504 209746 543516
rect 224862 543504 224868 543516
rect 209740 543476 224868 543504
rect 209740 543464 209746 543476
rect 224862 543464 224868 543476
rect 224920 543464 224926 543516
rect 231762 543464 231768 543516
rect 231820 543504 231826 543516
rect 264330 543504 264336 543516
rect 231820 543476 264336 543504
rect 231820 543464 231826 543476
rect 264330 543464 264336 543476
rect 264388 543464 264394 543516
rect 57514 543396 57520 543448
rect 57572 543436 57578 543448
rect 104526 543436 104532 543448
rect 57572 543408 104532 543436
rect 57572 543396 57578 543408
rect 104526 543396 104532 543408
rect 104584 543396 104590 543448
rect 123202 543396 123208 543448
rect 123260 543436 123266 543448
rect 207658 543436 207664 543448
rect 123260 543408 207664 543436
rect 123260 543396 123266 543408
rect 207658 543396 207664 543408
rect 207716 543396 207722 543448
rect 210970 543396 210976 543448
rect 211028 543436 211034 543448
rect 226978 543436 226984 543448
rect 211028 543408 226984 543436
rect 211028 543396 211034 543408
rect 226978 543396 226984 543408
rect 227036 543396 227042 543448
rect 233142 543396 233148 543448
rect 233200 543436 233206 543448
rect 266446 543436 266452 543448
rect 233200 543408 266452 543436
rect 233200 543396 233206 543408
rect 266446 543396 266452 543408
rect 266504 543396 266510 543448
rect 57606 543328 57612 543380
rect 57664 543368 57670 543380
rect 106642 543368 106648 543380
rect 57664 543340 106648 543368
rect 57664 543328 57670 543340
rect 106642 543328 106648 543340
rect 106700 543328 106706 543380
rect 119062 543328 119068 543380
rect 119120 543368 119126 543380
rect 204898 543368 204904 543380
rect 119120 543340 204904 543368
rect 119120 543328 119126 543340
rect 204898 543328 204904 543340
rect 204956 543328 204962 543380
rect 212350 543328 212356 543380
rect 212408 543368 212414 543380
rect 231118 543368 231124 543380
rect 212408 543340 231124 543368
rect 212408 543328 212414 543340
rect 231118 543328 231124 543340
rect 231176 543328 231182 543380
rect 233050 543328 233056 543380
rect 233108 543368 233114 543380
rect 268470 543368 268476 543380
rect 233108 543340 268476 543368
rect 233108 543328 233114 543340
rect 268470 543328 268476 543340
rect 268528 543328 268534 543380
rect 91002 543260 91008 543312
rect 91060 543300 91066 543312
rect 179230 543300 179236 543312
rect 91060 543272 179236 543300
rect 91060 543260 91066 543272
rect 179230 543260 179236 543272
rect 179288 543260 179294 543312
rect 215202 543260 215208 543312
rect 215260 543300 215266 543312
rect 235258 543300 235264 543312
rect 215260 543272 235264 543300
rect 215260 543260 215266 543272
rect 235258 543260 235264 543272
rect 235316 543260 235322 543312
rect 235902 543260 235908 543312
rect 235960 543300 235966 543312
rect 272610 543300 272616 543312
rect 235960 543272 272616 543300
rect 235960 543260 235966 543272
rect 272610 543260 272616 543272
rect 272668 543260 272674 543312
rect 57698 543192 57704 543244
rect 57756 543232 57762 543244
rect 108666 543232 108672 543244
rect 57756 543204 108672 543232
rect 57756 543192 57762 543204
rect 108666 543192 108672 543204
rect 108724 543192 108730 543244
rect 114922 543192 114928 543244
rect 114980 543232 114986 543244
rect 202138 543232 202144 543244
rect 114980 543204 202144 543232
rect 114980 543192 114986 543204
rect 202138 543192 202144 543204
rect 202196 543192 202202 543244
rect 211062 543192 211068 543244
rect 211120 543232 211126 543244
rect 229094 543232 229100 543244
rect 211120 543204 229100 543232
rect 211120 543192 211126 543204
rect 229094 543192 229100 543204
rect 229152 543192 229158 543244
rect 234522 543192 234528 543244
rect 234580 543232 234586 543244
rect 270586 543232 270592 543244
rect 234580 543204 270592 543232
rect 234580 543192 234586 543204
rect 270586 543192 270592 543204
rect 270644 543192 270650 543244
rect 93670 543124 93676 543176
rect 93728 543164 93734 543176
rect 183370 543164 183376 543176
rect 93728 543136 183376 543164
rect 93728 543124 93734 543136
rect 183370 543124 183376 543136
rect 183428 543124 183434 543176
rect 202782 543124 202788 543176
rect 202840 543164 202846 543176
rect 214558 543164 214564 543176
rect 202840 543136 214564 543164
rect 202840 543124 202846 543136
rect 214558 543124 214564 543136
rect 214616 543124 214622 543176
rect 216582 543124 216588 543176
rect 216640 543164 216646 543176
rect 237374 543164 237380 543176
rect 216640 543136 237380 543164
rect 216640 543124 216646 543136
rect 237374 543124 237380 543136
rect 237432 543124 237438 543176
rect 238662 543124 238668 543176
rect 238720 543164 238726 543176
rect 276750 543164 276756 543176
rect 238720 543136 276756 543164
rect 238720 543124 238726 543136
rect 276750 543124 276756 543136
rect 276808 543124 276814 543176
rect 57238 543056 57244 543108
rect 57296 543096 57302 543108
rect 79686 543096 79692 543108
rect 57296 543068 79692 543096
rect 57296 543056 57302 543068
rect 79686 543056 79692 543068
rect 79744 543056 79750 543108
rect 95050 543056 95056 543108
rect 95108 543096 95114 543108
rect 187510 543096 187516 543108
rect 95108 543068 187516 543096
rect 95108 543056 95114 543068
rect 187510 543056 187516 543068
rect 187568 543056 187574 543108
rect 204162 543056 204168 543108
rect 204220 543056 204226 543108
rect 213822 543056 213828 543108
rect 213880 543096 213886 543108
rect 233234 543096 233240 543108
rect 213880 543068 233240 543096
rect 213880 543056 213886 543068
rect 233234 543056 233240 543068
rect 233292 543056 233298 543108
rect 237282 543056 237288 543108
rect 237340 543096 237346 543108
rect 274726 543096 274732 543108
rect 237340 543068 274732 543096
rect 237340 543056 237346 543068
rect 274726 543056 274732 543068
rect 274784 543056 274790 543108
rect 67542 542988 67548 543040
rect 67600 543028 67606 543040
rect 98362 543028 98368 543040
rect 67600 543000 98368 543028
rect 67600 542988 67606 543000
rect 98362 542988 98368 543000
rect 98420 542988 98426 543040
rect 99282 542988 99288 543040
rect 99340 543028 99346 543040
rect 193766 543028 193772 543040
rect 99340 543000 193772 543028
rect 99340 542988 99346 543000
rect 193766 542988 193772 543000
rect 193824 542988 193830 543040
rect 204180 543028 204208 543056
rect 216582 543028 216588 543040
rect 204180 543000 216588 543028
rect 216582 542988 216588 543000
rect 216640 542988 216646 543040
rect 217870 542988 217876 543040
rect 217928 543028 217934 543040
rect 239398 543028 239404 543040
rect 217928 543000 239404 543028
rect 217928 542988 217934 543000
rect 239398 542988 239404 543000
rect 239456 542988 239462 543040
rect 240042 542988 240048 543040
rect 240100 543028 240106 543040
rect 278866 543028 278872 543040
rect 240100 543000 278872 543028
rect 240100 542988 240106 543000
rect 278866 542988 278872 543000
rect 278924 542988 278930 543040
rect 57330 542920 57336 542972
rect 57388 542960 57394 542972
rect 100386 542960 100392 542972
rect 57388 542932 100392 542960
rect 57388 542920 57394 542932
rect 100386 542920 100392 542932
rect 100444 542920 100450 542972
rect 108574 542920 108580 542972
rect 108632 542960 108638 542972
rect 143994 542960 144000 542972
rect 108632 542932 144000 542960
rect 108632 542920 108638 542932
rect 143994 542920 144000 542932
rect 144052 542920 144058 542972
rect 144178 542920 144184 542972
rect 144236 542960 144242 542972
rect 204162 542960 204168 542972
rect 144236 542932 204168 542960
rect 144236 542920 144242 542932
rect 204162 542920 204168 542932
rect 204220 542920 204226 542972
rect 226150 542920 226156 542972
rect 226208 542960 226214 542972
rect 256050 542960 256056 542972
rect 226208 542932 256056 542960
rect 226208 542920 226214 542932
rect 256050 542920 256056 542932
rect 256108 542920 256114 542972
rect 105538 542852 105544 542904
rect 105596 542892 105602 542904
rect 139854 542892 139860 542904
rect 105596 542864 139860 542892
rect 105596 542852 105602 542864
rect 139854 542852 139860 542864
rect 139912 542852 139918 542904
rect 140130 542852 140136 542904
rect 140188 542892 140194 542904
rect 195882 542892 195888 542904
rect 140188 542864 195888 542892
rect 140188 542852 140194 542864
rect 195882 542852 195888 542864
rect 195940 542852 195946 542904
rect 226242 542852 226248 542904
rect 226300 542892 226306 542904
rect 253934 542892 253940 542904
rect 226300 542864 253940 542892
rect 226300 542852 226306 542864
rect 253934 542852 253940 542864
rect 253992 542852 253998 542904
rect 104158 542784 104164 542836
rect 104216 542824 104222 542836
rect 137738 542824 137744 542836
rect 104216 542796 137744 542824
rect 104216 542784 104222 542796
rect 137738 542784 137744 542796
rect 137796 542784 137802 542836
rect 138658 542784 138664 542836
rect 138716 542824 138722 542836
rect 191742 542824 191748 542836
rect 138716 542796 191748 542824
rect 138716 542784 138722 542796
rect 191742 542784 191748 542796
rect 191800 542784 191806 542836
rect 223482 542784 223488 542836
rect 223540 542824 223546 542836
rect 249794 542824 249800 542836
rect 223540 542796 249800 542824
rect 223540 542784 223546 542796
rect 249794 542784 249800 542796
rect 249852 542784 249858 542836
rect 102778 542716 102784 542768
rect 102836 542756 102842 542768
rect 135714 542756 135720 542768
rect 102836 542728 135720 542756
rect 102836 542716 102842 542728
rect 135714 542716 135720 542728
rect 135772 542716 135778 542768
rect 137278 542716 137284 542768
rect 137336 542756 137342 542768
rect 185486 542756 185492 542768
rect 137336 542728 185492 542756
rect 137336 542716 137342 542728
rect 185486 542716 185492 542728
rect 185544 542716 185550 542768
rect 224678 542716 224684 542768
rect 224736 542756 224742 542768
rect 251910 542756 251916 542768
rect 224736 542728 251916 542756
rect 224736 542716 224742 542728
rect 251910 542716 251916 542728
rect 251968 542716 251974 542768
rect 70210 542648 70216 542700
rect 70268 542688 70274 542700
rect 73430 542688 73436 542700
rect 70268 542660 73436 542688
rect 70268 542648 70274 542660
rect 73430 542648 73436 542660
rect 73488 542648 73494 542700
rect 100018 542648 100024 542700
rect 100076 542688 100082 542700
rect 131482 542688 131488 542700
rect 100076 542660 131488 542688
rect 100076 542648 100082 542660
rect 131482 542648 131488 542660
rect 131540 542648 131546 542700
rect 131758 542648 131764 542700
rect 131816 542688 131822 542700
rect 177206 542688 177212 542700
rect 131816 542660 177212 542688
rect 131816 542648 131822 542660
rect 177206 542648 177212 542660
rect 177264 542648 177270 542700
rect 222102 542648 222108 542700
rect 222160 542688 222166 542700
rect 247770 542688 247776 542700
rect 222160 542660 247776 542688
rect 222160 542648 222166 542660
rect 247770 542648 247776 542660
rect 247828 542648 247834 542700
rect 101398 542580 101404 542632
rect 101456 542620 101462 542632
rect 133598 542620 133604 542632
rect 101456 542592 133604 542620
rect 101456 542580 101462 542592
rect 133598 542580 133604 542592
rect 133656 542580 133662 542632
rect 137462 542580 137468 542632
rect 137520 542620 137526 542632
rect 181346 542620 181352 542632
rect 137520 542592 181352 542620
rect 137520 542580 137526 542592
rect 181346 542580 181352 542592
rect 181404 542580 181410 542632
rect 220538 542580 220544 542632
rect 220596 542620 220602 542632
rect 245654 542620 245660 542632
rect 220596 542592 245660 542620
rect 220596 542580 220602 542592
rect 245654 542580 245660 542592
rect 245712 542580 245718 542632
rect 108298 542512 108304 542564
rect 108356 542552 108362 542564
rect 146018 542552 146024 542564
rect 108356 542524 146024 542552
rect 108356 542512 108362 542524
rect 146018 542512 146024 542524
rect 146076 542512 146082 542564
rect 152274 542552 152280 542564
rect 146956 542524 152280 542552
rect 106918 542444 106924 542496
rect 106976 542484 106982 542496
rect 141878 542484 141884 542496
rect 106976 542456 141884 542484
rect 106976 542444 106982 542456
rect 141878 542444 141884 542456
rect 141936 542444 141942 542496
rect 145469 542487 145527 542493
rect 145469 542453 145481 542487
rect 145515 542484 145527 542487
rect 146956 542484 146984 542524
rect 152274 542512 152280 542524
rect 152332 542512 152338 542564
rect 152461 542555 152519 542561
rect 152461 542521 152473 542555
rect 152507 542552 152519 542555
rect 154390 542552 154396 542564
rect 152507 542524 154396 542552
rect 152507 542521 152519 542524
rect 152461 542515 152519 542521
rect 154390 542512 154396 542524
rect 154448 542512 154454 542564
rect 166810 542552 166816 542564
rect 156616 542524 166816 542552
rect 145515 542456 146984 542484
rect 145515 542453 145527 542456
rect 145469 542447 145527 542453
rect 149698 542444 149704 542496
rect 149756 542484 149762 542496
rect 156616 542484 156644 542524
rect 166810 542512 166816 542524
rect 166868 542512 166874 542564
rect 217962 542512 217968 542564
rect 218020 542552 218026 542564
rect 241514 542552 241520 542564
rect 218020 542524 241520 542552
rect 218020 542512 218026 542524
rect 241514 542512 241520 542524
rect 241572 542512 241578 542564
rect 149756 542456 156644 542484
rect 149756 542444 149762 542456
rect 219342 542444 219348 542496
rect 219400 542484 219406 542496
rect 243538 542484 243544 542496
rect 219400 542456 243544 542484
rect 219400 542444 219406 542456
rect 243538 542444 243544 542456
rect 243596 542444 243602 542496
rect 137370 542376 137376 542428
rect 137428 542416 137434 542428
rect 150158 542416 150164 542428
rect 137428 542388 150164 542416
rect 137428 542376 137434 542388
rect 150158 542376 150164 542388
rect 150216 542376 150222 542428
rect 152369 542419 152427 542425
rect 152369 542385 152381 542419
rect 152415 542416 152427 542419
rect 160554 542416 160560 542428
rect 152415 542388 160560 542416
rect 152415 542385 152427 542388
rect 152369 542379 152427 542385
rect 160554 542376 160560 542388
rect 160612 542376 160618 542428
rect 281718 539520 281724 539572
rect 281776 539560 281782 539572
rect 464338 539560 464344 539572
rect 281776 539532 464344 539560
rect 281776 539520 281782 539532
rect 464338 539520 464344 539532
rect 464396 539520 464402 539572
rect 281718 538160 281724 538212
rect 281776 538200 281782 538212
rect 454678 538200 454684 538212
rect 281776 538172 454684 538200
rect 281776 538160 281782 538172
rect 454678 538160 454684 538172
rect 454736 538160 454742 538212
rect 281718 535372 281724 535424
rect 281776 535412 281782 535424
rect 453482 535412 453488 535424
rect 281776 535384 453488 535412
rect 281776 535372 281782 535384
rect 453482 535372 453488 535384
rect 453540 535372 453546 535424
rect 281718 534012 281724 534064
rect 281776 534052 281782 534064
rect 451918 534052 451924 534064
rect 281776 534024 451924 534052
rect 281776 534012 281782 534024
rect 451918 534012 451924 534024
rect 451976 534012 451982 534064
rect 281718 531224 281724 531276
rect 281776 531264 281782 531276
rect 450538 531264 450544 531276
rect 281776 531236 450544 531264
rect 281776 531224 281782 531236
rect 450538 531224 450544 531236
rect 450596 531224 450602 531276
rect 281718 529864 281724 529916
rect 281776 529904 281782 529916
rect 449158 529904 449164 529916
rect 281776 529876 449164 529904
rect 281776 529864 281782 529876
rect 449158 529864 449164 529876
rect 449216 529864 449222 529916
rect 281718 527076 281724 527128
rect 281776 527116 281782 527128
rect 447778 527116 447784 527128
rect 281776 527088 447784 527116
rect 281776 527076 281782 527088
rect 447778 527076 447784 527088
rect 447836 527076 447842 527128
rect 281718 525716 281724 525768
rect 281776 525756 281782 525768
rect 446398 525756 446404 525768
rect 281776 525728 446404 525756
rect 281776 525716 281782 525728
rect 446398 525716 446404 525728
rect 446456 525716 446462 525768
rect 281718 522928 281724 522980
rect 281776 522968 281782 522980
rect 443638 522968 443644 522980
rect 281776 522940 443644 522968
rect 281776 522928 281782 522940
rect 443638 522928 443644 522940
rect 443696 522928 443702 522980
rect 281718 521568 281724 521620
rect 281776 521608 281782 521620
rect 359550 521608 359556 521620
rect 281776 521580 359556 521608
rect 281776 521568 281782 521580
rect 359550 521568 359556 521580
rect 359608 521568 359614 521620
rect 281718 518848 281724 518900
rect 281776 518888 281782 518900
rect 359458 518888 359464 518900
rect 281776 518860 359464 518888
rect 281776 518848 281782 518860
rect 359458 518848 359464 518860
rect 359516 518848 359522 518900
rect 281718 517420 281724 517472
rect 281776 517460 281782 517472
rect 358170 517460 358176 517472
rect 281776 517432 358176 517460
rect 281776 517420 281782 517432
rect 358170 517420 358176 517432
rect 358228 517420 358234 517472
rect 281718 514700 281724 514752
rect 281776 514740 281782 514752
rect 356698 514740 356704 514752
rect 281776 514712 356704 514740
rect 281776 514700 281782 514712
rect 356698 514700 356704 514712
rect 356756 514700 356762 514752
rect 281718 513272 281724 513324
rect 281776 513312 281782 513324
rect 473354 513312 473360 513324
rect 281776 513284 473360 513312
rect 281776 513272 281782 513284
rect 473354 513272 473360 513284
rect 473412 513272 473418 513324
rect 281718 510552 281724 510604
rect 281776 510592 281782 510604
rect 471974 510592 471980 510604
rect 281776 510564 471980 510592
rect 281776 510552 281782 510564
rect 471974 510552 471980 510564
rect 472032 510552 472038 510604
rect 281718 509192 281724 509244
rect 281776 509232 281782 509244
rect 470594 509232 470600 509244
rect 281776 509204 470600 509232
rect 281776 509192 281782 509204
rect 470594 509192 470600 509204
rect 470652 509192 470658 509244
rect 281718 506404 281724 506456
rect 281776 506444 281782 506456
rect 469214 506444 469220 506456
rect 281776 506416 469220 506444
rect 281776 506404 281782 506416
rect 469214 506404 469220 506416
rect 469272 506404 469278 506456
rect 281718 505044 281724 505096
rect 281776 505084 281782 505096
rect 467926 505084 467932 505096
rect 281776 505056 467932 505084
rect 281776 505044 281782 505056
rect 467926 505044 467932 505056
rect 467984 505044 467990 505096
rect 281718 502256 281724 502308
rect 281776 502296 281782 502308
rect 467834 502296 467840 502308
rect 281776 502268 467840 502296
rect 281776 502256 281782 502268
rect 467834 502256 467840 502268
rect 467892 502256 467898 502308
rect 281718 500896 281724 500948
rect 281776 500936 281782 500948
rect 466454 500936 466460 500948
rect 281776 500908 466460 500936
rect 281776 500896 281782 500908
rect 466454 500896 466460 500908
rect 466512 500896 466518 500948
rect 281718 499468 281724 499520
rect 281776 499508 281782 499520
rect 465074 499508 465080 499520
rect 281776 499480 465080 499508
rect 281776 499468 281782 499480
rect 465074 499468 465080 499480
rect 465132 499468 465138 499520
rect 281718 496748 281724 496800
rect 281776 496788 281782 496800
rect 463694 496788 463700 496800
rect 281776 496760 463700 496788
rect 281776 496748 281782 496760
rect 463694 496748 463700 496760
rect 463752 496748 463758 496800
rect 281718 495388 281724 495440
rect 281776 495428 281782 495440
rect 462314 495428 462320 495440
rect 281776 495400 462320 495428
rect 281776 495388 281782 495400
rect 462314 495388 462320 495400
rect 462372 495388 462378 495440
rect 281718 492600 281724 492652
rect 281776 492640 281782 492652
rect 461026 492640 461032 492652
rect 281776 492612 461032 492640
rect 281776 492600 281782 492612
rect 461026 492600 461032 492612
rect 461084 492600 461090 492652
rect 281718 491240 281724 491292
rect 281776 491280 281782 491292
rect 460934 491280 460940 491292
rect 281776 491252 460940 491280
rect 281776 491240 281782 491252
rect 460934 491240 460940 491252
rect 460992 491240 460998 491292
rect 281718 488452 281724 488504
rect 281776 488492 281782 488504
rect 459554 488492 459560 488504
rect 281776 488464 459560 488492
rect 281776 488452 281782 488464
rect 459554 488452 459560 488464
rect 459612 488452 459618 488504
rect 281718 487092 281724 487144
rect 281776 487132 281782 487144
rect 458174 487132 458180 487144
rect 281776 487104 458180 487132
rect 281776 487092 281782 487104
rect 458174 487092 458180 487104
rect 458232 487092 458238 487144
rect 281718 484304 281724 484356
rect 281776 484344 281782 484356
rect 456794 484344 456800 484356
rect 281776 484316 456800 484344
rect 281776 484304 281782 484316
rect 456794 484304 456800 484316
rect 456852 484304 456858 484356
rect 281718 482944 281724 482996
rect 281776 482984 281782 482996
rect 455414 482984 455420 482996
rect 281776 482956 455420 482984
rect 281776 482944 281782 482956
rect 455414 482944 455420 482956
rect 455472 482944 455478 482996
rect 281718 480156 281724 480208
rect 281776 480196 281782 480208
rect 453390 480196 453396 480208
rect 281776 480168 453396 480196
rect 281776 480156 281782 480168
rect 453390 480156 453396 480168
rect 453448 480156 453454 480208
rect 281718 478796 281724 478848
rect 281776 478836 281782 478848
rect 358078 478836 358084 478848
rect 281776 478808 358084 478836
rect 281776 478796 281782 478808
rect 358078 478796 358084 478808
rect 358136 478796 358142 478848
rect 281718 476008 281724 476060
rect 281776 476048 281782 476060
rect 452654 476048 452660 476060
rect 281776 476020 452660 476048
rect 281776 476008 281782 476020
rect 452654 476008 452660 476020
rect 452712 476008 452718 476060
rect 281718 474648 281724 474700
rect 281776 474688 281782 474700
rect 358906 474688 358912 474700
rect 281776 474660 358912 474688
rect 281776 474648 281782 474660
rect 358906 474648 358912 474660
rect 358964 474648 358970 474700
rect 281718 471928 281724 471980
rect 281776 471968 281782 471980
rect 357526 471968 357532 471980
rect 281776 471940 357532 471968
rect 281776 471928 281782 471940
rect 357526 471928 357532 471940
rect 357584 471928 357590 471980
rect 281718 470500 281724 470552
rect 281776 470540 281782 470552
rect 356054 470540 356060 470552
rect 281776 470512 356060 470540
rect 281776 470500 281782 470512
rect 356054 470500 356060 470512
rect 356112 470500 356118 470552
rect 281718 467780 281724 467832
rect 281776 467820 281782 467832
rect 354674 467820 354680 467832
rect 281776 467792 354680 467820
rect 281776 467780 281782 467792
rect 354674 467780 354680 467792
rect 354732 467780 354738 467832
rect 281718 466352 281724 466404
rect 281776 466392 281782 466404
rect 353294 466392 353300 466404
rect 281776 466364 353300 466392
rect 281776 466352 281782 466364
rect 353294 466352 353300 466364
rect 353352 466352 353358 466404
rect 281718 463632 281724 463684
rect 281776 463672 281782 463684
rect 352006 463672 352012 463684
rect 281776 463644 352012 463672
rect 281776 463632 281782 463644
rect 352006 463632 352012 463644
rect 352064 463632 352070 463684
rect 281718 462272 281724 462324
rect 281776 462312 281782 462324
rect 352190 462312 352196 462324
rect 281776 462284 352196 462312
rect 281776 462272 281782 462284
rect 352190 462272 352196 462284
rect 352248 462272 352254 462324
rect 281718 459484 281724 459536
rect 281776 459524 281782 459536
rect 350534 459524 350540 459536
rect 281776 459496 350540 459524
rect 281776 459484 281782 459496
rect 350534 459484 350540 459496
rect 350592 459484 350598 459536
rect 281718 458124 281724 458176
rect 281776 458164 281782 458176
rect 349154 458164 349160 458176
rect 281776 458136 349160 458164
rect 281776 458124 281782 458136
rect 349154 458124 349160 458136
rect 349212 458124 349218 458176
rect 281718 455336 281724 455388
rect 281776 455376 281782 455388
rect 347774 455376 347780 455388
rect 281776 455348 347780 455376
rect 281776 455336 281782 455348
rect 347774 455336 347780 455348
rect 347832 455336 347838 455388
rect 281718 453976 281724 454028
rect 281776 454016 281782 454028
rect 346394 454016 346400 454028
rect 281776 453988 346400 454016
rect 281776 453976 281782 453988
rect 346394 453976 346400 453988
rect 346452 453976 346458 454028
rect 281718 452548 281724 452600
rect 281776 452588 281782 452600
rect 345014 452588 345020 452600
rect 281776 452560 345020 452588
rect 281776 452548 281782 452560
rect 345014 452548 345020 452560
rect 345072 452548 345078 452600
rect 281718 449828 281724 449880
rect 281776 449868 281782 449880
rect 343726 449868 343732 449880
rect 281776 449840 343732 449868
rect 281776 449828 281782 449840
rect 343726 449828 343732 449840
rect 343784 449828 343790 449880
rect 281718 448468 281724 448520
rect 281776 448508 281782 448520
rect 343634 448508 343640 448520
rect 281776 448480 343640 448508
rect 281776 448468 281782 448480
rect 343634 448468 343640 448480
rect 343692 448468 343698 448520
rect 281718 445680 281724 445732
rect 281776 445720 281782 445732
rect 342254 445720 342260 445732
rect 281776 445692 342260 445720
rect 281776 445680 281782 445692
rect 342254 445680 342260 445692
rect 342312 445680 342318 445732
rect 281718 444320 281724 444372
rect 281776 444360 281782 444372
rect 340874 444360 340880 444372
rect 281776 444332 340880 444360
rect 281776 444320 281782 444332
rect 340874 444320 340880 444332
rect 340932 444320 340938 444372
rect 281718 441532 281724 441584
rect 281776 441572 281782 441584
rect 339494 441572 339500 441584
rect 281776 441544 339500 441572
rect 281776 441532 281782 441544
rect 339494 441532 339500 441544
rect 339552 441532 339558 441584
rect 281718 440172 281724 440224
rect 281776 440212 281782 440224
rect 338114 440212 338120 440224
rect 281776 440184 338120 440212
rect 281776 440172 281782 440184
rect 338114 440172 338120 440184
rect 338172 440172 338178 440224
rect 281718 437384 281724 437436
rect 281776 437424 281782 437436
rect 336826 437424 336832 437436
rect 281776 437396 336832 437424
rect 281776 437384 281782 437396
rect 336826 437384 336832 437396
rect 336884 437384 336890 437436
rect 281718 436024 281724 436076
rect 281776 436064 281782 436076
rect 336734 436064 336740 436076
rect 281776 436036 336740 436064
rect 281776 436024 281782 436036
rect 336734 436024 336740 436036
rect 336792 436024 336798 436076
rect 281718 433236 281724 433288
rect 281776 433276 281782 433288
rect 335354 433276 335360 433288
rect 281776 433248 335360 433276
rect 281776 433236 281782 433248
rect 335354 433236 335360 433248
rect 335412 433236 335418 433288
rect 281718 431876 281724 431928
rect 281776 431916 281782 431928
rect 333974 431916 333980 431928
rect 281776 431888 333980 431916
rect 281776 431876 281782 431888
rect 333974 431876 333980 431888
rect 334032 431876 334038 431928
rect 281718 429088 281724 429140
rect 281776 429128 281782 429140
rect 332594 429128 332600 429140
rect 281776 429100 332600 429128
rect 281776 429088 281782 429100
rect 332594 429088 332600 429100
rect 332652 429088 332658 429140
rect 281718 427728 281724 427780
rect 281776 427768 281782 427780
rect 331214 427768 331220 427780
rect 281776 427740 331220 427768
rect 281776 427728 281782 427740
rect 331214 427728 331220 427740
rect 331272 427728 331278 427780
rect 281718 425008 281724 425060
rect 281776 425048 281782 425060
rect 329926 425048 329932 425060
rect 281776 425020 329932 425048
rect 281776 425008 281782 425020
rect 329926 425008 329932 425020
rect 329984 425008 329990 425060
rect 281718 423580 281724 423632
rect 281776 423620 281782 423632
rect 329834 423620 329840 423632
rect 281776 423592 329840 423620
rect 281776 423580 281782 423592
rect 329834 423580 329840 423592
rect 329892 423580 329898 423632
rect 281718 420860 281724 420912
rect 281776 420900 281782 420912
rect 328454 420900 328460 420912
rect 281776 420872 328460 420900
rect 281776 420860 281782 420872
rect 328454 420860 328460 420872
rect 328512 420860 328518 420912
rect 281718 419432 281724 419484
rect 281776 419472 281782 419484
rect 327074 419472 327080 419484
rect 281776 419444 327080 419472
rect 281776 419432 281782 419444
rect 327074 419432 327080 419444
rect 327132 419432 327138 419484
rect 281718 418072 281724 418124
rect 281776 418112 281782 418124
rect 325694 418112 325700 418124
rect 281776 418084 325700 418112
rect 281776 418072 281782 418084
rect 325694 418072 325700 418084
rect 325752 418072 325758 418124
rect 281718 415352 281724 415404
rect 281776 415392 281782 415404
rect 324314 415392 324320 415404
rect 281776 415364 324320 415392
rect 281776 415352 281782 415364
rect 324314 415352 324320 415364
rect 324372 415352 324378 415404
rect 281718 413924 281724 413976
rect 281776 413964 281782 413976
rect 322934 413964 322940 413976
rect 281776 413936 322940 413964
rect 281776 413924 281782 413936
rect 322934 413924 322940 413936
rect 322992 413924 322998 413976
rect 383562 413244 383568 413296
rect 383620 413284 383626 413296
rect 404998 413284 405004 413296
rect 383620 413256 405004 413284
rect 383620 413244 383626 413256
rect 404998 413244 405004 413256
rect 405056 413244 405062 413296
rect 404998 412632 405004 412684
rect 405056 412672 405062 412684
rect 513374 412672 513380 412684
rect 405056 412644 513380 412672
rect 405056 412632 405062 412644
rect 513374 412632 513380 412644
rect 513432 412632 513438 412684
rect 285306 412428 285312 412480
rect 285364 412468 285370 412480
rect 316034 412468 316040 412480
rect 285364 412440 316040 412468
rect 285364 412428 285370 412440
rect 316034 412428 316040 412440
rect 316092 412428 316098 412480
rect 281626 412360 281632 412412
rect 281684 412400 281690 412412
rect 324958 412400 324964 412412
rect 281684 412372 324964 412400
rect 281684 412360 281690 412372
rect 324958 412360 324964 412372
rect 325016 412360 325022 412412
rect 281534 412292 281540 412344
rect 281592 412332 281598 412344
rect 326338 412332 326344 412344
rect 281592 412304 326344 412332
rect 281592 412292 281598 412304
rect 326338 412292 326344 412304
rect 326396 412292 326402 412344
rect 281997 412267 282055 412273
rect 281997 412233 282009 412267
rect 282043 412264 282055 412267
rect 327718 412264 327724 412276
rect 282043 412236 327724 412264
rect 282043 412233 282055 412236
rect 281997 412227 282055 412233
rect 327718 412224 327724 412236
rect 327776 412224 327782 412276
rect 283098 412156 283104 412208
rect 283156 412196 283162 412208
rect 438578 412196 438584 412208
rect 283156 412168 438584 412196
rect 283156 412156 283162 412168
rect 438578 412156 438584 412168
rect 438636 412156 438642 412208
rect 283006 412088 283012 412140
rect 283064 412128 283070 412140
rect 438486 412128 438492 412140
rect 283064 412100 438492 412128
rect 283064 412088 283070 412100
rect 438486 412088 438492 412100
rect 438544 412088 438550 412140
rect 283190 412020 283196 412072
rect 283248 412060 283254 412072
rect 438670 412060 438676 412072
rect 283248 412032 438676 412060
rect 283248 412020 283254 412032
rect 438670 412020 438676 412032
rect 438728 412020 438734 412072
rect 283282 411952 283288 412004
rect 283340 411992 283346 412004
rect 445754 411992 445760 412004
rect 283340 411964 445760 411992
rect 283340 411952 283346 411964
rect 445754 411952 445760 411964
rect 445812 411952 445818 412004
rect 285398 411884 285404 411936
rect 285456 411924 285462 411936
rect 453298 411924 453304 411936
rect 285456 411896 453304 411924
rect 285456 411884 285462 411896
rect 453298 411884 453304 411896
rect 453356 411884 453362 411936
rect 281718 411340 281724 411392
rect 281776 411380 281782 411392
rect 281994 411380 282000 411392
rect 281776 411352 282000 411380
rect 281776 411340 281782 411352
rect 281994 411340 282000 411352
rect 282052 411340 282058 411392
rect 281994 411204 282000 411256
rect 282052 411244 282058 411256
rect 321554 411244 321560 411256
rect 282052 411216 321560 411244
rect 282052 411204 282058 411216
rect 321554 411204 321560 411216
rect 321612 411204 321618 411256
rect 285214 410796 285220 410848
rect 285272 410836 285278 410848
rect 438118 410836 438124 410848
rect 285272 410808 438124 410836
rect 285272 410796 285278 410808
rect 438118 410796 438124 410808
rect 438176 410796 438182 410848
rect 285122 410728 285128 410780
rect 285180 410768 285186 410780
rect 438210 410768 438216 410780
rect 285180 410740 438216 410768
rect 285180 410728 285186 410740
rect 438210 410728 438216 410740
rect 438268 410728 438274 410780
rect 285030 410660 285036 410712
rect 285088 410700 285094 410712
rect 438302 410700 438308 410712
rect 285088 410672 438308 410700
rect 285088 410660 285094 410672
rect 438302 410660 438308 410672
rect 438360 410660 438366 410712
rect 283374 410592 283380 410644
rect 283432 410632 283438 410644
rect 438762 410632 438768 410644
rect 283432 410604 438768 410632
rect 283432 410592 283438 410604
rect 438762 410592 438768 410604
rect 438820 410592 438826 410644
rect 281994 410564 282000 410576
rect 281955 410536 282000 410564
rect 281994 410524 282000 410536
rect 282052 410524 282058 410576
rect 282914 410524 282920 410576
rect 282972 410564 282978 410576
rect 438394 410564 438400 410576
rect 282972 410536 438400 410564
rect 282972 410524 282978 410536
rect 438394 410524 438400 410536
rect 438452 410524 438458 410576
rect 281534 404132 281540 404184
rect 281592 404172 281598 404184
rect 281994 404172 282000 404184
rect 281592 404144 282000 404172
rect 281592 404132 281598 404144
rect 281994 404132 282000 404144
rect 282052 404132 282058 404184
rect 281534 397060 281540 397112
rect 281592 397100 281598 397112
rect 283466 397100 283472 397112
rect 281592 397072 283472 397100
rect 281592 397060 281598 397072
rect 283466 397060 283472 397072
rect 283524 397060 283530 397112
rect 281902 378020 281908 378072
rect 281960 378060 281966 378072
rect 285398 378060 285404 378072
rect 281960 378032 285404 378060
rect 281960 378020 281966 378032
rect 285398 378020 285404 378032
rect 285456 378020 285462 378072
rect 282822 376660 282828 376712
rect 282880 376700 282886 376712
rect 294690 376700 294696 376712
rect 282880 376672 294696 376700
rect 282880 376660 282886 376672
rect 294690 376660 294696 376672
rect 294748 376660 294754 376712
rect 282822 373940 282828 373992
rect 282880 373980 282886 373992
rect 291838 373980 291844 373992
rect 282880 373952 291844 373980
rect 282880 373940 282886 373952
rect 291838 373940 291844 373952
rect 291896 373940 291902 373992
rect 282822 372512 282828 372564
rect 282880 372552 282886 372564
rect 290458 372552 290464 372564
rect 282880 372524 290464 372552
rect 282880 372512 282886 372524
rect 290458 372512 290464 372524
rect 290516 372512 290522 372564
rect 282362 371016 282368 371068
rect 282420 371056 282426 371068
rect 287698 371056 287704 371068
rect 282420 371028 287704 371056
rect 282420 371016 282426 371028
rect 287698 371016 287704 371028
rect 287756 371016 287762 371068
rect 282270 368024 282276 368076
rect 282328 368064 282334 368076
rect 286318 368064 286324 368076
rect 282328 368036 286324 368064
rect 282328 368024 282334 368036
rect 286318 368024 286324 368036
rect 286376 368024 286382 368076
rect 281718 365780 281724 365832
rect 281776 365820 281782 365832
rect 284938 365820 284944 365832
rect 281776 365792 284944 365820
rect 281776 365780 281782 365792
rect 284938 365780 284944 365792
rect 284996 365780 285002 365832
rect 282822 364284 282828 364336
rect 282880 364324 282886 364336
rect 294598 364324 294604 364336
rect 282880 364296 294604 364324
rect 282880 364284 282886 364296
rect 294598 364284 294604 364296
rect 294656 364284 294662 364336
rect 281902 362856 281908 362908
rect 281960 362896 281966 362908
rect 285306 362896 285312 362908
rect 281960 362868 285312 362896
rect 281960 362856 281966 362868
rect 285306 362856 285312 362868
rect 285364 362856 285370 362908
rect 281902 360136 281908 360188
rect 281960 360176 281966 360188
rect 285214 360176 285220 360188
rect 281960 360148 285220 360176
rect 281960 360136 281966 360148
rect 285214 360136 285220 360148
rect 285272 360136 285278 360188
rect 281718 357620 281724 357672
rect 281776 357660 281782 357672
rect 285122 357660 285128 357672
rect 281776 357632 285128 357660
rect 281776 357620 281782 357632
rect 285122 357620 285128 357632
rect 285180 357620 285186 357672
rect 282086 355852 282092 355904
rect 282144 355892 282150 355904
rect 285030 355892 285036 355904
rect 282144 355864 285036 355892
rect 282144 355852 282150 355864
rect 285030 355852 285036 355864
rect 285088 355852 285094 355904
rect 281534 346060 281540 346112
rect 281592 346100 281598 346112
rect 283282 346100 283288 346112
rect 281592 346072 283288 346100
rect 281592 346060 281598 346072
rect 283282 346060 283288 346072
rect 283340 346060 283346 346112
rect 282822 343544 282828 343596
rect 282880 343584 282886 343596
rect 302878 343584 302884 343596
rect 282880 343556 302884 343584
rect 282880 343544 282886 343556
rect 302878 343544 302884 343556
rect 302936 343544 302942 343596
rect 281534 341300 281540 341352
rect 281592 341340 281598 341352
rect 283374 341340 283380 341352
rect 281592 341312 283380 341340
rect 281592 341300 281598 341312
rect 283374 341300 283380 341312
rect 283432 341300 283438 341352
rect 281718 339260 281724 339312
rect 281776 339300 281782 339312
rect 284202 339300 284208 339312
rect 281776 339272 284208 339300
rect 281776 339260 281782 339272
rect 284202 339260 284208 339272
rect 284260 339260 284266 339312
rect 281534 337560 281540 337612
rect 281592 337600 281598 337612
rect 284110 337600 284116 337612
rect 281592 337572 284116 337600
rect 281592 337560 281598 337572
rect 284110 337560 284116 337572
rect 284168 337560 284174 337612
rect 281626 335180 281632 335232
rect 281684 335220 281690 335232
rect 284018 335220 284024 335232
rect 281684 335192 284024 335220
rect 281684 335180 281690 335192
rect 284018 335180 284024 335192
rect 284076 335180 284082 335232
rect 281534 333208 281540 333260
rect 281592 333248 281598 333260
rect 283926 333248 283932 333260
rect 281592 333220 283932 333248
rect 281592 333208 281598 333220
rect 283926 333208 283932 333220
rect 283984 333208 283990 333260
rect 281534 331100 281540 331152
rect 281592 331140 281598 331152
rect 283834 331140 283840 331152
rect 281592 331112 283840 331140
rect 281592 331100 281598 331112
rect 283834 331100 283840 331112
rect 283892 331100 283898 331152
rect 281534 329060 281540 329112
rect 281592 329100 281598 329112
rect 283742 329100 283748 329112
rect 281592 329072 283748 329100
rect 281592 329060 281598 329072
rect 283742 329060 283748 329072
rect 283800 329060 283806 329112
rect 281534 327020 281540 327072
rect 281592 327060 281598 327072
rect 283650 327060 283656 327072
rect 281592 327032 283656 327060
rect 281592 327020 281598 327032
rect 283650 327020 283656 327032
rect 283708 327020 283714 327072
rect 281534 325048 281540 325100
rect 281592 325088 281598 325100
rect 283558 325088 283564 325100
rect 281592 325060 283564 325088
rect 281592 325048 281598 325060
rect 283558 325048 283564 325060
rect 283616 325048 283622 325100
rect 135990 318996 135996 319048
rect 136048 319036 136054 319048
rect 136542 319036 136548 319048
rect 136048 319008 136548 319036
rect 136048 318996 136054 319008
rect 136542 318996 136548 319008
rect 136600 318996 136606 319048
rect 59354 318928 59360 318980
rect 59412 318968 59418 318980
rect 60274 318968 60280 318980
rect 59412 318940 60280 318968
rect 59412 318928 59418 318940
rect 60274 318928 60280 318940
rect 60332 318928 60338 318980
rect 60277 318835 60335 318841
rect 60277 318801 60289 318835
rect 60323 318832 60335 318835
rect 61013 318835 61071 318841
rect 61013 318832 61025 318835
rect 60323 318804 61025 318832
rect 60323 318801 60335 318804
rect 60277 318795 60335 318801
rect 61013 318801 61025 318804
rect 61059 318801 61071 318835
rect 145650 318832 145656 318844
rect 61013 318795 61071 318801
rect 138032 318804 145656 318832
rect 30282 318724 30288 318776
rect 30340 318764 30346 318776
rect 70946 318764 70952 318776
rect 30340 318736 70952 318764
rect 30340 318724 30346 318736
rect 70946 318724 70952 318736
rect 71004 318724 71010 318776
rect 115842 318724 115848 318776
rect 115900 318764 115906 318776
rect 138032 318764 138060 318804
rect 145650 318792 145656 318804
rect 145708 318792 145714 318844
rect 152461 318835 152519 318841
rect 152461 318832 152473 318835
rect 150268 318804 152473 318832
rect 115900 318736 138060 318764
rect 115900 318724 115906 318736
rect 138106 318724 138112 318776
rect 138164 318764 138170 318776
rect 138164 318736 145788 318764
rect 138164 318724 138170 318736
rect 31662 318656 31668 318708
rect 31720 318696 31726 318708
rect 71774 318696 71780 318708
rect 31720 318668 71780 318696
rect 31720 318656 31726 318668
rect 71774 318656 71780 318668
rect 71832 318656 71838 318708
rect 99650 318656 99656 318708
rect 99708 318696 99714 318708
rect 105170 318696 105176 318708
rect 99708 318668 105176 318696
rect 99708 318656 99714 318668
rect 105170 318656 105176 318668
rect 105228 318656 105234 318708
rect 117130 318656 117136 318708
rect 117188 318696 117194 318708
rect 142985 318699 143043 318705
rect 117188 318668 142936 318696
rect 117188 318656 117194 318668
rect 30190 318588 30196 318640
rect 30248 318628 30254 318640
rect 71314 318628 71320 318640
rect 30248 318600 71320 318628
rect 30248 318588 30254 318600
rect 71314 318588 71320 318600
rect 71372 318588 71378 318640
rect 118510 318588 118516 318640
rect 118568 318628 118574 318640
rect 142801 318631 142859 318637
rect 142801 318628 142813 318631
rect 118568 318600 142813 318628
rect 118568 318588 118574 318600
rect 142801 318597 142813 318600
rect 142847 318597 142859 318631
rect 142908 318628 142936 318668
rect 142985 318665 142997 318699
rect 143031 318696 143043 318699
rect 145653 318699 145711 318705
rect 145653 318696 145665 318699
rect 143031 318668 145665 318696
rect 143031 318665 143043 318668
rect 142985 318659 143043 318665
rect 145653 318665 145665 318668
rect 145699 318665 145711 318699
rect 145760 318696 145788 318736
rect 148594 318724 148600 318776
rect 148652 318764 148658 318776
rect 150268 318764 150296 318804
rect 152461 318801 152473 318804
rect 152507 318801 152519 318835
rect 152461 318795 152519 318801
rect 217612 318804 219388 318832
rect 148652 318736 150296 318764
rect 148652 318724 148658 318736
rect 150342 318724 150348 318776
rect 150400 318764 150406 318776
rect 175826 318764 175832 318776
rect 150400 318736 175832 318764
rect 150400 318724 150406 318736
rect 175826 318724 175832 318736
rect 175884 318724 175890 318776
rect 210970 318724 210976 318776
rect 211028 318764 211034 318776
rect 217612 318764 217640 318804
rect 211028 318736 217640 318764
rect 211028 318724 211034 318736
rect 217686 318724 217692 318776
rect 217744 318764 217750 318776
rect 219253 318767 219311 318773
rect 219253 318764 219265 318767
rect 217744 318736 219265 318764
rect 217744 318724 217750 318736
rect 219253 318733 219265 318736
rect 219299 318733 219311 318767
rect 219360 318764 219388 318804
rect 293218 318764 293224 318776
rect 219360 318736 293224 318764
rect 219253 318727 219311 318733
rect 293218 318724 293224 318736
rect 293276 318724 293282 318776
rect 313274 318724 313280 318776
rect 313332 318764 313338 318776
rect 404998 318764 405004 318776
rect 313332 318736 405004 318764
rect 313332 318724 313338 318736
rect 404998 318724 405004 318736
rect 405056 318764 405062 318776
rect 443086 318764 443092 318776
rect 405056 318736 443092 318764
rect 405056 318724 405062 318736
rect 443086 318724 443092 318736
rect 443144 318724 443150 318776
rect 149793 318699 149851 318705
rect 149793 318696 149805 318699
rect 145760 318668 149805 318696
rect 145653 318659 145711 318665
rect 149793 318665 149805 318668
rect 149839 318665 149851 318699
rect 149793 318659 149851 318665
rect 149882 318656 149888 318708
rect 149940 318696 149946 318708
rect 162118 318696 162124 318708
rect 149940 318668 162124 318696
rect 149940 318656 149946 318668
rect 162118 318656 162124 318668
rect 162176 318656 162182 318708
rect 163866 318656 163872 318708
rect 163924 318696 163930 318708
rect 246298 318696 246304 318708
rect 163924 318668 246304 318696
rect 163924 318656 163930 318668
rect 246298 318656 246304 318668
rect 246356 318656 246362 318708
rect 143629 318631 143687 318637
rect 143629 318628 143641 318631
rect 142908 318600 143641 318628
rect 142801 318591 142859 318597
rect 143629 318597 143641 318600
rect 143675 318597 143687 318631
rect 143629 318591 143687 318597
rect 145006 318588 145012 318640
rect 145064 318628 145070 318640
rect 152369 318631 152427 318637
rect 152369 318628 152381 318631
rect 145064 318600 152381 318628
rect 145064 318588 145070 318600
rect 152369 318597 152381 318600
rect 152415 318597 152427 318631
rect 152369 318591 152427 318597
rect 152461 318631 152519 318637
rect 152461 318597 152473 318631
rect 152507 318628 152519 318631
rect 155405 318631 155463 318637
rect 155405 318628 155417 318631
rect 152507 318600 155417 318628
rect 152507 318597 152519 318600
rect 152461 318591 152519 318597
rect 155405 318597 155417 318600
rect 155451 318597 155463 318631
rect 155405 318591 155463 318597
rect 155770 318588 155776 318640
rect 155828 318628 155834 318640
rect 178586 318628 178592 318640
rect 155828 318600 178592 318628
rect 155828 318588 155834 318600
rect 178586 318588 178592 318600
rect 178644 318588 178650 318640
rect 186774 318588 186780 318640
rect 186832 318628 186838 318640
rect 193858 318628 193864 318640
rect 186832 318600 193864 318628
rect 186832 318588 186838 318600
rect 193858 318588 193864 318600
rect 193916 318588 193922 318640
rect 198826 318588 198832 318640
rect 198884 318628 198890 318640
rect 291838 318628 291844 318640
rect 198884 318600 291844 318628
rect 198884 318588 198890 318600
rect 291838 318588 291844 318600
rect 291896 318588 291902 318640
rect 23382 318520 23388 318572
rect 23440 318560 23446 318572
rect 61013 318563 61071 318569
rect 23440 318532 60872 318560
rect 23440 318520 23446 318532
rect 27522 318452 27528 318504
rect 27580 318492 27586 318504
rect 60737 318495 60795 318501
rect 60737 318492 60749 318495
rect 27580 318464 60749 318492
rect 27580 318452 27586 318464
rect 60737 318461 60749 318464
rect 60783 318461 60795 318495
rect 60844 318492 60872 318532
rect 61013 318529 61025 318563
rect 61059 318560 61071 318563
rect 64598 318560 64604 318572
rect 61059 318532 64604 318560
rect 61059 318529 61071 318532
rect 61013 318523 61071 318529
rect 64598 318520 64604 318532
rect 64656 318520 64662 318572
rect 111794 318520 111800 318572
rect 111852 318560 111858 318572
rect 133138 318560 133144 318572
rect 111852 318532 133144 318560
rect 111852 318520 111858 318532
rect 133138 318520 133144 318532
rect 133196 318520 133202 318572
rect 134242 318520 134248 318572
rect 134300 318560 134306 318572
rect 169018 318560 169024 318572
rect 134300 318532 169024 318560
rect 134300 318520 134306 318532
rect 169018 318520 169024 318532
rect 169076 318520 169082 318572
rect 177298 318520 177304 318572
rect 177356 318560 177362 318572
rect 189074 318560 189080 318572
rect 177356 318532 189080 318560
rect 177356 318520 177362 318532
rect 189074 318520 189080 318532
rect 189132 318520 189138 318572
rect 193490 318520 193496 318572
rect 193548 318560 193554 318572
rect 289078 318560 289084 318572
rect 193548 318532 289084 318560
rect 193548 318520 193554 318532
rect 289078 318520 289084 318532
rect 289136 318520 289142 318572
rect 68646 318492 68652 318504
rect 60844 318464 68652 318492
rect 60737 318455 60795 318461
rect 68646 318452 68652 318464
rect 68704 318452 68710 318504
rect 82078 318452 82084 318504
rect 82136 318492 82142 318504
rect 90174 318492 90180 318504
rect 82136 318464 90180 318492
rect 82136 318452 82142 318464
rect 90174 318452 90180 318464
rect 90232 318452 90238 318504
rect 124766 318452 124772 318504
rect 124824 318492 124830 318504
rect 160741 318495 160799 318501
rect 160741 318492 160753 318495
rect 124824 318464 160753 318492
rect 124824 318452 124830 318464
rect 160741 318461 160753 318464
rect 160787 318461 160799 318495
rect 160741 318455 160799 318461
rect 170582 318452 170588 318504
rect 170640 318492 170646 318504
rect 271509 318495 271567 318501
rect 271509 318492 271521 318495
rect 170640 318464 271521 318492
rect 170640 318452 170646 318464
rect 271509 318461 271521 318464
rect 271555 318461 271567 318495
rect 271509 318455 271567 318461
rect 272886 318452 272892 318504
rect 272944 318492 272950 318504
rect 277305 318495 277363 318501
rect 277305 318492 277317 318495
rect 272944 318464 277317 318492
rect 272944 318452 272950 318464
rect 277305 318461 277317 318464
rect 277351 318461 277363 318495
rect 277305 318455 277363 318461
rect 22002 318384 22008 318436
rect 22060 318424 22066 318436
rect 67726 318424 67732 318436
rect 22060 318396 67732 318424
rect 22060 318384 22066 318396
rect 67726 318384 67732 318396
rect 67784 318384 67790 318436
rect 79318 318384 79324 318436
rect 79376 318424 79382 318436
rect 87506 318424 87512 318436
rect 79376 318396 87512 318424
rect 79376 318384 79382 318396
rect 87506 318384 87512 318396
rect 87564 318384 87570 318436
rect 108574 318384 108580 318436
rect 108632 318424 108638 318436
rect 128630 318424 128636 318436
rect 108632 318396 128636 318424
rect 108632 318384 108638 318396
rect 128630 318384 128636 318396
rect 128688 318384 128694 318436
rect 130194 318384 130200 318436
rect 130252 318424 130258 318436
rect 167638 318424 167644 318436
rect 130252 318396 167644 318424
rect 130252 318384 130258 318396
rect 167638 318384 167644 318396
rect 167696 318384 167702 318436
rect 171962 318384 171968 318436
rect 172020 318424 172026 318436
rect 279418 318424 279424 318436
rect 172020 318396 279424 318424
rect 172020 318384 172026 318396
rect 279418 318384 279424 318396
rect 279476 318384 279482 318436
rect 20622 318316 20628 318368
rect 20680 318356 20686 318368
rect 67358 318356 67364 318368
rect 20680 318328 67364 318356
rect 20680 318316 20686 318328
rect 67358 318316 67364 318328
rect 67416 318316 67422 318368
rect 82722 318316 82728 318368
rect 82780 318356 82786 318368
rect 90634 318356 90640 318368
rect 82780 318328 90640 318356
rect 82780 318316 82786 318328
rect 90634 318316 90640 318328
rect 90692 318316 90698 318368
rect 126146 318316 126152 318368
rect 126204 318356 126210 318368
rect 164878 318356 164884 318368
rect 126204 318328 164884 318356
rect 126204 318316 126210 318328
rect 164878 318316 164884 318328
rect 164936 318316 164942 318368
rect 165154 318316 165160 318368
rect 165212 318356 165218 318368
rect 169757 318359 169815 318365
rect 169757 318356 169769 318359
rect 165212 318328 169769 318356
rect 165212 318316 165218 318328
rect 169757 318325 169769 318328
rect 169803 318325 169815 318359
rect 169757 318319 169815 318325
rect 174630 318316 174636 318368
rect 174688 318356 174694 318368
rect 286318 318356 286324 318368
rect 174688 318328 286324 318356
rect 174688 318316 174694 318328
rect 286318 318316 286324 318328
rect 286376 318316 286382 318368
rect 21910 318248 21916 318300
rect 21968 318288 21974 318300
rect 60734 318288 60740 318300
rect 21968 318260 60740 318288
rect 21968 318248 21974 318260
rect 60734 318248 60740 318260
rect 60792 318248 60798 318300
rect 60829 318291 60887 318297
rect 60829 318257 60841 318291
rect 60875 318288 60887 318291
rect 70026 318288 70032 318300
rect 60875 318260 70032 318288
rect 60875 318257 60887 318260
rect 60829 318251 60887 318257
rect 70026 318248 70032 318260
rect 70084 318248 70090 318300
rect 75178 318248 75184 318300
rect 75236 318288 75242 318300
rect 87046 318288 87052 318300
rect 75236 318260 87052 318288
rect 75236 318248 75242 318260
rect 87046 318248 87052 318260
rect 87104 318248 87110 318300
rect 107286 318248 107292 318300
rect 107344 318288 107350 318300
rect 124401 318291 124459 318297
rect 124401 318288 124413 318291
rect 107344 318260 124413 318288
rect 107344 318248 107350 318260
rect 124401 318257 124413 318260
rect 124447 318257 124459 318291
rect 124401 318251 124459 318257
rect 127434 318248 127440 318300
rect 127492 318288 127498 318300
rect 166350 318288 166356 318300
rect 127492 318260 166356 318288
rect 127492 318248 127498 318260
rect 166350 318248 166356 318260
rect 166408 318248 166414 318300
rect 175918 318248 175924 318300
rect 175976 318288 175982 318300
rect 304258 318288 304264 318300
rect 175976 318260 304264 318288
rect 175976 318248 175982 318260
rect 304258 318248 304264 318260
rect 304316 318248 304322 318300
rect 60921 318223 60979 318229
rect 60921 318189 60933 318223
rect 60967 318220 60979 318223
rect 313274 318220 313280 318232
rect 60967 318192 313280 318220
rect 60967 318189 60979 318192
rect 60921 318183 60979 318189
rect 313274 318180 313280 318192
rect 313332 318180 313338 318232
rect 17862 318112 17868 318164
rect 17920 318152 17926 318164
rect 66438 318152 66444 318164
rect 17920 318124 66444 318152
rect 17920 318112 17926 318124
rect 66438 318112 66444 318124
rect 66496 318112 66502 318164
rect 87966 318152 87972 318164
rect 84028 318124 87972 318152
rect 13722 318044 13728 318096
rect 13780 318084 13786 318096
rect 60277 318087 60335 318093
rect 60277 318084 60289 318087
rect 13780 318056 60289 318084
rect 13780 318044 13786 318056
rect 60277 318053 60289 318056
rect 60323 318053 60335 318087
rect 60277 318047 60335 318053
rect 60366 318044 60372 318096
rect 60424 318084 60430 318096
rect 60645 318087 60703 318093
rect 60645 318084 60657 318087
rect 60424 318056 60657 318084
rect 60424 318044 60430 318056
rect 60645 318053 60657 318056
rect 60691 318053 60703 318087
rect 60645 318047 60703 318053
rect 60734 318044 60740 318096
rect 60792 318084 60798 318096
rect 68186 318084 68192 318096
rect 60792 318056 68192 318084
rect 60792 318044 60798 318056
rect 68186 318044 68192 318056
rect 68244 318044 68250 318096
rect 74442 318044 74448 318096
rect 74500 318084 74506 318096
rect 84028 318084 84056 318124
rect 87966 318112 87972 318124
rect 88024 318112 88030 318164
rect 122098 318112 122104 318164
rect 122156 318152 122162 318164
rect 152461 318155 152519 318161
rect 152461 318152 152473 318155
rect 122156 318124 152473 318152
rect 122156 318112 122162 318124
rect 152461 318121 152473 318124
rect 152507 318121 152519 318155
rect 152461 318115 152519 318121
rect 166994 318112 167000 318164
rect 167052 318152 167058 318164
rect 168282 318152 168288 318164
rect 167052 318124 168288 318152
rect 167052 318112 167058 318124
rect 168282 318112 168288 318124
rect 168340 318112 168346 318164
rect 169757 318155 169815 318161
rect 168668 318124 169708 318152
rect 74500 318056 84056 318084
rect 74500 318044 74506 318056
rect 87598 318044 87604 318096
rect 87656 318084 87662 318096
rect 89806 318084 89812 318096
rect 87656 318056 89812 318084
rect 87656 318044 87662 318056
rect 89806 318044 89812 318056
rect 89864 318044 89870 318096
rect 98730 318044 98736 318096
rect 98788 318084 98794 318096
rect 102410 318084 102416 318096
rect 98788 318056 102416 318084
rect 98788 318044 98794 318056
rect 102410 318044 102416 318056
rect 102468 318044 102474 318096
rect 102778 318044 102784 318096
rect 102836 318084 102842 318096
rect 103330 318084 103336 318096
rect 102836 318056 103336 318084
rect 102836 318044 102842 318056
rect 103330 318044 103336 318056
rect 103388 318044 103394 318096
rect 104986 318044 104992 318096
rect 105044 318084 105050 318096
rect 105722 318084 105728 318096
rect 105044 318056 105728 318084
rect 105044 318044 105050 318056
rect 105722 318044 105728 318056
rect 105780 318044 105786 318096
rect 107746 318044 107752 318096
rect 107804 318084 107810 318096
rect 108850 318084 108856 318096
rect 107804 318056 108856 318084
rect 107804 318044 107810 318056
rect 108850 318044 108856 318056
rect 108908 318044 108914 318096
rect 120718 318044 120724 318096
rect 120776 318084 120782 318096
rect 152645 318087 152703 318093
rect 152645 318084 152657 318087
rect 120776 318056 152657 318084
rect 120776 318044 120782 318056
rect 152645 318053 152657 318056
rect 152691 318053 152703 318087
rect 152645 318047 152703 318053
rect 152737 318087 152795 318093
rect 152737 318053 152749 318087
rect 152783 318084 152795 318087
rect 153838 318084 153844 318096
rect 152783 318056 153844 318084
rect 152783 318053 152795 318056
rect 152737 318047 152795 318053
rect 153838 318044 153844 318056
rect 153896 318044 153902 318096
rect 155310 318044 155316 318096
rect 155368 318084 155374 318096
rect 155770 318084 155776 318096
rect 155368 318056 155776 318084
rect 155368 318044 155374 318056
rect 155770 318044 155776 318056
rect 155828 318044 155834 318096
rect 167454 318044 167460 318096
rect 167512 318084 167518 318096
rect 168190 318084 168196 318096
rect 167512 318056 168196 318084
rect 167512 318044 167518 318056
rect 168190 318044 168196 318056
rect 168248 318044 168254 318096
rect 38470 317976 38476 318028
rect 38528 318016 38534 318028
rect 74534 318016 74540 318028
rect 38528 317988 74540 318016
rect 38528 317976 38534 317988
rect 74534 317976 74540 317988
rect 74592 317976 74598 318028
rect 88242 317976 88248 318028
rect 88300 318016 88306 318028
rect 92934 318016 92940 318028
rect 88300 317988 92940 318016
rect 88300 317976 88306 317988
rect 92934 317976 92940 317988
rect 92992 317976 92998 318028
rect 110414 317976 110420 318028
rect 110472 318016 110478 318028
rect 127618 318016 127624 318028
rect 110472 317988 127624 318016
rect 110472 317976 110478 317988
rect 127618 317976 127624 317988
rect 127676 317976 127682 318028
rect 138017 318019 138075 318025
rect 138017 317985 138029 318019
rect 138063 318016 138075 318019
rect 147493 318019 147551 318025
rect 147493 318016 147505 318019
rect 138063 317988 147505 318016
rect 138063 317985 138075 317988
rect 138017 317979 138075 317985
rect 147493 317985 147505 317988
rect 147539 317985 147551 318019
rect 147493 317979 147551 317985
rect 147769 318019 147827 318025
rect 147769 317985 147781 318019
rect 147815 318016 147827 318019
rect 151449 318019 151507 318025
rect 151449 318016 151461 318019
rect 147815 317988 151461 318016
rect 147815 317985 147827 317988
rect 147769 317979 147827 317985
rect 151449 317985 151461 317988
rect 151495 317985 151507 318019
rect 151449 317979 151507 317985
rect 152185 318019 152243 318025
rect 152185 317985 152197 318019
rect 152231 318016 152243 318019
rect 166258 318016 166264 318028
rect 152231 317988 166264 318016
rect 152231 317985 152243 317988
rect 152185 317979 152243 317985
rect 166258 317976 166264 317988
rect 166316 317976 166322 318028
rect 167914 317976 167920 318028
rect 167972 318016 167978 318028
rect 168668 318016 168696 318124
rect 168742 318044 168748 318096
rect 168800 318084 168806 318096
rect 169570 318084 169576 318096
rect 168800 318056 169576 318084
rect 168800 318044 168806 318056
rect 169570 318044 169576 318056
rect 169628 318044 169634 318096
rect 169680 318084 169708 318124
rect 169757 318121 169769 318155
rect 169803 318152 169815 318155
rect 248601 318155 248659 318161
rect 248601 318152 248613 318155
rect 169803 318124 248613 318152
rect 169803 318121 169815 318124
rect 169757 318115 169815 318121
rect 248601 318121 248613 318124
rect 248647 318121 248659 318155
rect 248601 318115 248659 318121
rect 248690 318112 248696 318164
rect 248748 318152 248754 318164
rect 249610 318152 249616 318164
rect 248748 318124 249616 318152
rect 248748 318112 248754 318124
rect 249610 318112 249616 318124
rect 249668 318112 249674 318164
rect 250070 318112 250076 318164
rect 250128 318152 250134 318164
rect 250990 318152 250996 318164
rect 250128 318124 250996 318152
rect 250128 318112 250134 318124
rect 250990 318112 250996 318124
rect 251048 318112 251054 318164
rect 251358 318112 251364 318164
rect 251416 318152 251422 318164
rect 252370 318152 252376 318164
rect 251416 318124 252376 318152
rect 251416 318112 251422 318124
rect 252370 318112 252376 318124
rect 252428 318112 252434 318164
rect 252738 318112 252744 318164
rect 252796 318152 252802 318164
rect 253658 318152 253664 318164
rect 252796 318124 253664 318152
rect 252796 318112 252802 318124
rect 253658 318112 253664 318124
rect 253716 318112 253722 318164
rect 254026 318112 254032 318164
rect 254084 318152 254090 318164
rect 255038 318152 255044 318164
rect 254084 318124 255044 318152
rect 254084 318112 254090 318124
rect 255038 318112 255044 318124
rect 255096 318112 255102 318164
rect 255406 318112 255412 318164
rect 255464 318152 255470 318164
rect 256418 318152 256424 318164
rect 255464 318124 256424 318152
rect 255464 318112 255470 318124
rect 256418 318112 256424 318124
rect 256476 318112 256482 318164
rect 256786 318112 256792 318164
rect 256844 318152 256850 318164
rect 257798 318152 257804 318164
rect 256844 318124 257804 318152
rect 256844 318112 256850 318124
rect 257798 318112 257804 318124
rect 257856 318112 257862 318164
rect 258074 318112 258080 318164
rect 258132 318152 258138 318164
rect 259178 318152 259184 318164
rect 258132 318124 259184 318152
rect 258132 318112 258138 318124
rect 259178 318112 259184 318124
rect 259236 318112 259242 318164
rect 259914 318112 259920 318164
rect 259972 318152 259978 318164
rect 260742 318152 260748 318164
rect 259972 318124 260748 318152
rect 259972 318112 259978 318124
rect 260742 318112 260748 318124
rect 260800 318112 260806 318164
rect 261846 318112 261852 318164
rect 261904 318152 261910 318164
rect 262122 318152 262128 318164
rect 261904 318124 262128 318152
rect 261904 318112 261910 318124
rect 262122 318112 262128 318124
rect 262180 318112 262186 318164
rect 263318 318112 263324 318164
rect 263376 318152 263382 318164
rect 263502 318152 263508 318164
rect 263376 318124 263508 318152
rect 263376 318112 263382 318124
rect 263502 318112 263508 318124
rect 263560 318112 263566 318164
rect 264698 318112 264704 318164
rect 264756 318152 264762 318164
rect 264882 318152 264888 318164
rect 264756 318124 264888 318152
rect 264756 318112 264762 318124
rect 264882 318112 264888 318124
rect 264940 318112 264946 318164
rect 265250 318112 265256 318164
rect 265308 318152 265314 318164
rect 266262 318152 266268 318164
rect 265308 318124 266268 318152
rect 265308 318112 265314 318124
rect 266262 318112 266268 318124
rect 266320 318112 266326 318164
rect 267090 318112 267096 318164
rect 267148 318152 267154 318164
rect 267550 318152 267556 318164
rect 267148 318124 267556 318152
rect 267148 318112 267154 318124
rect 267550 318112 267556 318124
rect 267608 318112 267614 318164
rect 268010 318112 268016 318164
rect 268068 318152 268074 318164
rect 269022 318152 269028 318164
rect 268068 318124 269028 318152
rect 268068 318112 268074 318124
rect 269022 318112 269028 318124
rect 269080 318112 269086 318164
rect 269298 318112 269304 318164
rect 269356 318152 269362 318164
rect 270402 318152 270408 318164
rect 269356 318124 270408 318152
rect 269356 318112 269362 318124
rect 270402 318112 270408 318124
rect 270460 318112 270466 318164
rect 270678 318112 270684 318164
rect 270736 318152 270742 318164
rect 271782 318152 271788 318164
rect 270736 318124 271788 318152
rect 270736 318112 270742 318124
rect 271782 318112 271788 318124
rect 271840 318112 271846 318164
rect 272518 318112 272524 318164
rect 272576 318152 272582 318164
rect 273070 318152 273076 318164
rect 272576 318124 273076 318152
rect 272576 318112 272582 318124
rect 273070 318112 273076 318124
rect 273128 318112 273134 318164
rect 273346 318112 273352 318164
rect 273404 318152 273410 318164
rect 274542 318152 274548 318164
rect 273404 318124 274548 318152
rect 273404 318112 273410 318124
rect 274542 318112 274548 318124
rect 274600 318112 274606 318164
rect 275646 318112 275652 318164
rect 275704 318152 275710 318164
rect 529382 318152 529388 318164
rect 275704 318124 529388 318152
rect 275704 318112 275710 318124
rect 529382 318112 529388 318124
rect 529440 318112 529446 318164
rect 268381 318087 268439 318093
rect 268381 318084 268393 318087
rect 169680 318056 268393 318084
rect 268381 318053 268393 318056
rect 268427 318053 268439 318087
rect 268381 318047 268439 318053
rect 268470 318044 268476 318096
rect 268528 318084 268534 318096
rect 268930 318084 268936 318096
rect 268528 318056 268936 318084
rect 268528 318044 268534 318056
rect 268930 318044 268936 318056
rect 268988 318044 268994 318096
rect 269758 318044 269764 318096
rect 269816 318084 269822 318096
rect 270310 318084 270316 318096
rect 269816 318056 270316 318084
rect 269816 318044 269822 318056
rect 270310 318044 270316 318056
rect 270368 318044 270374 318096
rect 271138 318044 271144 318096
rect 271196 318084 271202 318096
rect 271690 318084 271696 318096
rect 271196 318056 271696 318084
rect 271196 318044 271202 318056
rect 271690 318044 271696 318056
rect 271748 318044 271754 318096
rect 272058 318044 272064 318096
rect 272116 318084 272122 318096
rect 273162 318084 273168 318096
rect 272116 318056 273168 318084
rect 272116 318044 272122 318056
rect 273162 318044 273168 318056
rect 273220 318044 273226 318096
rect 273806 318044 273812 318096
rect 273864 318084 273870 318096
rect 274450 318084 274456 318096
rect 273864 318056 274456 318084
rect 273864 318044 273870 318056
rect 274450 318044 274456 318056
rect 274508 318044 274514 318096
rect 274726 318044 274732 318096
rect 274784 318084 274790 318096
rect 275922 318084 275928 318096
rect 274784 318056 275928 318084
rect 274784 318044 274790 318056
rect 275922 318044 275928 318056
rect 275980 318044 275986 318096
rect 276474 318044 276480 318096
rect 276532 318084 276538 318096
rect 277210 318084 277216 318096
rect 276532 318056 277216 318084
rect 276532 318044 276538 318056
rect 277210 318044 277216 318056
rect 277268 318044 277274 318096
rect 277305 318087 277363 318093
rect 277305 318053 277317 318087
rect 277351 318084 277363 318087
rect 529474 318084 529480 318096
rect 277351 318056 529480 318084
rect 277351 318053 277363 318056
rect 277305 318047 277363 318053
rect 529474 318044 529480 318056
rect 529532 318044 529538 318096
rect 167972 317988 168696 318016
rect 167972 317976 167978 317988
rect 169202 317976 169208 318028
rect 169260 318016 169266 318028
rect 169260 317988 180932 318016
rect 169260 317976 169266 317988
rect 37182 317908 37188 317960
rect 37240 317948 37246 317960
rect 73614 317948 73620 317960
rect 37240 317920 73620 317948
rect 37240 317908 37246 317920
rect 73614 317908 73620 317920
rect 73672 317908 73678 317960
rect 79410 317908 79416 317960
rect 79468 317948 79474 317960
rect 83458 317948 83464 317960
rect 79468 317920 83464 317948
rect 79468 317908 79474 317920
rect 83458 317908 83464 317920
rect 83516 317908 83522 317960
rect 85482 317908 85488 317960
rect 85540 317948 85546 317960
rect 92014 317948 92020 317960
rect 85540 317920 92020 317948
rect 85540 317908 85546 317920
rect 92014 317908 92020 317920
rect 92072 317908 92078 317960
rect 130654 317908 130660 317960
rect 130712 317948 130718 317960
rect 134610 317948 134616 317960
rect 130712 317920 134616 317948
rect 130712 317908 130718 317920
rect 134610 317908 134616 317920
rect 134668 317908 134674 317960
rect 134702 317908 134708 317960
rect 134760 317948 134766 317960
rect 143537 317951 143595 317957
rect 143537 317948 143549 317951
rect 134760 317920 143549 317948
rect 134760 317908 134766 317920
rect 143537 317917 143549 317920
rect 143583 317917 143595 317951
rect 143537 317911 143595 317917
rect 143629 317951 143687 317957
rect 143629 317917 143641 317951
rect 143675 317948 143687 317951
rect 146665 317951 146723 317957
rect 146665 317948 146677 317951
rect 143675 317920 146677 317948
rect 143675 317917 143687 317920
rect 143629 317911 143687 317917
rect 146665 317917 146677 317920
rect 146711 317917 146723 317951
rect 146665 317911 146723 317917
rect 146754 317908 146760 317960
rect 146812 317948 146818 317960
rect 147582 317948 147588 317960
rect 146812 317920 147588 317948
rect 146812 317908 146818 317920
rect 147582 317908 147588 317920
rect 147640 317908 147646 317960
rect 147674 317908 147680 317960
rect 147732 317948 147738 317960
rect 148870 317948 148876 317960
rect 147732 317920 148876 317948
rect 147732 317908 147738 317920
rect 148870 317908 148876 317920
rect 148928 317908 148934 317960
rect 149793 317951 149851 317957
rect 149793 317917 149805 317951
rect 149839 317948 149851 317951
rect 152369 317951 152427 317957
rect 149839 317920 152320 317948
rect 149839 317917 149851 317920
rect 149793 317911 149851 317917
rect 44082 317840 44088 317892
rect 44140 317880 44146 317892
rect 76282 317880 76288 317892
rect 44140 317852 76288 317880
rect 44140 317840 44146 317852
rect 76282 317840 76288 317852
rect 76340 317840 76346 317892
rect 89622 317840 89628 317892
rect 89680 317880 89686 317892
rect 93394 317880 93400 317892
rect 89680 317852 93400 317880
rect 89680 317840 89686 317852
rect 93394 317840 93400 317852
rect 93452 317840 93458 317892
rect 98270 317840 98276 317892
rect 98328 317880 98334 317892
rect 100110 317880 100116 317892
rect 98328 317852 100116 317880
rect 98328 317840 98334 317852
rect 100110 317840 100116 317852
rect 100168 317840 100174 317892
rect 127066 317840 127072 317892
rect 127124 317880 127130 317892
rect 128262 317880 128268 317892
rect 127124 317852 128268 317880
rect 127124 317840 127130 317852
rect 128262 317840 128268 317852
rect 128320 317840 128326 317892
rect 129274 317840 129280 317892
rect 129332 317880 129338 317892
rect 138017 317883 138075 317889
rect 138017 317880 138029 317883
rect 129332 317852 138029 317880
rect 129332 317840 129338 317852
rect 138017 317849 138029 317852
rect 138063 317849 138075 317883
rect 138017 317843 138075 317849
rect 138109 317883 138167 317889
rect 138109 317849 138121 317883
rect 138155 317880 138167 317883
rect 152185 317883 152243 317889
rect 152185 317880 152197 317883
rect 138155 317852 152197 317880
rect 138155 317849 138167 317852
rect 138109 317843 138167 317849
rect 152185 317849 152197 317852
rect 152231 317849 152243 317883
rect 152292 317880 152320 317920
rect 152369 317917 152381 317951
rect 152415 317948 152427 317951
rect 162121 317951 162179 317957
rect 162121 317948 162133 317951
rect 152415 317920 162133 317948
rect 152415 317917 152427 317920
rect 152369 317911 152427 317917
rect 162121 317917 162133 317920
rect 162167 317917 162179 317951
rect 162121 317911 162179 317917
rect 170122 317908 170128 317960
rect 170180 317948 170186 317960
rect 171042 317948 171048 317960
rect 170180 317920 171048 317948
rect 170180 317908 170186 317920
rect 171042 317908 171048 317920
rect 171100 317908 171106 317960
rect 172790 317908 172796 317960
rect 172848 317948 172854 317960
rect 173710 317948 173716 317960
rect 172848 317920 173716 317948
rect 172848 317908 172854 317920
rect 173710 317908 173716 317920
rect 173768 317908 173774 317960
rect 174170 317908 174176 317960
rect 174228 317948 174234 317960
rect 175090 317948 175096 317960
rect 174228 317920 175096 317948
rect 174228 317908 174234 317920
rect 175090 317908 175096 317920
rect 175148 317908 175154 317960
rect 176838 317908 176844 317960
rect 176896 317948 176902 317960
rect 177850 317948 177856 317960
rect 176896 317920 177856 317948
rect 176896 317908 176902 317920
rect 177850 317908 177856 317920
rect 177908 317908 177914 317960
rect 178218 317908 178224 317960
rect 178276 317948 178282 317960
rect 179230 317948 179236 317960
rect 178276 317920 179236 317948
rect 178276 317908 178282 317920
rect 179230 317908 179236 317920
rect 179288 317908 179294 317960
rect 179506 317908 179512 317960
rect 179564 317948 179570 317960
rect 180610 317948 180616 317960
rect 179564 317920 180616 317948
rect 179564 317908 179570 317920
rect 180610 317908 180616 317920
rect 180668 317908 180674 317960
rect 180904 317948 180932 317988
rect 182266 317976 182272 318028
rect 182324 318016 182330 318028
rect 183370 318016 183376 318028
rect 182324 317988 183376 318016
rect 182324 317976 182330 317988
rect 183370 317976 183376 317988
rect 183428 317976 183434 318028
rect 183554 317976 183560 318028
rect 183612 318016 183618 318028
rect 184750 318016 184756 318028
rect 183612 317988 184756 318016
rect 183612 317976 183618 317988
rect 184750 317976 184756 317988
rect 184808 317976 184814 318028
rect 184934 317976 184940 318028
rect 184992 318016 184998 318028
rect 186130 318016 186136 318028
rect 184992 317988 186136 318016
rect 184992 317976 184998 317988
rect 186130 317976 186136 317988
rect 186188 317976 186194 318028
rect 186314 317976 186320 318028
rect 186372 318016 186378 318028
rect 187418 318016 187424 318028
rect 186372 317988 187424 318016
rect 186372 317976 186378 317988
rect 187418 317976 187424 317988
rect 187476 317976 187482 318028
rect 188522 317976 188528 318028
rect 188580 318016 188586 318028
rect 188982 318016 188988 318028
rect 188580 317988 188988 318016
rect 188580 317976 188586 317988
rect 188982 317976 188988 317988
rect 189040 317976 189046 318028
rect 189902 317976 189908 318028
rect 189960 318016 189966 318028
rect 190362 318016 190368 318028
rect 189960 317988 190368 318016
rect 189960 317976 189966 317988
rect 190362 317976 190368 317988
rect 190420 317976 190426 318028
rect 191190 317976 191196 318028
rect 191248 318016 191254 318028
rect 191650 318016 191656 318028
rect 191248 317988 191656 318016
rect 191248 317976 191254 317988
rect 191650 317976 191656 317988
rect 191708 317976 191714 318028
rect 192110 317976 192116 318028
rect 192168 318016 192174 318028
rect 192938 318016 192944 318028
rect 192168 317988 192944 318016
rect 192168 317976 192174 317988
rect 192938 317976 192944 317988
rect 192996 317976 193002 318028
rect 193950 317976 193956 318028
rect 194008 318016 194014 318028
rect 194502 318016 194508 318028
rect 194008 317988 194508 318016
rect 194008 317976 194014 317988
rect 194502 317976 194508 317988
rect 194560 317976 194566 318028
rect 194778 317976 194784 318028
rect 194836 318016 194842 318028
rect 195698 318016 195704 318028
rect 194836 317988 195704 318016
rect 194836 317976 194842 317988
rect 195698 317976 195704 317988
rect 195756 317976 195762 318028
rect 196618 317976 196624 318028
rect 196676 318016 196682 318028
rect 197170 318016 197176 318028
rect 196676 317988 197176 318016
rect 196676 317976 196682 317988
rect 197170 317976 197176 317988
rect 197228 317976 197234 318028
rect 197538 317976 197544 318028
rect 197596 318016 197602 318028
rect 198458 318016 198464 318028
rect 197596 317988 198464 318016
rect 197596 317976 197602 317988
rect 198458 317976 198464 317988
rect 198516 317976 198522 318028
rect 199286 317976 199292 318028
rect 199344 318016 199350 318028
rect 200022 318016 200028 318028
rect 199344 317988 200028 318016
rect 199344 317976 199350 317988
rect 200022 317976 200028 317988
rect 200080 317976 200086 318028
rect 200206 317976 200212 318028
rect 200264 318016 200270 318028
rect 201218 318016 201224 318028
rect 200264 317988 201224 318016
rect 200264 317976 200270 317988
rect 201218 317976 201224 317988
rect 201276 317976 201282 318028
rect 201586 317976 201592 318028
rect 201644 318016 201650 318028
rect 202598 318016 202604 318028
rect 201644 317988 202604 318016
rect 201644 317976 201650 317988
rect 202598 317976 202604 317988
rect 202656 317976 202662 318028
rect 202874 317976 202880 318028
rect 202932 318016 202938 318028
rect 203978 318016 203984 318028
rect 202932 317988 203984 318016
rect 202932 317976 202938 317988
rect 203978 317976 203984 317988
rect 204036 317976 204042 318028
rect 205358 317976 205364 318028
rect 205416 318016 205422 318028
rect 205542 318016 205548 318028
rect 205416 317988 205548 318016
rect 205416 317976 205422 317988
rect 205542 317976 205548 317988
rect 205600 317976 205606 318028
rect 206002 317976 206008 318028
rect 206060 318016 206066 318028
rect 206830 318016 206836 318028
rect 206060 317988 206836 318016
rect 206060 317976 206066 317988
rect 206830 317976 206836 317988
rect 206888 317976 206894 318028
rect 207382 317976 207388 318028
rect 207440 318016 207446 318028
rect 208118 318016 208124 318028
rect 207440 317988 208124 318016
rect 207440 317976 207446 317988
rect 208118 317976 208124 317988
rect 208176 317976 208182 318028
rect 208762 317976 208768 318028
rect 208820 318016 208826 318028
rect 209590 318016 209596 318028
rect 208820 317988 209596 318016
rect 208820 317976 208826 317988
rect 209590 317976 209596 317988
rect 209648 317976 209654 318028
rect 210050 317976 210056 318028
rect 210108 318016 210114 318028
rect 211062 318016 211068 318028
rect 210108 317988 211068 318016
rect 210108 317976 210114 317988
rect 211062 317976 211068 317988
rect 211120 317976 211126 318028
rect 211430 317976 211436 318028
rect 211488 318016 211494 318028
rect 212442 318016 212448 318028
rect 211488 317988 212448 318016
rect 211488 317976 211494 317988
rect 212442 317976 212448 317988
rect 212500 317976 212506 318028
rect 213178 317976 213184 318028
rect 213236 318016 213242 318028
rect 213730 318016 213736 318028
rect 213236 317988 213736 318016
rect 213236 317976 213242 317988
rect 213730 317976 213736 317988
rect 213788 317976 213794 318028
rect 214098 317976 214104 318028
rect 214156 318016 214162 318028
rect 215110 318016 215116 318028
rect 214156 317988 215116 318016
rect 214156 317976 214162 317988
rect 215110 317976 215116 317988
rect 215168 317976 215174 318028
rect 215938 317976 215944 318028
rect 215996 318016 216002 318028
rect 216490 318016 216496 318028
rect 215996 317988 216496 318016
rect 215996 317976 216002 317988
rect 216490 317976 216496 317988
rect 216548 317976 216554 318028
rect 216766 317976 216772 318028
rect 216824 318016 216830 318028
rect 217962 318016 217968 318028
rect 216824 317988 217968 318016
rect 216824 317976 216830 317988
rect 217962 317976 217968 317988
rect 218020 317976 218026 318028
rect 219253 318019 219311 318025
rect 219253 317985 219265 318019
rect 219299 318016 219311 318019
rect 295978 318016 295984 318028
rect 219299 317988 295984 318016
rect 219299 317985 219311 317988
rect 219253 317979 219311 317985
rect 295978 317976 295984 317988
rect 296036 317976 296042 318028
rect 184198 317948 184204 317960
rect 180720 317920 180840 317948
rect 180904 317920 184204 317948
rect 152737 317883 152795 317889
rect 152737 317880 152749 317883
rect 152292 317852 152749 317880
rect 152185 317843 152243 317849
rect 152737 317849 152749 317852
rect 152783 317849 152795 317883
rect 152737 317843 152795 317849
rect 153102 317840 153108 317892
rect 153160 317880 153166 317892
rect 176010 317880 176016 317892
rect 153160 317852 176016 317880
rect 153160 317840 153166 317852
rect 176010 317840 176016 317852
rect 176068 317840 176074 317892
rect 180720 317880 180748 317920
rect 180628 317852 180748 317880
rect 180812 317880 180840 317920
rect 184198 317908 184204 317920
rect 184256 317908 184262 317960
rect 184290 317908 184296 317960
rect 184348 317948 184354 317960
rect 184348 317920 187096 317948
rect 184348 317908 184354 317920
rect 185578 317880 185584 317892
rect 180812 317852 185584 317880
rect 38562 317772 38568 317824
rect 38620 317812 38626 317824
rect 74074 317812 74080 317824
rect 38620 317784 74080 317812
rect 38620 317772 38626 317784
rect 74074 317772 74080 317784
rect 74132 317772 74138 317824
rect 84838 317772 84844 317824
rect 84896 317812 84902 317824
rect 91554 317812 91560 317824
rect 84896 317784 91560 317812
rect 84896 317772 84902 317784
rect 91554 317772 91560 317784
rect 91612 317772 91618 317824
rect 113082 317772 113088 317824
rect 113140 317812 113146 317824
rect 115937 317815 115995 317821
rect 115937 317812 115949 317815
rect 113140 317784 115949 317812
rect 113140 317772 113146 317784
rect 115937 317781 115949 317784
rect 115983 317781 115995 317815
rect 115937 317775 115995 317781
rect 127894 317772 127900 317824
rect 127952 317812 127958 317824
rect 148410 317812 148416 317824
rect 127952 317784 148416 317812
rect 127952 317772 127958 317784
rect 148410 317772 148416 317784
rect 148468 317772 148474 317824
rect 149054 317772 149060 317824
rect 149112 317812 149118 317824
rect 151357 317815 151415 317821
rect 151357 317812 151369 317815
rect 149112 317784 151369 317812
rect 149112 317772 149118 317784
rect 151357 317781 151369 317784
rect 151403 317781 151415 317815
rect 151357 317775 151415 317781
rect 151449 317815 151507 317821
rect 151449 317781 151461 317815
rect 151495 317812 151507 317815
rect 155218 317812 155224 317824
rect 151495 317784 155224 317812
rect 151495 317781 151507 317784
rect 151449 317775 151507 317781
rect 155218 317772 155224 317784
rect 155276 317772 155282 317824
rect 155313 317815 155371 317821
rect 155313 317781 155325 317815
rect 155359 317812 155371 317815
rect 173158 317812 173164 317824
rect 155359 317784 173164 317812
rect 155359 317781 155371 317784
rect 155313 317775 155371 317781
rect 173158 317772 173164 317784
rect 173216 317772 173222 317824
rect 173250 317772 173256 317824
rect 173308 317812 173314 317824
rect 180628 317812 180656 317852
rect 185578 317840 185584 317852
rect 185636 317840 185642 317892
rect 187068 317880 187096 317920
rect 187142 317908 187148 317960
rect 187200 317948 187206 317960
rect 187602 317948 187608 317960
rect 187200 317920 187608 317948
rect 187200 317908 187206 317920
rect 187602 317908 187608 317920
rect 187660 317908 187666 317960
rect 192570 317908 192576 317960
rect 192628 317948 192634 317960
rect 193122 317948 193128 317960
rect 192628 317920 193128 317948
rect 192628 317908 192634 317920
rect 193122 317908 193128 317920
rect 193180 317908 193186 317960
rect 195238 317908 195244 317960
rect 195296 317948 195302 317960
rect 195882 317948 195888 317960
rect 195296 317920 195888 317948
rect 195296 317908 195302 317920
rect 195882 317908 195888 317920
rect 195940 317908 195946 317960
rect 196158 317908 196164 317960
rect 196216 317948 196222 317960
rect 197262 317948 197268 317960
rect 196216 317920 197268 317948
rect 196216 317908 196222 317920
rect 197262 317908 197268 317920
rect 197320 317908 197326 317960
rect 200666 317908 200672 317960
rect 200724 317948 200730 317960
rect 201402 317948 201408 317960
rect 200724 317920 201408 317948
rect 200724 317908 200730 317920
rect 201402 317908 201408 317920
rect 201460 317908 201466 317960
rect 203334 317908 203340 317960
rect 203392 317948 203398 317960
rect 204162 317948 204168 317960
rect 203392 317920 204168 317948
rect 203392 317908 203398 317920
rect 204162 317908 204168 317920
rect 204220 317908 204226 317960
rect 207842 317908 207848 317960
rect 207900 317948 207906 317960
rect 208302 317948 208308 317960
rect 207900 317920 208308 317948
rect 207900 317908 207906 317920
rect 208302 317908 208308 317920
rect 208360 317908 208366 317960
rect 212810 317908 212816 317960
rect 212868 317948 212874 317960
rect 213822 317948 213828 317960
rect 212868 317920 213828 317948
rect 212868 317908 212874 317920
rect 213822 317908 213828 317920
rect 213880 317908 213886 317960
rect 215478 317908 215484 317960
rect 215536 317948 215542 317960
rect 216582 317948 216588 317960
rect 215536 317920 216588 317948
rect 215536 317908 215542 317920
rect 216582 317908 216588 317920
rect 216640 317908 216646 317960
rect 217226 317908 217232 317960
rect 217284 317948 217290 317960
rect 217870 317948 217876 317960
rect 217284 317920 217876 317948
rect 217284 317908 217290 317920
rect 217870 317908 217876 317920
rect 217928 317908 217934 317960
rect 218146 317908 218152 317960
rect 218204 317948 218210 317960
rect 219342 317948 219348 317960
rect 218204 317920 219348 317948
rect 218204 317908 218210 317920
rect 219342 317908 219348 317920
rect 219400 317908 219406 317960
rect 219986 317908 219992 317960
rect 220044 317948 220050 317960
rect 220630 317948 220636 317960
rect 220044 317920 220636 317948
rect 220044 317908 220050 317920
rect 220630 317908 220636 317920
rect 220688 317908 220694 317960
rect 220814 317908 220820 317960
rect 220872 317948 220878 317960
rect 222010 317948 222016 317960
rect 220872 317920 222016 317948
rect 220872 317908 220878 317920
rect 222010 317908 222016 317920
rect 222068 317908 222074 317960
rect 222654 317908 222660 317960
rect 222712 317948 222718 317960
rect 223390 317948 223396 317960
rect 222712 317920 223396 317948
rect 222712 317908 222718 317920
rect 223390 317908 223396 317920
rect 223448 317908 223454 317960
rect 223574 317908 223580 317960
rect 223632 317948 223638 317960
rect 224862 317948 224868 317960
rect 223632 317920 224868 317948
rect 223632 317908 223638 317920
rect 224862 317908 224868 317920
rect 224920 317908 224926 317960
rect 225322 317908 225328 317960
rect 225380 317948 225386 317960
rect 226150 317948 226156 317960
rect 225380 317920 226156 317948
rect 225380 317908 225386 317920
rect 226150 317908 226156 317920
rect 226208 317908 226214 317960
rect 226702 317908 226708 317960
rect 226760 317948 226766 317960
rect 227530 317948 227536 317960
rect 226760 317920 227536 317948
rect 226760 317908 226766 317920
rect 227530 317908 227536 317920
rect 227588 317908 227594 317960
rect 227990 317908 227996 317960
rect 228048 317948 228054 317960
rect 228910 317948 228916 317960
rect 228048 317920 228916 317948
rect 228048 317908 228054 317920
rect 228910 317908 228916 317920
rect 228968 317908 228974 317960
rect 229005 317951 229063 317957
rect 229005 317917 229017 317951
rect 229051 317948 229063 317951
rect 296070 317948 296076 317960
rect 229051 317920 296076 317948
rect 229051 317917 229063 317920
rect 229005 317911 229063 317917
rect 296070 317908 296076 317920
rect 296128 317908 296134 317960
rect 253106 317880 253112 317892
rect 187068 317852 253112 317880
rect 253106 317840 253112 317852
rect 253164 317840 253170 317892
rect 253198 317840 253204 317892
rect 253256 317880 253262 317892
rect 253842 317880 253848 317892
rect 253256 317852 253848 317880
rect 253256 317840 253262 317852
rect 253842 317840 253848 317852
rect 253900 317840 253906 317892
rect 254486 317840 254492 317892
rect 254544 317880 254550 317892
rect 255222 317880 255228 317892
rect 254544 317852 255228 317880
rect 254544 317840 254550 317852
rect 255222 317840 255228 317852
rect 255280 317840 255286 317892
rect 255866 317840 255872 317892
rect 255924 317880 255930 317892
rect 256602 317880 256608 317892
rect 255924 317852 256608 317880
rect 255924 317840 255930 317852
rect 256602 317840 256608 317852
rect 256660 317840 256666 317892
rect 257246 317840 257252 317892
rect 257304 317880 257310 317892
rect 257982 317880 257988 317892
rect 257304 317852 257988 317880
rect 257304 317840 257310 317852
rect 257982 317840 257988 317852
rect 258040 317840 258046 317892
rect 258534 317840 258540 317892
rect 258592 317880 258598 317892
rect 259362 317880 259368 317892
rect 258592 317852 259368 317880
rect 258592 317840 258598 317852
rect 259362 317840 259368 317852
rect 259420 317840 259426 317892
rect 260834 317840 260840 317892
rect 260892 317880 260898 317892
rect 261938 317880 261944 317892
rect 260892 317852 261944 317880
rect 260892 317840 260898 317852
rect 261938 317840 261944 317852
rect 261996 317840 262002 317892
rect 263962 317840 263968 317892
rect 264020 317880 264026 317892
rect 264882 317880 264888 317892
rect 264020 317852 264888 317880
rect 264020 317840 264026 317852
rect 264882 317840 264888 317852
rect 264940 317840 264946 317892
rect 266630 317840 266636 317892
rect 266688 317880 266694 317892
rect 267642 317880 267648 317892
rect 266688 317852 267648 317880
rect 266688 317840 266694 317852
rect 267642 317840 267648 317852
rect 267700 317840 267706 317892
rect 268381 317883 268439 317889
rect 268381 317849 268393 317883
rect 268427 317880 268439 317883
rect 271138 317880 271144 317892
rect 268427 317852 271144 317880
rect 268427 317849 268439 317852
rect 268381 317843 268439 317849
rect 271138 317840 271144 317852
rect 271196 317840 271202 317892
rect 271509 317883 271567 317889
rect 271509 317849 271521 317883
rect 271555 317880 271567 317883
rect 275278 317880 275284 317892
rect 271555 317852 275284 317880
rect 271555 317849 271567 317852
rect 271509 317843 271567 317849
rect 275278 317840 275284 317852
rect 275336 317840 275342 317892
rect 276106 317840 276112 317892
rect 276164 317880 276170 317892
rect 277302 317880 277308 317892
rect 276164 317852 277308 317880
rect 276164 317840 276170 317852
rect 277302 317840 277308 317852
rect 277360 317840 277366 317892
rect 277854 317840 277860 317892
rect 277912 317880 277918 317892
rect 278590 317880 278596 317892
rect 277912 317852 278596 317880
rect 277912 317840 277918 317852
rect 278590 317840 278596 317852
rect 278648 317840 278654 317892
rect 278774 317840 278780 317892
rect 278832 317880 278838 317892
rect 280062 317880 280068 317892
rect 278832 317852 280068 317880
rect 278832 317840 278838 317852
rect 280062 317840 280068 317852
rect 280120 317840 280126 317892
rect 173308 317784 180656 317812
rect 173308 317772 173314 317784
rect 180886 317772 180892 317824
rect 180944 317812 180950 317824
rect 181990 317812 181996 317824
rect 180944 317784 181996 317812
rect 180944 317772 180950 317784
rect 181990 317772 181996 317784
rect 182048 317772 182054 317824
rect 185394 317772 185400 317824
rect 185452 317812 185458 317824
rect 189718 317812 189724 317824
rect 185452 317784 189724 317812
rect 185452 317772 185458 317784
rect 189718 317772 189724 317784
rect 189776 317772 189782 317824
rect 189905 317815 189963 317821
rect 189905 317781 189917 317815
rect 189951 317812 189963 317815
rect 250438 317812 250444 317824
rect 189951 317784 250444 317812
rect 189951 317781 189963 317784
rect 189905 317775 189963 317781
rect 250438 317772 250444 317784
rect 250496 317772 250502 317824
rect 261294 317772 261300 317824
rect 261352 317812 261358 317824
rect 262122 317812 262128 317824
rect 261352 317784 262128 317812
rect 261352 317772 261358 317784
rect 262122 317772 262128 317784
rect 262180 317772 262186 317824
rect 275186 317772 275192 317824
rect 275244 317812 275250 317824
rect 275830 317812 275836 317824
rect 275244 317784 275836 317812
rect 275244 317772 275250 317784
rect 275830 317772 275836 317784
rect 275888 317772 275894 317824
rect 277394 317772 277400 317824
rect 277452 317812 277458 317824
rect 278682 317812 278688 317824
rect 277452 317784 278688 317812
rect 277452 317772 277458 317784
rect 278682 317772 278688 317784
rect 278740 317772 278746 317824
rect 45462 317704 45468 317756
rect 45520 317744 45526 317756
rect 76742 317744 76748 317756
rect 45520 317716 76748 317744
rect 45520 317704 45526 317716
rect 76742 317704 76748 317716
rect 76800 317704 76806 317756
rect 99190 317704 99196 317756
rect 99248 317744 99254 317756
rect 100018 317744 100024 317756
rect 99248 317716 100024 317744
rect 99248 317704 99254 317716
rect 100018 317704 100024 317716
rect 100076 317704 100082 317756
rect 101030 317704 101036 317756
rect 101088 317744 101094 317756
rect 102778 317744 102784 317756
rect 101088 317716 102784 317744
rect 101088 317704 101094 317716
rect 102778 317704 102784 317716
rect 102836 317704 102842 317756
rect 106826 317704 106832 317756
rect 106884 317744 106890 317756
rect 107470 317744 107476 317756
rect 106884 317716 107476 317744
rect 106884 317704 106890 317716
rect 107470 317704 107476 317716
rect 107528 317704 107534 317756
rect 108206 317704 108212 317756
rect 108264 317744 108270 317756
rect 108942 317744 108948 317756
rect 108264 317716 108948 317744
rect 108264 317704 108270 317716
rect 108942 317704 108948 317716
rect 109000 317704 109006 317756
rect 125597 317747 125655 317753
rect 125597 317744 125609 317747
rect 118896 317716 125609 317744
rect 50982 317636 50988 317688
rect 51040 317676 51046 317688
rect 78950 317676 78956 317688
rect 51040 317648 78956 317676
rect 51040 317636 51046 317648
rect 78950 317636 78956 317648
rect 79008 317636 79014 317688
rect 100570 317636 100576 317688
rect 100628 317676 100634 317688
rect 104158 317676 104164 317688
rect 100628 317648 104164 317676
rect 100628 317636 100634 317648
rect 104158 317636 104164 317648
rect 104216 317636 104222 317688
rect 115937 317679 115995 317685
rect 115937 317645 115949 317679
rect 115983 317676 115995 317679
rect 118896 317676 118924 317716
rect 125597 317713 125609 317716
rect 125643 317713 125655 317747
rect 138569 317747 138627 317753
rect 125597 317707 125655 317713
rect 128372 317716 138520 317744
rect 115983 317648 118924 317676
rect 115983 317645 115995 317648
rect 115937 317639 115995 317645
rect 119430 317636 119436 317688
rect 119488 317676 119494 317688
rect 126977 317679 127035 317685
rect 126977 317676 126989 317679
rect 119488 317648 126989 317676
rect 119488 317636 119494 317648
rect 126977 317645 126989 317648
rect 127023 317645 127035 317679
rect 128372 317676 128400 317716
rect 126977 317639 127035 317645
rect 127084 317648 128400 317676
rect 46842 317568 46848 317620
rect 46900 317608 46906 317620
rect 77202 317608 77208 317620
rect 46900 317580 77208 317608
rect 46900 317568 46906 317580
rect 77202 317568 77208 317580
rect 77260 317568 77266 317620
rect 77938 317568 77944 317620
rect 77996 317608 78002 317620
rect 85298 317608 85304 317620
rect 77996 317580 85304 317608
rect 77996 317568 78002 317580
rect 85298 317568 85304 317580
rect 85356 317568 85362 317620
rect 91002 317568 91008 317620
rect 91060 317608 91066 317620
rect 94222 317608 94228 317620
rect 91060 317580 94228 317608
rect 91060 317568 91066 317580
rect 94222 317568 94228 317580
rect 94280 317568 94286 317620
rect 102318 317568 102324 317620
rect 102376 317608 102382 317620
rect 104250 317608 104256 317620
rect 102376 317580 104256 317608
rect 102376 317568 102382 317580
rect 104250 317568 104256 317580
rect 104308 317568 104314 317620
rect 106366 317568 106372 317620
rect 106424 317608 106430 317620
rect 107562 317608 107568 317620
rect 106424 317580 107568 317608
rect 106424 317568 106430 317580
rect 107562 317568 107568 317580
rect 107620 317568 107626 317620
rect 123478 317568 123484 317620
rect 123536 317608 123542 317620
rect 124122 317608 124128 317620
rect 123536 317580 124128 317608
rect 123536 317568 123542 317580
rect 124122 317568 124128 317580
rect 124180 317568 124186 317620
rect 125597 317611 125655 317617
rect 125597 317577 125609 317611
rect 125643 317608 125655 317611
rect 127084 317608 127112 317648
rect 131942 317636 131948 317688
rect 132000 317676 132006 317688
rect 138014 317676 138020 317688
rect 132000 317648 138020 317676
rect 132000 317636 132006 317648
rect 138014 317636 138020 317648
rect 138072 317636 138078 317688
rect 138492 317676 138520 317716
rect 138569 317713 138581 317747
rect 138615 317744 138627 317747
rect 147677 317747 147735 317753
rect 147677 317744 147689 317747
rect 138615 317716 147689 317744
rect 138615 317713 138627 317716
rect 138569 317707 138627 317713
rect 147677 317713 147689 317716
rect 147723 317713 147735 317747
rect 152274 317744 152280 317756
rect 147677 317707 147735 317713
rect 147784 317716 152280 317744
rect 140774 317676 140780 317688
rect 138492 317648 140780 317676
rect 140774 317636 140780 317648
rect 140832 317636 140838 317688
rect 140869 317679 140927 317685
rect 140869 317645 140881 317679
rect 140915 317676 140927 317679
rect 145558 317676 145564 317688
rect 140915 317648 145564 317676
rect 140915 317645 140927 317648
rect 140869 317639 140927 317645
rect 145558 317636 145564 317648
rect 145616 317636 145622 317688
rect 145653 317679 145711 317685
rect 145653 317645 145665 317679
rect 145699 317676 145711 317679
rect 147784 317676 147812 317716
rect 152274 317704 152280 317716
rect 152332 317704 152338 317756
rect 152461 317747 152519 317753
rect 152461 317713 152473 317747
rect 152507 317744 152519 317747
rect 159450 317744 159456 317756
rect 152507 317716 159456 317744
rect 152507 317713 152519 317716
rect 152461 317707 152519 317713
rect 159450 317704 159456 317716
rect 159508 317704 159514 317756
rect 160370 317744 160376 317756
rect 159560 317716 160376 317744
rect 145699 317648 147812 317676
rect 147861 317679 147919 317685
rect 145699 317645 145711 317648
rect 145653 317639 145711 317645
rect 147861 317645 147873 317679
rect 147907 317676 147919 317679
rect 152550 317676 152556 317688
rect 147907 317648 152556 317676
rect 147907 317645 147919 317648
rect 147861 317639 147919 317645
rect 152550 317636 152556 317648
rect 152608 317636 152614 317688
rect 152645 317679 152703 317685
rect 152645 317645 152657 317679
rect 152691 317676 152703 317679
rect 159560 317676 159588 317716
rect 160370 317704 160376 317716
rect 160428 317704 160434 317756
rect 162486 317704 162492 317756
rect 162544 317744 162550 317756
rect 180058 317744 180064 317756
rect 162544 317716 180064 317744
rect 162544 317704 162550 317716
rect 180058 317704 180064 317716
rect 180116 317704 180122 317756
rect 188062 317704 188068 317756
rect 188120 317744 188126 317756
rect 248509 317747 248567 317753
rect 248509 317744 248521 317747
rect 188120 317716 248521 317744
rect 188120 317704 188126 317716
rect 248509 317713 248521 317716
rect 248555 317713 248567 317747
rect 248509 317707 248567 317713
rect 248601 317747 248659 317753
rect 248601 317713 248613 317747
rect 248647 317744 248659 317747
rect 253290 317744 253296 317756
rect 248647 317716 253296 317744
rect 248647 317713 248659 317716
rect 248601 317707 248659 317713
rect 253290 317704 253296 317716
rect 253348 317704 253354 317756
rect 262582 317704 262588 317756
rect 262640 317744 262646 317756
rect 263502 317744 263508 317756
rect 262640 317716 263508 317744
rect 262640 317704 262646 317716
rect 263502 317704 263508 317716
rect 263560 317704 263566 317756
rect 152691 317648 159588 317676
rect 162121 317679 162179 317685
rect 152691 317645 152703 317648
rect 152645 317639 152703 317645
rect 162121 317645 162133 317679
rect 162167 317676 162179 317679
rect 171778 317676 171784 317688
rect 162167 317648 171784 317676
rect 162167 317645 162179 317648
rect 162121 317639 162179 317645
rect 171778 317636 171784 317648
rect 171836 317636 171842 317688
rect 182818 317676 182824 317688
rect 171888 317648 182824 317676
rect 135441 317611 135499 317617
rect 135441 317608 135453 317611
rect 125643 317580 127112 317608
rect 131132 317580 135453 317608
rect 125643 317577 125655 317580
rect 125597 317571 125655 317577
rect 53742 317500 53748 317552
rect 53800 317540 53806 317552
rect 79870 317540 79876 317552
rect 53800 317512 79876 317540
rect 53800 317500 53806 317512
rect 79870 317500 79876 317512
rect 79928 317500 79934 317552
rect 82170 317500 82176 317552
rect 82228 317540 82234 317552
rect 88886 317540 88892 317552
rect 82228 317512 88892 317540
rect 82228 317500 82234 317512
rect 88886 317500 88892 317512
rect 88944 317500 88950 317552
rect 92382 317500 92388 317552
rect 92440 317540 92446 317552
rect 94682 317540 94688 317552
rect 92440 317512 94688 317540
rect 92440 317500 92446 317512
rect 94682 317500 94688 317512
rect 94740 317500 94746 317552
rect 97442 317500 97448 317552
rect 97500 317540 97506 317552
rect 97902 317540 97908 317552
rect 97500 317512 97908 317540
rect 97500 317500 97506 317512
rect 97902 317500 97908 317512
rect 97960 317500 97966 317552
rect 109494 317500 109500 317552
rect 109552 317540 109558 317552
rect 110138 317540 110144 317552
rect 109552 317512 110144 317540
rect 109552 317500 109558 317512
rect 110138 317500 110144 317512
rect 110196 317500 110202 317552
rect 130378 317540 130384 317552
rect 128740 317512 130384 317540
rect 57882 317432 57888 317484
rect 57940 317472 57946 317484
rect 81710 317472 81716 317484
rect 57940 317444 81716 317472
rect 57940 317432 57946 317444
rect 81710 317432 81716 317444
rect 81768 317432 81774 317484
rect 86218 317432 86224 317484
rect 86276 317472 86282 317484
rect 88426 317472 88432 317484
rect 86276 317444 88432 317472
rect 86276 317432 86282 317444
rect 88426 317432 88432 317444
rect 88484 317432 88490 317484
rect 90358 317432 90364 317484
rect 90416 317472 90422 317484
rect 91094 317472 91100 317484
rect 90416 317444 91100 317472
rect 90416 317432 90422 317444
rect 91094 317432 91100 317444
rect 91152 317432 91158 317484
rect 93762 317432 93768 317484
rect 93820 317472 93826 317484
rect 95142 317472 95148 317484
rect 93820 317444 95148 317472
rect 93820 317432 93826 317444
rect 95142 317432 95148 317444
rect 95200 317432 95206 317484
rect 96982 317432 96988 317484
rect 97040 317472 97046 317484
rect 97718 317472 97724 317484
rect 97040 317444 97724 317472
rect 97040 317432 97046 317444
rect 97718 317432 97724 317444
rect 97776 317432 97782 317484
rect 103698 317432 103704 317484
rect 103756 317472 103762 317484
rect 104710 317472 104716 317484
rect 103756 317444 104716 317472
rect 103756 317432 103762 317444
rect 104710 317432 104716 317444
rect 104768 317432 104774 317484
rect 109034 317432 109040 317484
rect 109092 317472 109098 317484
rect 110322 317472 110328 317484
rect 109092 317444 110328 317472
rect 109092 317432 109098 317444
rect 110322 317432 110328 317444
rect 110380 317432 110386 317484
rect 110874 317432 110880 317484
rect 110932 317472 110938 317484
rect 111610 317472 111616 317484
rect 110932 317444 111616 317472
rect 110932 317432 110938 317444
rect 111610 317432 111616 317444
rect 111668 317432 111674 317484
rect 112254 317432 112260 317484
rect 112312 317472 112318 317484
rect 112990 317472 112996 317484
rect 112312 317444 112996 317472
rect 112312 317432 112318 317444
rect 112990 317432 112996 317444
rect 113048 317432 113054 317484
rect 113542 317432 113548 317484
rect 113600 317472 113606 317484
rect 114370 317472 114376 317484
rect 113600 317444 114376 317472
rect 113600 317432 113606 317444
rect 114370 317432 114376 317444
rect 114428 317432 114434 317484
rect 114922 317432 114928 317484
rect 114980 317472 114986 317484
rect 115842 317472 115848 317484
rect 114980 317444 115848 317472
rect 114980 317432 114986 317444
rect 115842 317432 115848 317444
rect 115900 317432 115906 317484
rect 116210 317432 116216 317484
rect 116268 317472 116274 317484
rect 116946 317472 116952 317484
rect 116268 317444 116952 317472
rect 116268 317432 116274 317444
rect 116946 317432 116952 317444
rect 117004 317432 117010 317484
rect 118970 317432 118976 317484
rect 119028 317472 119034 317484
rect 119890 317472 119896 317484
rect 119028 317444 119896 317472
rect 119028 317432 119034 317444
rect 119890 317432 119896 317444
rect 119948 317432 119954 317484
rect 120258 317432 120264 317484
rect 120316 317472 120322 317484
rect 121270 317472 121276 317484
rect 120316 317444 121276 317472
rect 120316 317432 120322 317444
rect 121270 317432 121276 317444
rect 121328 317432 121334 317484
rect 121638 317432 121644 317484
rect 121696 317472 121702 317484
rect 122650 317472 122656 317484
rect 121696 317444 122656 317472
rect 121696 317432 121702 317444
rect 122650 317432 122656 317444
rect 122708 317432 122714 317484
rect 123018 317432 123024 317484
rect 123076 317472 123082 317484
rect 123938 317472 123944 317484
rect 123076 317444 123944 317472
rect 123076 317432 123082 317444
rect 123938 317432 123944 317444
rect 123996 317432 124002 317484
rect 124306 317432 124312 317484
rect 124364 317472 124370 317484
rect 125410 317472 125416 317484
rect 124364 317444 125416 317472
rect 124364 317432 124370 317444
rect 125410 317432 125416 317444
rect 125468 317432 125474 317484
rect 125686 317432 125692 317484
rect 125744 317472 125750 317484
rect 126882 317472 126888 317484
rect 125744 317444 126888 317472
rect 125744 317432 125750 317444
rect 126882 317432 126888 317444
rect 126940 317432 126946 317484
rect 126977 317475 127035 317481
rect 126977 317441 126989 317475
rect 127023 317472 127035 317475
rect 128740 317472 128768 317512
rect 130378 317500 130384 317512
rect 130436 317500 130442 317552
rect 127023 317444 128768 317472
rect 127023 317441 127035 317444
rect 126977 317435 127035 317441
rect 128814 317432 128820 317484
rect 128872 317472 128878 317484
rect 129642 317472 129648 317484
rect 128872 317444 129648 317472
rect 128872 317432 128878 317444
rect 129642 317432 129648 317444
rect 129700 317432 129706 317484
rect 129734 317432 129740 317484
rect 129792 317472 129798 317484
rect 131022 317472 131028 317484
rect 129792 317444 131028 317472
rect 129792 317432 129798 317444
rect 131022 317432 131028 317444
rect 131080 317432 131086 317484
rect 126606 317364 126612 317416
rect 126664 317404 126670 317416
rect 131132 317404 131160 317580
rect 135441 317577 135453 317580
rect 135487 317577 135499 317611
rect 135441 317571 135499 317577
rect 137922 317568 137928 317620
rect 137980 317608 137986 317620
rect 147401 317611 147459 317617
rect 147401 317608 147413 317611
rect 137980 317580 147413 317608
rect 137980 317568 137986 317580
rect 147401 317577 147413 317580
rect 147447 317577 147459 317611
rect 147401 317571 147459 317577
rect 147493 317611 147551 317617
rect 147493 317577 147505 317611
rect 147539 317608 147551 317611
rect 148318 317608 148324 317620
rect 147539 317580 148324 317608
rect 147539 317577 147551 317580
rect 147493 317571 147551 317577
rect 148318 317568 148324 317580
rect 148376 317568 148382 317620
rect 148413 317611 148471 317617
rect 148413 317577 148425 317611
rect 148459 317608 148471 317611
rect 156598 317608 156604 317620
rect 148459 317580 156604 317608
rect 148459 317577 148471 317580
rect 148413 317571 148471 317577
rect 156598 317568 156604 317580
rect 156656 317568 156662 317620
rect 156690 317568 156696 317620
rect 156748 317608 156754 317620
rect 157058 317608 157064 317620
rect 156748 317580 157064 317608
rect 156748 317568 156754 317580
rect 157058 317568 157064 317580
rect 157116 317568 157122 317620
rect 157518 317568 157524 317620
rect 157576 317608 157582 317620
rect 158622 317608 158628 317620
rect 157576 317580 158628 317608
rect 157576 317568 157582 317580
rect 158622 317568 158628 317580
rect 158680 317568 158686 317620
rect 158898 317568 158904 317620
rect 158956 317608 158962 317620
rect 160002 317608 160008 317620
rect 158956 317580 160008 317608
rect 158956 317568 158962 317580
rect 160002 317568 160008 317580
rect 160060 317568 160066 317620
rect 166074 317568 166080 317620
rect 166132 317608 166138 317620
rect 166810 317608 166816 317620
rect 166132 317580 166816 317608
rect 166132 317568 166138 317580
rect 166810 317568 166816 317580
rect 166868 317568 166874 317620
rect 133322 317500 133328 317552
rect 133380 317540 133386 317552
rect 137833 317543 137891 317549
rect 133380 317512 137784 317540
rect 133380 317500 133386 317512
rect 131482 317432 131488 317484
rect 131540 317472 131546 317484
rect 132402 317472 132408 317484
rect 131540 317444 132408 317472
rect 131540 317432 131546 317444
rect 132402 317432 132408 317444
rect 132460 317432 132466 317484
rect 132862 317432 132868 317484
rect 132920 317472 132926 317484
rect 133782 317472 133788 317484
rect 132920 317444 133788 317472
rect 132920 317432 132926 317444
rect 133782 317432 133788 317444
rect 133840 317432 133846 317484
rect 137756 317472 137784 317512
rect 137833 317509 137845 317543
rect 137879 317540 137891 317543
rect 138109 317543 138167 317549
rect 138109 317540 138121 317543
rect 137879 317512 138121 317540
rect 137879 317509 137891 317512
rect 137833 317503 137891 317509
rect 138109 317509 138121 317512
rect 138155 317509 138167 317543
rect 138109 317503 138167 317509
rect 138290 317500 138296 317552
rect 138348 317540 138354 317552
rect 139302 317540 139308 317552
rect 138348 317512 139308 317540
rect 138348 317500 138354 317512
rect 139302 317500 139308 317512
rect 139360 317500 139366 317552
rect 140685 317543 140743 317549
rect 140685 317540 140697 317543
rect 139412 317512 140697 317540
rect 138569 317475 138627 317481
rect 138569 317472 138581 317475
rect 137756 317444 138581 317472
rect 138569 317441 138581 317444
rect 138615 317441 138627 317475
rect 138569 317435 138627 317441
rect 138658 317432 138664 317484
rect 138716 317472 138722 317484
rect 139210 317472 139216 317484
rect 138716 317444 139216 317472
rect 138716 317432 138722 317444
rect 139210 317432 139216 317444
rect 139268 317432 139274 317484
rect 139412 317472 139440 317512
rect 140685 317509 140697 317512
rect 140731 317509 140743 317543
rect 140685 317503 140743 317509
rect 142246 317500 142252 317552
rect 142304 317540 142310 317552
rect 143442 317540 143448 317552
rect 142304 317512 143448 317540
rect 142304 317500 142310 317512
rect 143442 317500 143448 317512
rect 143500 317500 143506 317552
rect 143537 317543 143595 317549
rect 143537 317509 143549 317543
rect 143583 317540 143595 317543
rect 147953 317543 148011 317549
rect 147953 317540 147965 317543
rect 143583 317512 147965 317540
rect 143583 317509 143595 317512
rect 143537 317503 143595 317509
rect 147953 317509 147965 317512
rect 147999 317509 148011 317543
rect 151078 317540 151084 317552
rect 147953 317503 148011 317509
rect 148060 317512 151084 317540
rect 139320 317444 139440 317472
rect 126664 317376 131160 317404
rect 126664 317364 126670 317376
rect 135898 317364 135904 317416
rect 135956 317404 135962 317416
rect 137833 317407 137891 317413
rect 137833 317404 137845 317407
rect 135956 317376 137845 317404
rect 135956 317364 135962 317376
rect 137833 317373 137845 317376
rect 137879 317373 137891 317407
rect 137833 317367 137891 317373
rect 135441 317339 135499 317345
rect 135441 317305 135453 317339
rect 135487 317336 135499 317339
rect 139320 317336 139348 317444
rect 140038 317432 140044 317484
rect 140096 317472 140102 317484
rect 140590 317472 140596 317484
rect 140096 317444 140596 317472
rect 140096 317432 140102 317444
rect 140590 317432 140596 317444
rect 140648 317432 140654 317484
rect 141418 317432 141424 317484
rect 141476 317472 141482 317484
rect 141970 317472 141976 317484
rect 141476 317444 141976 317472
rect 141476 317432 141482 317444
rect 141970 317432 141976 317444
rect 142028 317432 142034 317484
rect 142706 317432 142712 317484
rect 142764 317472 142770 317484
rect 143350 317472 143356 317484
rect 142764 317444 143356 317472
rect 142764 317432 142770 317444
rect 143350 317432 143356 317444
rect 143408 317432 143414 317484
rect 144086 317432 144092 317484
rect 144144 317472 144150 317484
rect 144730 317472 144736 317484
rect 144144 317444 144736 317472
rect 144144 317432 144150 317444
rect 144730 317432 144736 317444
rect 144788 317432 144794 317484
rect 145466 317432 145472 317484
rect 145524 317472 145530 317484
rect 146202 317472 146208 317484
rect 145524 317444 146208 317472
rect 145524 317432 145530 317444
rect 146202 317432 146208 317444
rect 146260 317432 146266 317484
rect 146294 317432 146300 317484
rect 146352 317472 146358 317484
rect 147490 317472 147496 317484
rect 146352 317444 147496 317472
rect 146352 317432 146358 317444
rect 147490 317432 147496 317444
rect 147548 317432 147554 317484
rect 147585 317475 147643 317481
rect 147585 317441 147597 317475
rect 147631 317472 147643 317475
rect 148060 317472 148088 317512
rect 151078 317500 151084 317512
rect 151136 317500 151142 317552
rect 151357 317543 151415 317549
rect 151357 317509 151369 317543
rect 151403 317540 151415 317543
rect 155313 317543 155371 317549
rect 155313 317540 155325 317543
rect 151403 317512 155325 317540
rect 151403 317509 151415 317512
rect 151357 317503 151415 317509
rect 155313 317509 155325 317512
rect 155359 317509 155371 317543
rect 155313 317503 155371 317509
rect 155405 317543 155463 317549
rect 155405 317509 155417 317543
rect 155451 317540 155463 317543
rect 155451 317512 156000 317540
rect 155451 317509 155463 317512
rect 155405 317503 155463 317509
rect 147631 317444 148088 317472
rect 147631 317441 147643 317444
rect 147585 317435 147643 317441
rect 148134 317432 148140 317484
rect 148192 317472 148198 317484
rect 148962 317472 148968 317484
rect 148192 317444 148968 317472
rect 148192 317432 148198 317444
rect 148962 317432 148968 317444
rect 149020 317432 149026 317484
rect 149514 317432 149520 317484
rect 149572 317472 149578 317484
rect 150158 317472 150164 317484
rect 149572 317444 150164 317472
rect 149572 317432 149578 317444
rect 150158 317432 150164 317444
rect 150216 317432 150222 317484
rect 150802 317432 150808 317484
rect 150860 317472 150866 317484
rect 151722 317472 151728 317484
rect 150860 317444 151728 317472
rect 150860 317432 150866 317444
rect 151722 317432 151728 317444
rect 151780 317432 151786 317484
rect 152182 317432 152188 317484
rect 152240 317472 152246 317484
rect 153102 317472 153108 317484
rect 152240 317444 153108 317472
rect 152240 317432 152246 317444
rect 153102 317432 153108 317444
rect 153160 317432 153166 317484
rect 153470 317432 153476 317484
rect 153528 317472 153534 317484
rect 154482 317472 154488 317484
rect 153528 317444 154488 317472
rect 153528 317432 153534 317444
rect 154482 317432 154488 317444
rect 154540 317432 154546 317484
rect 154850 317432 154856 317484
rect 154908 317472 154914 317484
rect 155862 317472 155868 317484
rect 154908 317444 155868 317472
rect 154908 317432 154914 317444
rect 155862 317432 155868 317444
rect 155920 317432 155926 317484
rect 155972 317472 156000 317512
rect 156230 317500 156236 317552
rect 156288 317540 156294 317552
rect 157242 317540 157248 317552
rect 156288 317512 157248 317540
rect 156288 317500 156294 317512
rect 157242 317500 157248 317512
rect 157300 317500 157306 317552
rect 157904 317512 159312 317540
rect 157904 317472 157932 317512
rect 155972 317444 157932 317472
rect 157978 317432 157984 317484
rect 158036 317472 158042 317484
rect 158530 317472 158536 317484
rect 158036 317444 158536 317472
rect 158036 317432 158042 317444
rect 158530 317432 158536 317444
rect 158588 317432 158594 317484
rect 147401 317407 147459 317413
rect 147401 317373 147413 317407
rect 147447 317404 147459 317407
rect 147861 317407 147919 317413
rect 147861 317404 147873 317407
rect 147447 317376 147873 317404
rect 147447 317373 147459 317376
rect 147401 317367 147459 317373
rect 147861 317373 147873 317376
rect 147907 317373 147919 317407
rect 159284 317404 159312 317512
rect 160278 317500 160284 317552
rect 160336 317540 160342 317552
rect 161382 317540 161388 317552
rect 160336 317512 161388 317540
rect 160336 317500 160342 317512
rect 161382 317500 161388 317512
rect 161440 317500 161446 317552
rect 162026 317500 162032 317552
rect 162084 317540 162090 317552
rect 162670 317540 162676 317552
rect 162084 317512 162676 317540
rect 162084 317500 162090 317512
rect 162670 317500 162676 317512
rect 162728 317500 162734 317552
rect 163406 317500 163412 317552
rect 163464 317540 163470 317552
rect 164050 317540 164056 317552
rect 163464 317512 164056 317540
rect 163464 317500 163470 317512
rect 164050 317500 164056 317512
rect 164108 317500 164114 317552
rect 164326 317500 164332 317552
rect 164384 317540 164390 317552
rect 165522 317540 165528 317552
rect 164384 317512 165528 317540
rect 164384 317500 164390 317512
rect 165522 317500 165528 317512
rect 165580 317500 165586 317552
rect 166534 317500 166540 317552
rect 166592 317540 166598 317552
rect 171888 317540 171916 317648
rect 182818 317636 182824 317648
rect 182876 317636 182882 317688
rect 189074 317636 189080 317688
rect 189132 317676 189138 317688
rect 189810 317676 189816 317688
rect 189132 317648 189816 317676
rect 189132 317636 189138 317648
rect 189810 317636 189816 317648
rect 189868 317636 189874 317688
rect 190730 317636 190736 317688
rect 190788 317676 190794 317688
rect 191742 317676 191748 317688
rect 190788 317648 191748 317676
rect 190788 317636 190794 317648
rect 191742 317636 191748 317648
rect 191800 317636 191806 317688
rect 204714 317636 204720 317688
rect 204772 317676 204778 317688
rect 205542 317676 205548 317688
rect 204772 317648 205548 317676
rect 204772 317636 204778 317648
rect 205542 317636 205548 317648
rect 205600 317636 205606 317688
rect 271230 317676 271236 317688
rect 209700 317648 271236 317676
rect 182726 317568 182732 317620
rect 182784 317608 182790 317620
rect 189905 317611 189963 317617
rect 189905 317608 189917 317611
rect 182784 317580 189917 317608
rect 182784 317568 182790 317580
rect 189905 317577 189917 317580
rect 189951 317577 189963 317611
rect 189905 317571 189963 317577
rect 166592 317512 171916 317540
rect 166592 317500 166598 317512
rect 204254 317500 204260 317552
rect 204312 317540 204318 317552
rect 209700 317540 209728 317648
rect 271230 317636 271236 317648
rect 271288 317636 271294 317688
rect 218606 317568 218612 317620
rect 218664 317608 218670 317620
rect 219250 317608 219256 317620
rect 218664 317580 219256 317608
rect 218664 317568 218670 317580
rect 219250 317568 219256 317580
rect 219308 317568 219314 317620
rect 219526 317568 219532 317620
rect 219584 317608 219590 317620
rect 220722 317608 220728 317620
rect 219584 317580 220728 317608
rect 219584 317568 219590 317580
rect 220722 317568 220728 317580
rect 220780 317568 220786 317620
rect 221274 317568 221280 317620
rect 221332 317608 221338 317620
rect 221918 317608 221924 317620
rect 221332 317580 221924 317608
rect 221332 317568 221338 317580
rect 221918 317568 221924 317580
rect 221976 317568 221982 317620
rect 222194 317568 222200 317620
rect 222252 317608 222258 317620
rect 223482 317608 223488 317620
rect 222252 317580 223488 317608
rect 222252 317568 222258 317580
rect 223482 317568 223488 317580
rect 223540 317568 223546 317620
rect 224402 317568 224408 317620
rect 224460 317608 224466 317620
rect 229005 317611 229063 317617
rect 229005 317608 229017 317611
rect 224460 317580 229017 317608
rect 224460 317568 224466 317580
rect 229005 317577 229017 317580
rect 229051 317577 229063 317611
rect 229005 317571 229063 317577
rect 229370 317568 229376 317620
rect 229428 317608 229434 317620
rect 230198 317608 230204 317620
rect 229428 317580 230204 317608
rect 229428 317568 229434 317580
rect 230198 317568 230204 317580
rect 230256 317568 230262 317620
rect 230750 317568 230756 317620
rect 230808 317608 230814 317620
rect 231670 317608 231676 317620
rect 230808 317580 231676 317608
rect 230808 317568 230814 317580
rect 231670 317568 231676 317580
rect 231728 317568 231734 317620
rect 232038 317568 232044 317620
rect 232096 317608 232102 317620
rect 232958 317608 232964 317620
rect 232096 317580 232964 317608
rect 232096 317568 232102 317580
rect 232958 317568 232964 317580
rect 233016 317568 233022 317620
rect 233418 317568 233424 317620
rect 233476 317608 233482 317620
rect 234430 317608 234436 317620
rect 233476 317580 234436 317608
rect 233476 317568 233482 317580
rect 234430 317568 234436 317580
rect 234488 317568 234494 317620
rect 234798 317568 234804 317620
rect 234856 317608 234862 317620
rect 235718 317608 235724 317620
rect 234856 317580 235724 317608
rect 234856 317568 234862 317580
rect 235718 317568 235724 317580
rect 235776 317568 235782 317620
rect 236086 317568 236092 317620
rect 236144 317608 236150 317620
rect 237190 317608 237196 317620
rect 236144 317580 237196 317608
rect 236144 317568 236150 317580
rect 237190 317568 237196 317580
rect 237248 317568 237254 317620
rect 237466 317568 237472 317620
rect 237524 317608 237530 317620
rect 238478 317608 238484 317620
rect 237524 317580 238484 317608
rect 237524 317568 237530 317580
rect 238478 317568 238484 317580
rect 238536 317568 238542 317620
rect 238846 317568 238852 317620
rect 238904 317608 238910 317620
rect 239950 317608 239956 317620
rect 238904 317580 239956 317608
rect 238904 317568 238910 317580
rect 239950 317568 239956 317580
rect 240008 317568 240014 317620
rect 240134 317568 240140 317620
rect 240192 317608 240198 317620
rect 241238 317608 241244 317620
rect 240192 317580 241244 317608
rect 240192 317568 240198 317580
rect 241238 317568 241244 317580
rect 241296 317568 241302 317620
rect 241974 317568 241980 317620
rect 242032 317608 242038 317620
rect 242618 317608 242624 317620
rect 242032 317580 242624 317608
rect 242032 317568 242038 317580
rect 242618 317568 242624 317580
rect 242676 317568 242682 317620
rect 243262 317568 243268 317620
rect 243320 317608 243326 317620
rect 244182 317608 244188 317620
rect 243320 317580 244188 317608
rect 243320 317568 243326 317580
rect 244182 317568 244188 317580
rect 244240 317568 244246 317620
rect 246022 317568 246028 317620
rect 246080 317608 246086 317620
rect 246942 317608 246948 317620
rect 246080 317580 246948 317608
rect 246080 317568 246086 317580
rect 246942 317568 246948 317580
rect 247000 317568 247006 317620
rect 247310 317568 247316 317620
rect 247368 317608 247374 317620
rect 248230 317608 248236 317620
rect 247368 317580 248236 317608
rect 247368 317568 247374 317580
rect 248230 317568 248236 317580
rect 248288 317568 248294 317620
rect 248509 317611 248567 317617
rect 248509 317577 248521 317611
rect 248555 317608 248567 317611
rect 255958 317608 255964 317620
rect 248555 317580 255964 317608
rect 248555 317577 248567 317580
rect 248509 317571 248567 317577
rect 255958 317568 255964 317580
rect 256016 317568 256022 317620
rect 204312 317512 209728 317540
rect 204312 317500 204318 317512
rect 224034 317500 224040 317552
rect 224092 317540 224098 317552
rect 224678 317540 224684 317552
rect 224092 317512 224684 317540
rect 224092 317500 224098 317512
rect 224678 317500 224684 317512
rect 224736 317500 224742 317552
rect 229830 317500 229836 317552
rect 229888 317540 229894 317552
rect 230382 317540 230388 317552
rect 229888 317512 230388 317540
rect 229888 317500 229894 317512
rect 230382 317500 230388 317512
rect 230440 317500 230446 317552
rect 232498 317500 232504 317552
rect 232556 317540 232562 317552
rect 233142 317540 233148 317552
rect 232556 317512 233148 317540
rect 232556 317500 232562 317512
rect 233142 317500 233148 317512
rect 233200 317500 233206 317552
rect 235258 317500 235264 317552
rect 235316 317540 235322 317552
rect 235902 317540 235908 317552
rect 235316 317512 235908 317540
rect 235316 317500 235322 317512
rect 235902 317500 235908 317512
rect 235960 317500 235966 317552
rect 236546 317500 236552 317552
rect 236604 317540 236610 317552
rect 237098 317540 237104 317552
rect 236604 317512 237104 317540
rect 236604 317500 236610 317512
rect 237098 317500 237104 317512
rect 237156 317500 237162 317552
rect 237926 317500 237932 317552
rect 237984 317540 237990 317552
rect 238662 317540 238668 317552
rect 237984 317512 238668 317540
rect 237984 317500 237990 317512
rect 238662 317500 238668 317512
rect 238720 317500 238726 317552
rect 239214 317500 239220 317552
rect 239272 317540 239278 317552
rect 239858 317540 239864 317552
rect 239272 317512 239864 317540
rect 239272 317500 239278 317512
rect 239858 317500 239864 317512
rect 239916 317500 239922 317552
rect 240594 317500 240600 317552
rect 240652 317540 240658 317552
rect 241422 317540 241428 317552
rect 240652 317512 241428 317540
rect 240652 317500 240658 317512
rect 241422 317500 241428 317512
rect 241480 317500 241486 317552
rect 241514 317500 241520 317552
rect 241572 317540 241578 317552
rect 242710 317540 242716 317552
rect 241572 317512 242716 317540
rect 241572 317500 241578 317512
rect 242710 317500 242716 317512
rect 242768 317500 242774 317552
rect 244642 317500 244648 317552
rect 244700 317540 244706 317552
rect 245562 317540 245568 317552
rect 244700 317512 245568 317540
rect 244700 317500 244706 317512
rect 245562 317500 245568 317512
rect 245620 317500 245626 317552
rect 259454 317500 259460 317552
rect 259512 317540 259518 317552
rect 260558 317540 260564 317552
rect 259512 317512 260564 317540
rect 259512 317500 259518 317512
rect 260558 317500 260564 317512
rect 260616 317500 260622 317552
rect 159358 317432 159364 317484
rect 159416 317472 159422 317484
rect 159910 317472 159916 317484
rect 159416 317444 159916 317472
rect 159416 317432 159422 317444
rect 159910 317432 159916 317444
rect 159968 317432 159974 317484
rect 160738 317432 160744 317484
rect 160796 317472 160802 317484
rect 161290 317472 161296 317484
rect 160796 317444 161296 317472
rect 160796 317432 160802 317444
rect 161290 317432 161296 317444
rect 161348 317432 161354 317484
rect 161566 317432 161572 317484
rect 161624 317472 161630 317484
rect 162762 317472 162768 317484
rect 161624 317444 162768 317472
rect 161624 317432 161630 317444
rect 162762 317432 162768 317444
rect 162820 317432 162826 317484
rect 162946 317432 162952 317484
rect 163004 317472 163010 317484
rect 164142 317472 164148 317484
rect 163004 317444 164148 317472
rect 163004 317432 163010 317444
rect 164142 317432 164148 317444
rect 164200 317432 164206 317484
rect 164694 317432 164700 317484
rect 164752 317472 164758 317484
rect 165430 317472 165436 317484
rect 164752 317444 165436 317472
rect 164752 317432 164758 317444
rect 165430 317432 165436 317444
rect 165488 317432 165494 317484
rect 165614 317432 165620 317484
rect 165672 317472 165678 317484
rect 166902 317472 166908 317484
rect 165672 317444 166908 317472
rect 165672 317432 165678 317444
rect 166902 317432 166908 317444
rect 166960 317432 166966 317484
rect 171502 317432 171508 317484
rect 171560 317472 171566 317484
rect 172330 317472 172336 317484
rect 171560 317444 172336 317472
rect 171560 317432 171566 317444
rect 172330 317432 172336 317444
rect 172388 317432 172394 317484
rect 175550 317432 175556 317484
rect 175608 317472 175614 317484
rect 176470 317472 176476 317484
rect 175608 317444 176476 317472
rect 175608 317432 175614 317444
rect 176470 317432 176476 317444
rect 176528 317432 176534 317484
rect 179966 317432 179972 317484
rect 180024 317472 180030 317484
rect 180518 317472 180524 317484
rect 180024 317444 180524 317472
rect 180024 317432 180030 317444
rect 180518 317432 180524 317444
rect 180576 317432 180582 317484
rect 197998 317432 198004 317484
rect 198056 317472 198062 317484
rect 198642 317472 198648 317484
rect 198056 317444 198648 317472
rect 198056 317432 198062 317444
rect 198642 317432 198648 317444
rect 198700 317432 198706 317484
rect 201954 317432 201960 317484
rect 202012 317472 202018 317484
rect 202782 317472 202788 317484
rect 202012 317444 202788 317472
rect 202012 317432 202018 317444
rect 202782 317432 202788 317444
rect 202840 317432 202846 317484
rect 159284 317376 159404 317404
rect 147861 317367 147919 317373
rect 159376 317348 159404 317376
rect 135487 317308 139348 317336
rect 135487 317305 135499 317308
rect 135441 317299 135499 317305
rect 159358 317296 159364 317348
rect 159416 317296 159422 317348
rect 60734 315936 60740 315988
rect 60792 315976 60798 315988
rect 61102 315976 61108 315988
rect 60792 315948 61108 315976
rect 60792 315936 60798 315948
rect 61102 315936 61108 315948
rect 61160 315936 61166 315988
rect 64874 315936 64880 315988
rect 64932 315976 64938 315988
rect 65702 315976 65708 315988
rect 64932 315948 65708 315976
rect 64932 315936 64938 315948
rect 65702 315936 65708 315948
rect 65760 315936 65766 315988
rect 69106 315936 69112 315988
rect 69164 315976 69170 315988
rect 69382 315976 69388 315988
rect 69164 315948 69388 315976
rect 69164 315936 69170 315948
rect 69382 315936 69388 315948
rect 69440 315936 69446 315988
rect 80146 315936 80152 315988
rect 80204 315976 80210 315988
rect 80974 315976 80980 315988
rect 80204 315948 80980 315976
rect 80204 315936 80210 315948
rect 80974 315936 80980 315948
rect 81032 315936 81038 315988
rect 81526 315936 81532 315988
rect 81584 315976 81590 315988
rect 82262 315976 82268 315988
rect 81584 315948 82268 315976
rect 81584 315936 81590 315948
rect 82262 315936 82268 315948
rect 82320 315936 82326 315988
rect 84286 315936 84292 315988
rect 84344 315976 84350 315988
rect 84470 315976 84476 315988
rect 84344 315948 84476 315976
rect 84344 315936 84350 315948
rect 84470 315936 84476 315948
rect 84528 315936 84534 315988
rect 85574 315936 85580 315988
rect 85632 315976 85638 315988
rect 86310 315976 86316 315988
rect 85632 315948 86316 315976
rect 85632 315936 85638 315948
rect 86310 315936 86316 315948
rect 86368 315936 86374 315988
rect 92566 315936 92572 315988
rect 92624 315976 92630 315988
rect 93486 315976 93492 315988
rect 92624 315948 93492 315976
rect 92624 315936 92630 315948
rect 93486 315936 93492 315948
rect 93544 315936 93550 315988
rect 74994 315868 75000 315920
rect 75052 315908 75058 315920
rect 75454 315908 75460 315920
rect 75052 315880 75460 315908
rect 75052 315868 75058 315880
rect 75454 315868 75460 315880
rect 75512 315868 75518 315920
rect 77570 315868 77576 315920
rect 77628 315908 77634 315920
rect 78214 315908 78220 315920
rect 77628 315880 78220 315908
rect 77628 315868 77634 315880
rect 78214 315868 78220 315880
rect 78272 315868 78278 315920
rect 117866 315868 117872 315920
rect 117924 315908 117930 315920
rect 118510 315908 118516 315920
rect 117924 315880 118516 315908
rect 117924 315868 117930 315880
rect 118510 315868 118516 315880
rect 118568 315868 118574 315920
rect 82906 315664 82912 315716
rect 82964 315704 82970 315716
rect 83550 315704 83556 315716
rect 82964 315676 83556 315704
rect 82964 315664 82970 315676
rect 83550 315664 83556 315676
rect 83608 315664 83614 315716
rect 128354 315392 128360 315444
rect 128412 315432 128418 315444
rect 129550 315432 129556 315444
rect 128412 315404 129556 315432
rect 128412 315392 128418 315404
rect 129550 315392 129556 315404
rect 129608 315392 129614 315444
rect 66806 313896 66812 313948
rect 66864 313936 66870 313948
rect 66990 313936 66996 313948
rect 66864 313908 66996 313936
rect 66864 313896 66870 313908
rect 66990 313896 66996 313908
rect 67048 313896 67054 313948
rect 135073 311967 135131 311973
rect 135073 311933 135085 311967
rect 135119 311964 135131 311967
rect 135162 311964 135168 311976
rect 135119 311936 135168 311964
rect 135119 311933 135131 311936
rect 135073 311927 135131 311933
rect 135162 311924 135168 311936
rect 135220 311924 135226 311976
rect 137738 311856 137744 311908
rect 137796 311896 137802 311908
rect 137922 311896 137928 311908
rect 137796 311868 137928 311896
rect 137796 311856 137802 311868
rect 137922 311856 137928 311868
rect 137980 311856 137986 311908
rect 140774 311788 140780 311840
rect 140832 311828 140838 311840
rect 140958 311828 140964 311840
rect 140832 311800 140964 311828
rect 140832 311788 140838 311800
rect 140958 311788 140964 311800
rect 141016 311788 141022 311840
rect 78858 309136 78864 309188
rect 78916 309176 78922 309188
rect 79042 309176 79048 309188
rect 78916 309148 79048 309176
rect 78916 309136 78922 309148
rect 79042 309136 79048 309148
rect 79100 309136 79106 309188
rect 86034 309136 86040 309188
rect 86092 309176 86098 309188
rect 86126 309176 86132 309188
rect 86092 309148 86132 309176
rect 86092 309136 86098 309148
rect 86126 309136 86132 309148
rect 86184 309136 86190 309188
rect 135070 309176 135076 309188
rect 135031 309148 135076 309176
rect 135070 309136 135076 309148
rect 135128 309136 135134 309188
rect 160738 309176 160744 309188
rect 160699 309148 160744 309176
rect 160738 309136 160744 309148
rect 160796 309136 160802 309188
rect 66809 309111 66867 309117
rect 66809 309077 66821 309111
rect 66855 309108 66867 309111
rect 66990 309108 66996 309120
rect 66855 309080 66996 309108
rect 66855 309077 66867 309080
rect 66809 309071 66867 309077
rect 66990 309068 66996 309080
rect 67048 309068 67054 309120
rect 74442 309108 74448 309120
rect 74403 309080 74448 309108
rect 74442 309068 74448 309080
rect 74500 309068 74506 309120
rect 77570 309108 77576 309120
rect 77531 309080 77576 309108
rect 77570 309068 77576 309080
rect 77628 309068 77634 309120
rect 95418 309108 95424 309120
rect 95379 309080 95424 309108
rect 95418 309068 95424 309080
rect 95476 309068 95482 309120
rect 124401 307887 124459 307893
rect 124401 307853 124413 307887
rect 124447 307884 124459 307887
rect 124490 307884 124496 307896
rect 124447 307856 124496 307884
rect 124447 307853 124459 307856
rect 124401 307847 124459 307853
rect 124490 307844 124496 307856
rect 124548 307844 124554 307896
rect 85945 307751 86003 307757
rect 85945 307717 85957 307751
rect 85991 307748 86003 307751
rect 86034 307748 86040 307760
rect 85991 307720 86040 307748
rect 85991 307717 86003 307720
rect 85945 307711 86003 307717
rect 86034 307708 86040 307720
rect 86092 307708 86098 307760
rect 124217 307751 124275 307757
rect 124217 307717 124229 307751
rect 124263 307748 124275 307751
rect 124398 307748 124404 307760
rect 124263 307720 124404 307748
rect 124263 307717 124275 307720
rect 124217 307711 124275 307717
rect 124398 307708 124404 307720
rect 124456 307708 124462 307760
rect 136634 307028 136640 307080
rect 136692 307068 136698 307080
rect 137922 307068 137928 307080
rect 136692 307040 137928 307068
rect 136692 307028 136698 307040
rect 137922 307028 137928 307040
rect 137980 307028 137986 307080
rect 139394 307028 139400 307080
rect 139452 307068 139458 307080
rect 140682 307068 140688 307080
rect 139452 307040 140688 307068
rect 139452 307028 139458 307040
rect 140682 307028 140688 307040
rect 140740 307028 140746 307080
rect 140866 307028 140872 307080
rect 140924 307068 140930 307080
rect 142062 307068 142068 307080
rect 140924 307040 142068 307068
rect 140924 307028 140930 307040
rect 142062 307028 142068 307040
rect 142120 307028 142126 307080
rect 143626 307028 143632 307080
rect 143684 307068 143690 307080
rect 144822 307068 144828 307080
rect 143684 307040 144828 307068
rect 143684 307028 143690 307040
rect 144822 307028 144828 307040
rect 144880 307028 144886 307080
rect 74994 302376 75000 302388
rect 74955 302348 75000 302376
rect 74994 302336 75000 302348
rect 75052 302336 75058 302388
rect 134978 302240 134984 302252
rect 134939 302212 134984 302240
rect 134978 302200 134984 302212
rect 135036 302200 135042 302252
rect 80241 301563 80299 301569
rect 80241 301529 80253 301563
rect 80287 301560 80299 301563
rect 80422 301560 80428 301572
rect 80287 301532 80428 301560
rect 80287 301529 80299 301532
rect 80241 301523 80299 301529
rect 80422 301520 80428 301532
rect 80480 301520 80486 301572
rect 66806 299520 66812 299532
rect 66767 299492 66812 299520
rect 66806 299480 66812 299492
rect 66864 299480 66870 299532
rect 74442 299520 74448 299532
rect 74403 299492 74448 299520
rect 74442 299480 74448 299492
rect 74500 299480 74506 299532
rect 74994 299520 75000 299532
rect 74955 299492 75000 299520
rect 74994 299480 75000 299492
rect 75052 299480 75058 299532
rect 77570 299520 77576 299532
rect 77531 299492 77576 299520
rect 77570 299480 77576 299492
rect 77628 299480 77634 299532
rect 95421 299523 95479 299529
rect 95421 299489 95433 299523
rect 95467 299520 95479 299523
rect 95694 299520 95700 299532
rect 95467 299492 95700 299520
rect 95467 299489 95479 299492
rect 95421 299483 95479 299489
rect 95694 299480 95700 299492
rect 95752 299480 95758 299532
rect 134978 299520 134984 299532
rect 134939 299492 134984 299520
rect 134978 299480 134984 299492
rect 135036 299480 135042 299532
rect 74905 299387 74963 299393
rect 74905 299353 74917 299387
rect 74951 299384 74963 299387
rect 74994 299384 75000 299396
rect 74951 299356 75000 299384
rect 74951 299353 74963 299356
rect 74905 299347 74963 299353
rect 74994 299344 75000 299356
rect 75052 299344 75058 299396
rect 124214 298188 124220 298240
rect 124272 298228 124278 298240
rect 124272 298200 124317 298228
rect 124272 298188 124278 298200
rect 85942 298160 85948 298172
rect 85903 298132 85948 298160
rect 85942 298120 85948 298132
rect 86000 298120 86006 298172
rect 74442 298092 74448 298104
rect 74403 298064 74448 298092
rect 74442 298052 74448 298064
rect 74500 298052 74506 298104
rect 124214 298052 124220 298104
rect 124272 298092 124278 298104
rect 124401 298095 124459 298101
rect 124401 298092 124413 298095
rect 124272 298064 124413 298092
rect 124272 298052 124278 298064
rect 124401 298061 124413 298064
rect 124447 298061 124459 298095
rect 124401 298055 124459 298061
rect 80238 296732 80244 296744
rect 80199 296704 80244 296732
rect 80238 296692 80244 296704
rect 80296 296692 80302 296744
rect 140774 296692 140780 296744
rect 140832 296732 140838 296744
rect 140958 296732 140964 296744
rect 140832 296704 140964 296732
rect 140832 296692 140838 296704
rect 140958 296692 140964 296704
rect 141016 296692 141022 296744
rect 66622 294584 66628 294636
rect 66680 294624 66686 294636
rect 66806 294624 66812 294636
rect 66680 294596 66812 294624
rect 66680 294584 66686 294596
rect 66806 294584 66812 294596
rect 66864 294584 66870 294636
rect 72237 292655 72295 292661
rect 72237 292621 72249 292655
rect 72283 292652 72295 292655
rect 72326 292652 72332 292664
rect 72283 292624 72332 292652
rect 72283 292621 72295 292624
rect 72237 292615 72295 292621
rect 72326 292612 72332 292624
rect 72384 292612 72390 292664
rect 85942 292612 85948 292664
rect 86000 292612 86006 292664
rect 85960 292528 85988 292612
rect 85942 292476 85948 292528
rect 86000 292476 86006 292528
rect 124398 292448 124404 292460
rect 124359 292420 124404 292448
rect 124398 292408 124404 292420
rect 124456 292408 124462 292460
rect 72234 289864 72240 289876
rect 72195 289836 72240 289864
rect 72234 289824 72240 289836
rect 72292 289824 72298 289876
rect 74902 289864 74908 289876
rect 74863 289836 74908 289864
rect 74902 289824 74908 289836
rect 74960 289824 74966 289876
rect 134889 289799 134947 289805
rect 134889 289765 134901 289799
rect 134935 289796 134947 289799
rect 135162 289796 135168 289808
rect 134935 289768 135168 289796
rect 134935 289765 134947 289768
rect 134889 289759 134947 289765
rect 135162 289756 135168 289768
rect 135220 289756 135226 289808
rect 74902 289728 74908 289740
rect 74863 289700 74908 289728
rect 74902 289688 74908 289700
rect 74960 289688 74966 289740
rect 80238 288260 80244 288312
rect 80296 288260 80302 288312
rect 80256 288232 80284 288260
rect 80422 288232 80428 288244
rect 80256 288204 80428 288232
rect 80422 288192 80428 288204
rect 80480 288192 80486 288244
rect 81710 283608 81716 283620
rect 81671 283580 81716 283608
rect 81710 283568 81716 283580
rect 81768 283568 81774 283620
rect 124398 282956 124404 283008
rect 124456 282956 124462 283008
rect 77570 282928 77576 282940
rect 77531 282900 77576 282928
rect 77570 282888 77576 282900
rect 77628 282888 77634 282940
rect 124416 282872 124444 282956
rect 150158 282888 150164 282940
rect 150216 282928 150222 282940
rect 150342 282928 150348 282940
rect 150216 282900 150348 282928
rect 150216 282888 150222 282900
rect 150342 282888 150348 282900
rect 150400 282888 150406 282940
rect 124398 282820 124404 282872
rect 124456 282820 124462 282872
rect 74442 280208 74448 280220
rect 74403 280180 74448 280208
rect 74442 280168 74448 280180
rect 74500 280168 74506 280220
rect 74905 280211 74963 280217
rect 74905 280177 74917 280211
rect 74951 280208 74963 280211
rect 74994 280208 75000 280220
rect 74951 280180 75000 280208
rect 74951 280177 74963 280180
rect 74905 280171 74963 280177
rect 74994 280168 75000 280180
rect 75052 280168 75058 280220
rect 134886 280208 134892 280220
rect 134847 280180 134892 280208
rect 134886 280168 134892 280180
rect 134944 280168 134950 280220
rect 66530 280140 66536 280152
rect 66491 280112 66536 280140
rect 66530 280100 66536 280112
rect 66588 280100 66594 280152
rect 72234 280140 72240 280152
rect 72195 280112 72240 280140
rect 72234 280100 72240 280112
rect 72292 280100 72298 280152
rect 95602 280140 95608 280152
rect 95563 280112 95608 280140
rect 95602 280100 95608 280112
rect 95660 280100 95666 280152
rect 124398 280140 124404 280152
rect 124359 280112 124404 280140
rect 124398 280100 124404 280112
rect 124456 280100 124462 280152
rect 85850 278808 85856 278860
rect 85908 278848 85914 278860
rect 85942 278848 85948 278860
rect 85908 278820 85948 278848
rect 85908 278808 85914 278820
rect 85942 278808 85948 278820
rect 86000 278808 86006 278860
rect 81710 278780 81716 278792
rect 81671 278752 81716 278780
rect 81710 278740 81716 278752
rect 81768 278740 81774 278792
rect 85850 278672 85856 278724
rect 85908 278712 85914 278724
rect 86034 278712 86040 278724
rect 85908 278684 86040 278712
rect 85908 278672 85914 278684
rect 86034 278672 86040 278684
rect 86092 278672 86098 278724
rect 86034 277312 86040 277364
rect 86092 277352 86098 277364
rect 86126 277352 86132 277364
rect 86092 277324 86132 277352
rect 86092 277312 86098 277324
rect 86126 277312 86132 277324
rect 86184 277312 86190 277364
rect 124398 273952 124404 273964
rect 124359 273924 124404 273952
rect 124398 273912 124404 273924
rect 124456 273912 124462 273964
rect 66533 270555 66591 270561
rect 66533 270521 66545 270555
rect 66579 270552 66591 270555
rect 66622 270552 66628 270564
rect 66579 270524 66628 270552
rect 66579 270521 66591 270524
rect 66533 270515 66591 270521
rect 66622 270512 66628 270524
rect 66680 270512 66686 270564
rect 72234 270552 72240 270564
rect 72195 270524 72240 270552
rect 72234 270512 72240 270524
rect 72292 270512 72298 270564
rect 77570 270552 77576 270564
rect 77531 270524 77576 270552
rect 77570 270512 77576 270524
rect 77628 270512 77634 270564
rect 95605 270555 95663 270561
rect 95605 270521 95617 270555
rect 95651 270552 95663 270555
rect 95694 270552 95700 270564
rect 95651 270524 95700 270552
rect 95651 270521 95663 270524
rect 95605 270515 95663 270521
rect 95694 270512 95700 270524
rect 95752 270512 95758 270564
rect 134889 270487 134947 270493
rect 134889 270453 134901 270487
rect 134935 270484 134947 270487
rect 134978 270484 134984 270496
rect 134935 270456 134984 270484
rect 134935 270453 134947 270456
rect 134889 270447 134947 270453
rect 134978 270444 134984 270456
rect 135036 270444 135042 270496
rect 74258 269084 74264 269136
rect 74316 269124 74322 269136
rect 74442 269124 74448 269136
rect 74316 269096 74448 269124
rect 74316 269084 74322 269096
rect 74442 269084 74448 269096
rect 74500 269084 74506 269136
rect 124306 263616 124312 263628
rect 124267 263588 124312 263616
rect 124306 263576 124312 263588
rect 124364 263576 124370 263628
rect 140774 263576 140780 263628
rect 140832 263616 140838 263628
rect 140958 263616 140964 263628
rect 140832 263588 140964 263616
rect 140832 263576 140838 263588
rect 140958 263576 140964 263588
rect 141016 263576 141022 263628
rect 150158 263576 150164 263628
rect 150216 263616 150222 263628
rect 150342 263616 150348 263628
rect 150216 263588 150348 263616
rect 150216 263576 150222 263588
rect 150342 263576 150348 263588
rect 150400 263576 150406 263628
rect 134886 260896 134892 260908
rect 134847 260868 134892 260896
rect 134886 260856 134892 260868
rect 134944 260856 134950 260908
rect 66530 260828 66536 260840
rect 66491 260800 66536 260828
rect 66530 260788 66536 260800
rect 66588 260788 66594 260840
rect 72234 260828 72240 260840
rect 72195 260800 72240 260828
rect 72234 260788 72240 260800
rect 72292 260788 72298 260840
rect 74994 260828 75000 260840
rect 74955 260800 75000 260828
rect 74994 260788 75000 260800
rect 75052 260788 75058 260840
rect 77570 260828 77576 260840
rect 77531 260800 77576 260828
rect 77570 260788 77576 260800
rect 77628 260788 77634 260840
rect 80330 260788 80336 260840
rect 80388 260828 80394 260840
rect 80422 260828 80428 260840
rect 80388 260800 80428 260828
rect 80388 260788 80394 260800
rect 80422 260788 80428 260800
rect 80480 260788 80486 260840
rect 95602 260828 95608 260840
rect 95563 260800 95608 260828
rect 95602 260788 95608 260800
rect 95660 260788 95666 260840
rect 124306 259468 124312 259480
rect 124267 259440 124312 259468
rect 124306 259428 124312 259440
rect 124364 259428 124370 259480
rect 124306 253920 124312 253972
rect 124364 253920 124370 253972
rect 124324 253824 124352 253920
rect 124398 253824 124404 253836
rect 124324 253796 124404 253824
rect 124398 253784 124404 253796
rect 124456 253784 124462 253836
rect 66533 251243 66591 251249
rect 66533 251209 66545 251243
rect 66579 251240 66591 251243
rect 66622 251240 66628 251252
rect 66579 251212 66628 251240
rect 66579 251209 66591 251212
rect 66533 251203 66591 251209
rect 66622 251200 66628 251212
rect 66680 251200 66686 251252
rect 72234 251240 72240 251252
rect 72195 251212 72240 251240
rect 72234 251200 72240 251212
rect 72292 251200 72298 251252
rect 74994 251240 75000 251252
rect 74955 251212 75000 251240
rect 74994 251200 75000 251212
rect 75052 251200 75058 251252
rect 77570 251240 77576 251252
rect 77531 251212 77576 251240
rect 77570 251200 77576 251212
rect 77628 251200 77634 251252
rect 81802 251200 81808 251252
rect 81860 251240 81866 251252
rect 81894 251240 81900 251252
rect 81860 251212 81900 251240
rect 81860 251200 81866 251212
rect 81894 251200 81900 251212
rect 81952 251200 81958 251252
rect 95605 251243 95663 251249
rect 95605 251209 95617 251243
rect 95651 251240 95663 251243
rect 95694 251240 95700 251252
rect 95651 251212 95700 251240
rect 95651 251209 95663 251212
rect 95605 251203 95663 251209
rect 95694 251200 95700 251212
rect 95752 251200 95758 251252
rect 85942 251132 85948 251184
rect 86000 251172 86006 251184
rect 86126 251172 86132 251184
rect 86000 251144 86132 251172
rect 86000 251132 86006 251144
rect 86126 251132 86132 251144
rect 86184 251132 86190 251184
rect 134889 251175 134947 251181
rect 134889 251141 134901 251175
rect 134935 251172 134947 251175
rect 134978 251172 134984 251184
rect 134935 251144 134984 251172
rect 134935 251141 134947 251144
rect 134889 251135 134947 251141
rect 134978 251132 134984 251144
rect 135036 251132 135042 251184
rect 74258 249772 74264 249824
rect 74316 249812 74322 249824
rect 74442 249812 74448 249824
rect 74316 249784 74448 249812
rect 74316 249772 74322 249784
rect 74442 249772 74448 249784
rect 74500 249772 74506 249824
rect 124398 244372 124404 244384
rect 124324 244344 124404 244372
rect 124324 244248 124352 244344
rect 124398 244332 124404 244344
rect 124456 244332 124462 244384
rect 140774 244264 140780 244316
rect 140832 244304 140838 244316
rect 140958 244304 140964 244316
rect 140832 244276 140964 244304
rect 140832 244264 140838 244276
rect 140958 244264 140964 244276
rect 141016 244264 141022 244316
rect 150158 244264 150164 244316
rect 150216 244304 150222 244316
rect 150342 244304 150348 244316
rect 150216 244276 150348 244304
rect 150216 244264 150222 244276
rect 150342 244264 150348 244276
rect 150400 244264 150406 244316
rect 124306 244196 124312 244248
rect 124364 244196 124370 244248
rect 134886 241516 134892 241528
rect 134847 241488 134892 241516
rect 134886 241476 134892 241488
rect 134944 241476 134950 241528
rect 77662 234648 77668 234660
rect 77588 234620 77668 234648
rect 77588 234592 77616 234620
rect 77662 234608 77668 234620
rect 77720 234608 77726 234660
rect 85942 234648 85948 234660
rect 85868 234620 85948 234648
rect 85868 234592 85896 234620
rect 85942 234608 85948 234620
rect 86000 234608 86006 234660
rect 124306 234608 124312 234660
rect 124364 234608 124370 234660
rect 134886 234608 134892 234660
rect 134944 234608 134950 234660
rect 77570 234540 77576 234592
rect 77628 234540 77634 234592
rect 85850 234540 85856 234592
rect 85908 234540 85914 234592
rect 124324 234512 124352 234608
rect 124398 234512 124404 234524
rect 124324 234484 124404 234512
rect 124398 234472 124404 234484
rect 124456 234472 124462 234524
rect 134904 234512 134932 234608
rect 134978 234512 134984 234524
rect 134904 234484 134984 234512
rect 134978 234472 134984 234484
rect 135036 234472 135042 234524
rect 66346 231820 66352 231872
rect 66404 231860 66410 231872
rect 66622 231860 66628 231872
rect 66404 231832 66628 231860
rect 66404 231820 66410 231832
rect 66622 231820 66628 231832
rect 66680 231820 66686 231872
rect 72050 231820 72056 231872
rect 72108 231860 72114 231872
rect 72234 231860 72240 231872
rect 72108 231832 72240 231860
rect 72108 231820 72114 231832
rect 72234 231820 72240 231832
rect 72292 231820 72298 231872
rect 74810 231820 74816 231872
rect 74868 231860 74874 231872
rect 74994 231860 75000 231872
rect 74868 231832 75000 231860
rect 74868 231820 74874 231832
rect 74994 231820 75000 231832
rect 75052 231820 75058 231872
rect 80330 231820 80336 231872
rect 80388 231860 80394 231872
rect 80422 231860 80428 231872
rect 80388 231832 80428 231860
rect 80388 231820 80394 231832
rect 80422 231820 80428 231832
rect 80480 231820 80486 231872
rect 81802 231820 81808 231872
rect 81860 231860 81866 231872
rect 81894 231860 81900 231872
rect 81860 231832 81900 231860
rect 81860 231820 81866 231832
rect 81894 231820 81900 231832
rect 81952 231820 81958 231872
rect 95418 231820 95424 231872
rect 95476 231860 95482 231872
rect 95694 231860 95700 231872
rect 95476 231832 95700 231860
rect 95476 231820 95482 231832
rect 95694 231820 95700 231832
rect 95752 231820 95758 231872
rect 74258 230460 74264 230512
rect 74316 230500 74322 230512
rect 74442 230500 74448 230512
rect 74316 230472 74448 230500
rect 74316 230460 74322 230472
rect 74442 230460 74448 230472
rect 74500 230460 74506 230512
rect 124306 224992 124312 225004
rect 124267 224964 124312 224992
rect 124306 224952 124312 224964
rect 124364 224952 124370 225004
rect 134886 224992 134892 225004
rect 134847 224964 134892 224992
rect 134886 224952 134892 224964
rect 134944 224952 134950 225004
rect 140774 224952 140780 225004
rect 140832 224992 140838 225004
rect 140958 224992 140964 225004
rect 140832 224964 140964 224992
rect 140832 224952 140838 224964
rect 140958 224952 140964 224964
rect 141016 224952 141022 225004
rect 150158 224952 150164 225004
rect 150216 224992 150222 225004
rect 150342 224992 150348 225004
rect 150216 224964 150348 224992
rect 150216 224952 150222 224964
rect 150342 224952 150348 224964
rect 150400 224952 150406 225004
rect 124306 222204 124312 222216
rect 124267 222176 124312 222204
rect 124306 222164 124312 222176
rect 124364 222164 124370 222216
rect 134886 222204 134892 222216
rect 134847 222176 134892 222204
rect 134886 222164 134892 222176
rect 134944 222164 134950 222216
rect 124306 215296 124312 215348
rect 124364 215296 124370 215348
rect 134886 215296 134892 215348
rect 134944 215296 134950 215348
rect 124324 215200 124352 215296
rect 124398 215200 124404 215212
rect 124324 215172 124404 215200
rect 124398 215160 124404 215172
rect 124456 215160 124462 215212
rect 134904 215200 134932 215296
rect 134978 215200 134984 215212
rect 134904 215172 134984 215200
rect 134978 215160 134984 215172
rect 135036 215160 135042 215212
rect 66346 212508 66352 212560
rect 66404 212548 66410 212560
rect 66622 212548 66628 212560
rect 66404 212520 66628 212548
rect 66404 212508 66410 212520
rect 66622 212508 66628 212520
rect 66680 212508 66686 212560
rect 72050 212508 72056 212560
rect 72108 212548 72114 212560
rect 72234 212548 72240 212560
rect 72108 212520 72240 212548
rect 72108 212508 72114 212520
rect 72234 212508 72240 212520
rect 72292 212508 72298 212560
rect 74810 212508 74816 212560
rect 74868 212548 74874 212560
rect 74994 212548 75000 212560
rect 74868 212520 75000 212548
rect 74868 212508 74874 212520
rect 74994 212508 75000 212520
rect 75052 212508 75058 212560
rect 77570 212508 77576 212560
rect 77628 212548 77634 212560
rect 77754 212548 77760 212560
rect 77628 212520 77760 212548
rect 77628 212508 77634 212520
rect 77754 212508 77760 212520
rect 77812 212508 77818 212560
rect 80330 212508 80336 212560
rect 80388 212548 80394 212560
rect 80422 212548 80428 212560
rect 80388 212520 80428 212548
rect 80388 212508 80394 212520
rect 80422 212508 80428 212520
rect 80480 212508 80486 212560
rect 81802 212508 81808 212560
rect 81860 212548 81866 212560
rect 81894 212548 81900 212560
rect 81860 212520 81900 212548
rect 81860 212508 81866 212520
rect 81894 212508 81900 212520
rect 81952 212508 81958 212560
rect 95418 212508 95424 212560
rect 95476 212548 95482 212560
rect 95694 212548 95700 212560
rect 95476 212520 95700 212548
rect 95476 212508 95482 212520
rect 95694 212508 95700 212520
rect 95752 212508 95758 212560
rect 124306 205680 124312 205692
rect 124267 205652 124312 205680
rect 124306 205640 124312 205652
rect 124364 205640 124370 205692
rect 134886 205680 134892 205692
rect 134847 205652 134892 205680
rect 134886 205640 134892 205652
rect 134944 205640 134950 205692
rect 140774 205640 140780 205692
rect 140832 205680 140838 205692
rect 140958 205680 140964 205692
rect 140832 205652 140964 205680
rect 140832 205640 140838 205652
rect 140958 205640 140964 205652
rect 141016 205640 141022 205692
rect 150158 205640 150164 205692
rect 150216 205680 150222 205692
rect 150342 205680 150348 205692
rect 150216 205652 150348 205680
rect 150216 205640 150222 205652
rect 150342 205640 150348 205652
rect 150400 205640 150406 205692
rect 85942 202852 85948 202904
rect 86000 202892 86006 202904
rect 86126 202892 86132 202904
rect 86000 202864 86132 202892
rect 86000 202852 86006 202864
rect 86126 202852 86132 202864
rect 86184 202852 86190 202904
rect 124306 202892 124312 202904
rect 124267 202864 124312 202892
rect 124306 202852 124312 202864
rect 124364 202852 124370 202904
rect 134886 202892 134892 202904
rect 134847 202864 134892 202892
rect 134886 202852 134892 202864
rect 134944 202852 134950 202904
rect 80330 202784 80336 202836
rect 80388 202824 80394 202836
rect 80422 202824 80428 202836
rect 80388 202796 80428 202824
rect 80388 202784 80394 202796
rect 80422 202784 80428 202796
rect 80480 202784 80486 202836
rect 74258 201424 74264 201476
rect 74316 201464 74322 201476
rect 74442 201464 74448 201476
rect 74316 201436 74448 201464
rect 74316 201424 74322 201436
rect 74442 201424 74448 201436
rect 74500 201424 74506 201476
rect 77662 196024 77668 196036
rect 77588 195996 77668 196024
rect 77588 195968 77616 195996
rect 77662 195984 77668 195996
rect 77720 195984 77726 196036
rect 85942 196024 85948 196036
rect 85868 195996 85948 196024
rect 85868 195968 85896 195996
rect 85942 195984 85948 195996
rect 86000 195984 86006 196036
rect 124306 195984 124312 196036
rect 124364 195984 124370 196036
rect 134886 195984 134892 196036
rect 134944 195984 134950 196036
rect 77570 195916 77576 195968
rect 77628 195916 77634 195968
rect 85850 195916 85856 195968
rect 85908 195916 85914 195968
rect 124324 195888 124352 195984
rect 124398 195888 124404 195900
rect 124324 195860 124404 195888
rect 124398 195848 124404 195860
rect 124456 195848 124462 195900
rect 134904 195888 134932 195984
rect 134978 195888 134984 195900
rect 134904 195860 134984 195888
rect 134978 195848 134984 195860
rect 135036 195848 135042 195900
rect 66346 193196 66352 193248
rect 66404 193236 66410 193248
rect 66622 193236 66628 193248
rect 66404 193208 66628 193236
rect 66404 193196 66410 193208
rect 66622 193196 66628 193208
rect 66680 193196 66686 193248
rect 72050 193196 72056 193248
rect 72108 193236 72114 193248
rect 72234 193236 72240 193248
rect 72108 193208 72240 193236
rect 72108 193196 72114 193208
rect 72234 193196 72240 193208
rect 72292 193196 72298 193248
rect 74810 193196 74816 193248
rect 74868 193236 74874 193248
rect 74994 193236 75000 193248
rect 74868 193208 75000 193236
rect 74868 193196 74874 193208
rect 74994 193196 75000 193208
rect 75052 193196 75058 193248
rect 81802 193196 81808 193248
rect 81860 193236 81866 193248
rect 81894 193236 81900 193248
rect 81860 193208 81900 193236
rect 81860 193196 81866 193208
rect 81894 193196 81900 193208
rect 81952 193196 81958 193248
rect 95418 193196 95424 193248
rect 95476 193236 95482 193248
rect 95694 193236 95700 193248
rect 95476 193208 95700 193236
rect 95476 193196 95482 193208
rect 95694 193196 95700 193208
rect 95752 193196 95758 193248
rect 160554 193196 160560 193248
rect 160612 193236 160618 193248
rect 160738 193236 160744 193248
rect 160612 193208 160744 193236
rect 160612 193196 160618 193208
rect 160738 193196 160744 193208
rect 160796 193196 160802 193248
rect 124306 186368 124312 186380
rect 124267 186340 124312 186368
rect 124306 186328 124312 186340
rect 124364 186328 124370 186380
rect 140774 186328 140780 186380
rect 140832 186368 140838 186380
rect 140958 186368 140964 186380
rect 140832 186340 140964 186368
rect 140832 186328 140838 186340
rect 140958 186328 140964 186340
rect 141016 186328 141022 186380
rect 150158 186328 150164 186380
rect 150216 186368 150222 186380
rect 150342 186368 150348 186380
rect 150216 186340 150348 186368
rect 150216 186328 150222 186340
rect 150342 186328 150348 186340
rect 150400 186328 150406 186380
rect 85942 183540 85948 183592
rect 86000 183580 86006 183592
rect 86126 183580 86132 183592
rect 86000 183552 86132 183580
rect 86000 183540 86006 183552
rect 86126 183540 86132 183552
rect 86184 183540 86190 183592
rect 124306 183580 124312 183592
rect 124267 183552 124312 183580
rect 124306 183540 124312 183552
rect 124364 183540 124370 183592
rect 134794 183540 134800 183592
rect 134852 183580 134858 183592
rect 135070 183580 135076 183592
rect 134852 183552 135076 183580
rect 134852 183540 134858 183552
rect 135070 183540 135076 183552
rect 135128 183540 135134 183592
rect 80330 183472 80336 183524
rect 80388 183512 80394 183524
rect 80422 183512 80428 183524
rect 80388 183484 80428 183512
rect 80388 183472 80394 183484
rect 80422 183472 80428 183484
rect 80480 183472 80486 183524
rect 74258 182112 74264 182164
rect 74316 182152 74322 182164
rect 74442 182152 74448 182164
rect 74316 182124 74448 182152
rect 74316 182112 74322 182124
rect 74442 182112 74448 182124
rect 74500 182112 74506 182164
rect 135070 176740 135076 176792
rect 135128 176740 135134 176792
rect 77478 176672 77484 176724
rect 77536 176712 77542 176724
rect 85942 176712 85948 176724
rect 77536 176684 77616 176712
rect 77536 176672 77542 176684
rect 77588 176656 77616 176684
rect 85868 176684 85948 176712
rect 85868 176656 85896 176684
rect 85942 176672 85948 176684
rect 86000 176672 86006 176724
rect 124306 176672 124312 176724
rect 124364 176672 124370 176724
rect 77570 176604 77576 176656
rect 77628 176604 77634 176656
rect 85850 176604 85856 176656
rect 85908 176604 85914 176656
rect 124324 176576 124352 176672
rect 124398 176576 124404 176588
rect 124324 176548 124404 176576
rect 124398 176536 124404 176548
rect 124456 176536 124462 176588
rect 134978 176536 134984 176588
rect 135036 176576 135042 176588
rect 135088 176576 135116 176740
rect 135036 176548 135116 176576
rect 135036 176536 135042 176548
rect 66346 173884 66352 173936
rect 66404 173924 66410 173936
rect 66622 173924 66628 173936
rect 66404 173896 66628 173924
rect 66404 173884 66410 173896
rect 66622 173884 66628 173896
rect 66680 173884 66686 173936
rect 72050 173884 72056 173936
rect 72108 173924 72114 173936
rect 72234 173924 72240 173936
rect 72108 173896 72240 173924
rect 72108 173884 72114 173896
rect 72234 173884 72240 173896
rect 72292 173884 72298 173936
rect 74810 173884 74816 173936
rect 74868 173924 74874 173936
rect 74994 173924 75000 173936
rect 74868 173896 75000 173924
rect 74868 173884 74874 173896
rect 74994 173884 75000 173896
rect 75052 173884 75058 173936
rect 81802 173884 81808 173936
rect 81860 173924 81866 173936
rect 81894 173924 81900 173936
rect 81860 173896 81900 173924
rect 81860 173884 81866 173896
rect 81894 173884 81900 173896
rect 81952 173884 81958 173936
rect 95418 173884 95424 173936
rect 95476 173924 95482 173936
rect 95694 173924 95700 173936
rect 95476 173896 95700 173924
rect 95476 173884 95482 173896
rect 95694 173884 95700 173896
rect 95752 173884 95758 173936
rect 140958 173884 140964 173936
rect 141016 173924 141022 173936
rect 141142 173924 141148 173936
rect 141016 173896 141148 173924
rect 141016 173884 141022 173896
rect 141142 173884 141148 173896
rect 141200 173884 141206 173936
rect 150066 173884 150072 173936
rect 150124 173924 150130 173936
rect 150342 173924 150348 173936
rect 150124 173896 150348 173924
rect 150124 173884 150130 173896
rect 150342 173884 150348 173896
rect 150400 173884 150406 173936
rect 124306 167056 124312 167068
rect 124267 167028 124312 167056
rect 124306 167016 124312 167028
rect 124364 167016 124370 167068
rect 140774 167016 140780 167068
rect 140832 167056 140838 167068
rect 140958 167056 140964 167068
rect 140832 167028 140964 167056
rect 140832 167016 140838 167028
rect 140958 167016 140964 167028
rect 141016 167016 141022 167068
rect 150158 167016 150164 167068
rect 150216 167056 150222 167068
rect 150342 167056 150348 167068
rect 150216 167028 150348 167056
rect 150216 167016 150222 167028
rect 150342 167016 150348 167028
rect 150400 167016 150406 167068
rect 78858 166948 78864 167000
rect 78916 166948 78922 167000
rect 134794 166948 134800 167000
rect 134852 166988 134858 167000
rect 134978 166988 134984 167000
rect 134852 166960 134984 166988
rect 134852 166948 134858 166960
rect 134978 166948 134984 166960
rect 135036 166948 135042 167000
rect 78876 166864 78904 166948
rect 78858 166812 78864 166864
rect 78916 166812 78922 166864
rect 124306 164268 124312 164280
rect 124267 164240 124312 164268
rect 124306 164228 124312 164240
rect 124364 164228 124370 164280
rect 66346 164160 66352 164212
rect 66404 164200 66410 164212
rect 66530 164200 66536 164212
rect 66404 164172 66536 164200
rect 66404 164160 66410 164172
rect 66530 164160 66536 164172
rect 66588 164160 66594 164212
rect 95418 164160 95424 164212
rect 95476 164200 95482 164212
rect 95602 164200 95608 164212
rect 95476 164172 95608 164200
rect 95476 164160 95482 164172
rect 95602 164160 95608 164172
rect 95660 164160 95666 164212
rect 140866 164200 140872 164212
rect 140827 164172 140872 164200
rect 140866 164160 140872 164172
rect 140924 164160 140930 164212
rect 150250 164200 150256 164212
rect 150211 164172 150256 164200
rect 150250 164160 150256 164172
rect 150308 164160 150314 164212
rect 74442 162840 74448 162852
rect 74403 162812 74448 162840
rect 74442 162800 74448 162812
rect 74500 162800 74506 162852
rect 78858 162840 78864 162852
rect 78819 162812 78864 162840
rect 78858 162800 78864 162812
rect 78916 162800 78922 162852
rect 135070 157468 135076 157480
rect 135031 157440 135076 157468
rect 135070 157428 135076 157440
rect 135128 157428 135134 157480
rect 124306 157360 124312 157412
rect 124364 157360 124370 157412
rect 80238 157292 80244 157344
rect 80296 157332 80302 157344
rect 80422 157332 80428 157344
rect 80296 157304 80428 157332
rect 80296 157292 80302 157304
rect 80422 157292 80428 157304
rect 80480 157292 80486 157344
rect 81710 157292 81716 157344
rect 81768 157332 81774 157344
rect 81894 157332 81900 157344
rect 81768 157304 81900 157332
rect 81768 157292 81774 157304
rect 81894 157292 81900 157304
rect 81952 157292 81958 157344
rect 85850 157292 85856 157344
rect 85908 157332 85914 157344
rect 86034 157332 86040 157344
rect 85908 157304 86040 157332
rect 85908 157292 85914 157304
rect 86034 157292 86040 157304
rect 86092 157292 86098 157344
rect 124324 157264 124352 157360
rect 140866 157332 140872 157344
rect 140827 157304 140872 157332
rect 140866 157292 140872 157304
rect 140924 157292 140930 157344
rect 150250 157332 150256 157344
rect 150211 157304 150256 157332
rect 150250 157292 150256 157304
rect 150308 157292 150314 157344
rect 124398 157264 124404 157276
rect 124324 157236 124404 157264
rect 124398 157224 124404 157236
rect 124456 157224 124462 157276
rect 135070 154612 135076 154624
rect 135031 154584 135076 154612
rect 135070 154572 135076 154584
rect 135128 154572 135134 154624
rect 80330 154504 80336 154556
rect 80388 154544 80394 154556
rect 80422 154544 80428 154556
rect 80388 154516 80428 154544
rect 80388 154504 80394 154516
rect 80422 154504 80428 154516
rect 80480 154504 80486 154556
rect 81802 154504 81808 154556
rect 81860 154544 81866 154556
rect 81894 154544 81900 154556
rect 81860 154516 81900 154544
rect 81860 154504 81866 154516
rect 81894 154504 81900 154516
rect 81952 154504 81958 154556
rect 124398 154504 124404 154556
rect 124456 154544 124462 154556
rect 124582 154544 124588 154556
rect 124456 154516 124588 154544
rect 124456 154504 124462 154516
rect 124582 154504 124588 154516
rect 124640 154504 124646 154556
rect 74442 153252 74448 153264
rect 74403 153224 74448 153252
rect 74442 153212 74448 153224
rect 74500 153212 74506 153264
rect 78858 153252 78864 153264
rect 78819 153224 78864 153252
rect 78858 153212 78864 153224
rect 78916 153212 78922 153264
rect 135070 147676 135076 147688
rect 135031 147648 135076 147676
rect 135070 147636 135076 147648
rect 135128 147636 135134 147688
rect 140774 147636 140780 147688
rect 140832 147676 140838 147688
rect 140958 147676 140964 147688
rect 140832 147648 140964 147676
rect 140832 147636 140838 147648
rect 140958 147636 140964 147648
rect 141016 147636 141022 147688
rect 150158 147636 150164 147688
rect 150216 147676 150222 147688
rect 150342 147676 150348 147688
rect 150216 147648 150348 147676
rect 150216 147636 150222 147648
rect 150342 147636 150348 147648
rect 150400 147636 150406 147688
rect 135070 144956 135076 144968
rect 135031 144928 135076 144956
rect 135070 144916 135076 144928
rect 135128 144916 135134 144968
rect 85850 144848 85856 144900
rect 85908 144888 85914 144900
rect 85942 144888 85948 144900
rect 85908 144860 85948 144888
rect 85908 144848 85914 144860
rect 85942 144848 85948 144860
rect 86000 144848 86006 144900
rect 140866 144888 140872 144900
rect 140827 144860 140872 144888
rect 140866 144848 140872 144860
rect 140924 144848 140930 144900
rect 150250 144888 150256 144900
rect 150211 144860 150256 144888
rect 150250 144848 150256 144860
rect 150308 144848 150314 144900
rect 74442 143528 74448 143540
rect 74403 143500 74448 143528
rect 74442 143488 74448 143500
rect 74500 143488 74506 143540
rect 74994 143528 75000 143540
rect 74955 143500 75000 143528
rect 74994 143488 75000 143500
rect 75052 143488 75058 143540
rect 78766 140020 78772 140072
rect 78824 140020 78830 140072
rect 78784 139992 78812 140020
rect 78858 139992 78864 140004
rect 78784 139964 78864 139992
rect 78858 139952 78864 139964
rect 78916 139952 78922 140004
rect 135070 138088 135076 138100
rect 134996 138060 135076 138088
rect 80330 137980 80336 138032
rect 80388 137980 80394 138032
rect 81802 137980 81808 138032
rect 81860 137980 81866 138032
rect 124306 137980 124312 138032
rect 124364 137980 124370 138032
rect 80348 137952 80376 137980
rect 80422 137952 80428 137964
rect 80348 137924 80428 137952
rect 80422 137912 80428 137924
rect 80480 137912 80486 137964
rect 81820 137952 81848 137980
rect 81894 137952 81900 137964
rect 81820 137924 81900 137952
rect 81894 137912 81900 137924
rect 81952 137912 81958 137964
rect 124324 137952 124352 137980
rect 134996 137964 135024 138060
rect 135070 138048 135076 138060
rect 135128 138048 135134 138100
rect 124398 137952 124404 137964
rect 124324 137924 124404 137952
rect 124398 137912 124404 137924
rect 124456 137912 124462 137964
rect 134978 137912 134984 137964
rect 135036 137912 135042 137964
rect 140866 137952 140872 137964
rect 140827 137924 140872 137952
rect 140866 137912 140872 137924
rect 140924 137912 140930 137964
rect 150250 137952 150256 137964
rect 150211 137924 150256 137952
rect 150250 137912 150256 137924
rect 150308 137912 150314 137964
rect 77570 135328 77576 135380
rect 77628 135328 77634 135380
rect 77588 135244 77616 135328
rect 77570 135192 77576 135244
rect 77628 135192 77634 135244
rect 124398 135192 124404 135244
rect 124456 135232 124462 135244
rect 124582 135232 124588 135244
rect 124456 135204 124588 135232
rect 124456 135192 124462 135204
rect 124582 135192 124588 135204
rect 124640 135192 124646 135244
rect 74442 133940 74448 133952
rect 74403 133912 74448 133940
rect 74442 133900 74448 133912
rect 74500 133900 74506 133952
rect 74994 133940 75000 133952
rect 74955 133912 75000 133940
rect 74994 133900 75000 133912
rect 75052 133900 75058 133952
rect 77662 133832 77668 133884
rect 77720 133872 77726 133884
rect 77846 133872 77852 133884
rect 77720 133844 77852 133872
rect 77720 133832 77726 133844
rect 77846 133832 77852 133844
rect 77904 133832 77910 133884
rect 134978 128324 134984 128376
rect 135036 128324 135042 128376
rect 140774 128324 140780 128376
rect 140832 128364 140838 128376
rect 140958 128364 140964 128376
rect 140832 128336 140964 128364
rect 140832 128324 140838 128336
rect 140958 128324 140964 128336
rect 141016 128324 141022 128376
rect 150158 128324 150164 128376
rect 150216 128364 150222 128376
rect 150342 128364 150348 128376
rect 150216 128336 150348 128364
rect 150216 128324 150222 128336
rect 150342 128324 150348 128336
rect 150400 128324 150406 128376
rect 134996 128296 135024 128324
rect 135070 128296 135076 128308
rect 134996 128268 135076 128296
rect 135070 128256 135076 128268
rect 135128 128256 135134 128308
rect 78766 125536 78772 125588
rect 78824 125536 78830 125588
rect 85850 125536 85856 125588
rect 85908 125576 85914 125588
rect 85942 125576 85948 125588
rect 85908 125548 85948 125576
rect 85908 125536 85914 125548
rect 85942 125536 85948 125548
rect 86000 125536 86006 125588
rect 140866 125576 140872 125588
rect 140827 125548 140872 125576
rect 140866 125536 140872 125548
rect 140924 125536 140930 125588
rect 150250 125576 150256 125588
rect 150211 125548 150256 125576
rect 150250 125536 150256 125548
rect 150308 125536 150314 125588
rect 78784 125440 78812 125536
rect 78858 125440 78864 125452
rect 78784 125412 78864 125440
rect 78858 125400 78864 125412
rect 78916 125400 78922 125452
rect 77478 124108 77484 124160
rect 77536 124148 77542 124160
rect 77570 124148 77576 124160
rect 77536 124120 77576 124148
rect 77536 124108 77542 124120
rect 77570 124108 77576 124120
rect 77628 124108 77634 124160
rect 134981 124151 135039 124157
rect 134981 124117 134993 124151
rect 135027 124148 135039 124151
rect 135070 124148 135076 124160
rect 135027 124120 135076 124148
rect 135027 124117 135039 124120
rect 134981 124111 135039 124117
rect 135070 124108 135076 124120
rect 135128 124108 135134 124160
rect 72234 122788 72240 122800
rect 72195 122760 72240 122788
rect 72234 122748 72240 122760
rect 72292 122748 72298 122800
rect 74994 122788 75000 122800
rect 74955 122760 75000 122788
rect 74994 122748 75000 122760
rect 75052 122748 75058 122800
rect 80330 118668 80336 118720
rect 80388 118668 80394 118720
rect 81802 118668 81808 118720
rect 81860 118668 81866 118720
rect 124306 118668 124312 118720
rect 124364 118668 124370 118720
rect 80348 118640 80376 118668
rect 80422 118640 80428 118652
rect 80348 118612 80428 118640
rect 80422 118600 80428 118612
rect 80480 118600 80486 118652
rect 81820 118640 81848 118668
rect 81894 118640 81900 118652
rect 81820 118612 81900 118640
rect 81894 118600 81900 118612
rect 81952 118600 81958 118652
rect 124324 118640 124352 118668
rect 124398 118640 124404 118652
rect 124324 118612 124404 118640
rect 124398 118600 124404 118612
rect 124456 118600 124462 118652
rect 140866 118640 140872 118652
rect 140827 118612 140872 118640
rect 140866 118600 140872 118612
rect 140924 118600 140930 118652
rect 150250 118640 150256 118652
rect 150211 118612 150256 118640
rect 150250 118600 150256 118612
rect 150308 118600 150314 118652
rect 74994 117280 75000 117292
rect 74955 117252 75000 117280
rect 74994 117240 75000 117252
rect 75052 117240 75058 117292
rect 124398 115880 124404 115932
rect 124456 115920 124462 115932
rect 124582 115920 124588 115932
rect 124456 115892 124588 115920
rect 124456 115880 124462 115892
rect 124582 115880 124588 115892
rect 124640 115880 124646 115932
rect 134978 114560 134984 114572
rect 134939 114532 134984 114560
rect 134978 114520 134984 114532
rect 135036 114520 135042 114572
rect 77570 114492 77576 114504
rect 77531 114464 77576 114492
rect 77570 114452 77576 114464
rect 77628 114452 77634 114504
rect 72234 113200 72240 113212
rect 72195 113172 72240 113200
rect 72234 113160 72240 113172
rect 72292 113160 72298 113212
rect 134978 109012 134984 109064
rect 135036 109012 135042 109064
rect 140774 109012 140780 109064
rect 140832 109052 140838 109064
rect 140958 109052 140964 109064
rect 140832 109024 140964 109052
rect 140832 109012 140838 109024
rect 140958 109012 140964 109024
rect 141016 109012 141022 109064
rect 150158 109012 150164 109064
rect 150216 109052 150222 109064
rect 150342 109052 150348 109064
rect 150216 109024 150348 109052
rect 150216 109012 150222 109024
rect 150342 109012 150348 109024
rect 150400 109012 150406 109064
rect 134996 108984 135024 109012
rect 135070 108984 135076 108996
rect 134996 108956 135076 108984
rect 135070 108944 135076 108956
rect 135128 108944 135134 108996
rect 85942 106292 85948 106344
rect 86000 106332 86006 106344
rect 86034 106332 86040 106344
rect 86000 106304 86040 106332
rect 86000 106292 86006 106304
rect 86034 106292 86040 106304
rect 86092 106292 86098 106344
rect 140866 106264 140872 106276
rect 140827 106236 140872 106264
rect 140866 106224 140872 106236
rect 140924 106224 140930 106276
rect 150250 106264 150256 106276
rect 150211 106236 150256 106264
rect 150250 106224 150256 106236
rect 150308 106224 150314 106276
rect 77570 104904 77576 104916
rect 77531 104876 77576 104904
rect 77570 104864 77576 104876
rect 77628 104864 77634 104916
rect 74442 104836 74448 104848
rect 74403 104808 74448 104836
rect 74442 104796 74448 104808
rect 74500 104796 74506 104848
rect 78766 104836 78772 104848
rect 78727 104808 78772 104836
rect 78766 104796 78772 104808
rect 78824 104796 78830 104848
rect 85942 104836 85948 104848
rect 85903 104808 85948 104836
rect 85942 104796 85948 104808
rect 86000 104796 86006 104848
rect 134981 104839 135039 104845
rect 134981 104805 134993 104839
rect 135027 104836 135039 104839
rect 135070 104836 135076 104848
rect 135027 104808 135076 104836
rect 135027 104805 135039 104808
rect 134981 104799 135039 104805
rect 135070 104796 135076 104808
rect 135128 104796 135134 104848
rect 72237 102119 72295 102125
rect 72237 102085 72249 102119
rect 72283 102116 72295 102119
rect 72326 102116 72332 102128
rect 72283 102088 72332 102116
rect 72283 102085 72295 102088
rect 72237 102079 72295 102085
rect 72326 102076 72332 102088
rect 72384 102076 72390 102128
rect 124306 99356 124312 99408
rect 124364 99356 124370 99408
rect 124324 99328 124352 99356
rect 124398 99328 124404 99340
rect 124324 99300 124404 99328
rect 124398 99288 124404 99300
rect 124456 99288 124462 99340
rect 140866 99328 140872 99340
rect 140827 99300 140872 99328
rect 140866 99288 140872 99300
rect 140924 99288 140930 99340
rect 150250 99328 150256 99340
rect 150211 99300 150256 99328
rect 150250 99288 150256 99300
rect 150308 99288 150314 99340
rect 124398 96568 124404 96620
rect 124456 96608 124462 96620
rect 124582 96608 124588 96620
rect 124456 96580 124588 96608
rect 124456 96568 124462 96580
rect 124582 96568 124588 96580
rect 124640 96568 124646 96620
rect 74442 95248 74448 95260
rect 74403 95220 74448 95248
rect 74442 95208 74448 95220
rect 74500 95208 74506 95260
rect 78769 95251 78827 95257
rect 78769 95217 78781 95251
rect 78815 95248 78827 95251
rect 78950 95248 78956 95260
rect 78815 95220 78956 95248
rect 78815 95217 78827 95220
rect 78769 95211 78827 95217
rect 78950 95208 78956 95220
rect 79008 95208 79014 95260
rect 85945 95251 86003 95257
rect 85945 95217 85957 95251
rect 85991 95248 86003 95251
rect 86034 95248 86040 95260
rect 85991 95220 86040 95248
rect 85991 95217 86003 95220
rect 85945 95211 86003 95217
rect 86034 95208 86040 95220
rect 86092 95208 86098 95260
rect 74994 93820 75000 93832
rect 74955 93792 75000 93820
rect 74994 93780 75000 93792
rect 75052 93780 75058 93832
rect 72234 92528 72240 92540
rect 72195 92500 72240 92528
rect 72234 92488 72240 92500
rect 72292 92488 72298 92540
rect 140774 89700 140780 89752
rect 140832 89740 140838 89752
rect 140958 89740 140964 89752
rect 140832 89712 140964 89740
rect 140832 89700 140838 89712
rect 140958 89700 140964 89712
rect 141016 89700 141022 89752
rect 150158 89700 150164 89752
rect 150216 89740 150222 89752
rect 150342 89740 150348 89752
rect 150216 89712 150348 89740
rect 150216 89700 150222 89712
rect 150342 89700 150348 89712
rect 150400 89700 150406 89752
rect 134978 89672 134984 89684
rect 134939 89644 134984 89672
rect 134978 89632 134984 89644
rect 135036 89632 135042 89684
rect 66349 86955 66407 86961
rect 66349 86921 66361 86955
rect 66395 86952 66407 86955
rect 66438 86952 66444 86964
rect 66395 86924 66444 86952
rect 66395 86921 66407 86924
rect 66349 86915 66407 86921
rect 66438 86912 66444 86924
rect 66496 86912 66502 86964
rect 85853 86955 85911 86961
rect 85853 86921 85865 86955
rect 85899 86952 85911 86955
rect 85942 86952 85948 86964
rect 85899 86924 85948 86952
rect 85899 86921 85911 86924
rect 85853 86915 85911 86921
rect 85942 86912 85948 86924
rect 86000 86912 86006 86964
rect 95421 86955 95479 86961
rect 95421 86921 95433 86955
rect 95467 86952 95479 86955
rect 95510 86952 95516 86964
rect 95467 86924 95516 86952
rect 95467 86921 95479 86924
rect 95421 86915 95479 86921
rect 95510 86912 95516 86924
rect 95568 86912 95574 86964
rect 140866 86952 140872 86964
rect 140827 86924 140872 86952
rect 140866 86912 140872 86924
rect 140924 86912 140930 86964
rect 150250 86952 150256 86964
rect 150211 86924 150256 86952
rect 150250 86912 150256 86924
rect 150308 86912 150314 86964
rect 160738 86884 160744 86896
rect 160699 86856 160744 86884
rect 160738 86844 160744 86856
rect 160796 86844 160802 86896
rect 78766 85552 78772 85604
rect 78824 85592 78830 85604
rect 78950 85592 78956 85604
rect 78824 85564 78956 85592
rect 78824 85552 78830 85564
rect 78950 85552 78956 85564
rect 79008 85552 79014 85604
rect 74994 84300 75000 84312
rect 74955 84272 75000 84300
rect 74994 84260 75000 84272
rect 75052 84260 75058 84312
rect 74994 84164 75000 84176
rect 74955 84136 75000 84164
rect 74994 84124 75000 84136
rect 75052 84124 75058 84176
rect 134702 82084 134708 82136
rect 134760 82124 134766 82136
rect 135070 82124 135076 82136
rect 134760 82096 135076 82124
rect 134760 82084 134766 82096
rect 135070 82084 135076 82096
rect 135128 82084 135134 82136
rect 81710 80152 81716 80164
rect 81636 80124 81716 80152
rect 81636 80028 81664 80124
rect 81710 80112 81716 80124
rect 81768 80112 81774 80164
rect 124306 80044 124312 80096
rect 124364 80044 124370 80096
rect 81618 79976 81624 80028
rect 81676 79976 81682 80028
rect 124324 79948 124352 80044
rect 124398 79948 124404 79960
rect 124324 79920 124404 79948
rect 124398 79908 124404 79920
rect 124456 79908 124462 79960
rect 66346 77296 66352 77308
rect 66307 77268 66352 77296
rect 66346 77256 66352 77268
rect 66404 77256 66410 77308
rect 85850 77296 85856 77308
rect 85811 77268 85856 77296
rect 85850 77256 85856 77268
rect 85908 77256 85914 77308
rect 95418 77296 95424 77308
rect 95379 77268 95424 77296
rect 95418 77256 95424 77268
rect 95476 77256 95482 77308
rect 140869 77299 140927 77305
rect 140869 77265 140881 77299
rect 140915 77296 140927 77299
rect 140958 77296 140964 77308
rect 140915 77268 140964 77296
rect 140915 77265 140927 77268
rect 140869 77259 140927 77265
rect 140958 77256 140964 77268
rect 141016 77256 141022 77308
rect 150253 77299 150311 77305
rect 150253 77265 150265 77299
rect 150299 77296 150311 77299
rect 150342 77296 150348 77308
rect 150299 77268 150348 77296
rect 150299 77265 150311 77268
rect 150253 77259 150311 77265
rect 150342 77256 150348 77268
rect 150400 77256 150406 77308
rect 160738 77296 160744 77308
rect 160699 77268 160744 77296
rect 160738 77256 160744 77268
rect 160796 77256 160802 77308
rect 81618 77228 81624 77240
rect 81579 77200 81624 77228
rect 81618 77188 81624 77200
rect 81676 77188 81682 77240
rect 66346 77160 66352 77172
rect 66307 77132 66352 77160
rect 66346 77120 66352 77132
rect 66404 77120 66410 77172
rect 95418 77160 95424 77172
rect 95379 77132 95424 77160
rect 95418 77120 95424 77132
rect 95476 77120 95482 77172
rect 140869 77163 140927 77169
rect 140869 77129 140881 77163
rect 140915 77160 140927 77163
rect 140958 77160 140964 77172
rect 140915 77132 140964 77160
rect 140915 77129 140927 77132
rect 140869 77123 140927 77129
rect 140958 77120 140964 77132
rect 141016 77120 141022 77172
rect 78766 75896 78772 75948
rect 78824 75936 78830 75948
rect 78858 75936 78864 75948
rect 78824 75908 78864 75936
rect 78824 75896 78830 75908
rect 78858 75896 78864 75908
rect 78916 75896 78922 75948
rect 74994 74536 75000 74588
rect 75052 74576 75058 74588
rect 75052 74548 75097 74576
rect 75052 74536 75058 74548
rect 74813 71111 74871 71117
rect 74813 71077 74825 71111
rect 74859 71108 74871 71111
rect 74994 71108 75000 71120
rect 74859 71080 75000 71108
rect 74859 71077 74871 71080
rect 74813 71071 74871 71077
rect 74994 71068 75000 71080
rect 75052 71068 75058 71120
rect 134978 70496 134984 70508
rect 134904 70468 134984 70496
rect 80330 70388 80336 70440
rect 80388 70388 80394 70440
rect 80348 70304 80376 70388
rect 134904 70372 134932 70468
rect 134978 70456 134984 70468
rect 135036 70456 135042 70508
rect 150158 70388 150164 70440
rect 150216 70428 150222 70440
rect 150216 70400 150296 70428
rect 150216 70388 150222 70400
rect 150268 70372 150296 70400
rect 134886 70320 134892 70372
rect 134944 70320 134950 70372
rect 150250 70320 150256 70372
rect 150308 70320 150314 70372
rect 66349 70295 66407 70301
rect 66349 70261 66361 70295
rect 66395 70292 66407 70295
rect 66438 70292 66444 70304
rect 66395 70264 66444 70292
rect 66395 70261 66407 70264
rect 66349 70255 66407 70261
rect 66438 70252 66444 70264
rect 66496 70252 66502 70304
rect 80330 70252 80336 70304
rect 80388 70252 80394 70304
rect 81621 70295 81679 70301
rect 81621 70261 81633 70295
rect 81667 70292 81679 70295
rect 81710 70292 81716 70304
rect 81667 70264 81716 70292
rect 81667 70261 81679 70264
rect 81621 70255 81679 70261
rect 81710 70252 81716 70264
rect 81768 70252 81774 70304
rect 95421 70295 95479 70301
rect 95421 70261 95433 70295
rect 95467 70292 95479 70295
rect 95510 70292 95516 70304
rect 95467 70264 95516 70292
rect 95467 70261 95479 70264
rect 95421 70255 95479 70261
rect 95510 70252 95516 70264
rect 95568 70252 95574 70304
rect 77570 67708 77576 67720
rect 77496 67680 77576 67708
rect 77496 67652 77524 67680
rect 77570 67668 77576 67680
rect 77628 67668 77634 67720
rect 77478 67600 77484 67652
rect 77536 67600 77542 67652
rect 140866 67640 140872 67652
rect 140827 67612 140872 67640
rect 140866 67600 140872 67612
rect 140924 67600 140930 67652
rect 74810 66280 74816 66292
rect 74771 66252 74816 66280
rect 74810 66240 74816 66252
rect 74868 66240 74874 66292
rect 124398 66240 124404 66292
rect 124456 66280 124462 66292
rect 124582 66280 124588 66292
rect 124456 66252 124588 66280
rect 124456 66240 124462 66252
rect 124582 66240 124588 66252
rect 124640 66240 124646 66292
rect 72142 66172 72148 66224
rect 72200 66212 72206 66224
rect 72418 66212 72424 66224
rect 72200 66184 72424 66212
rect 72200 66172 72206 66184
rect 72418 66172 72424 66184
rect 72476 66172 72482 66224
rect 74442 66212 74448 66224
rect 74403 66184 74448 66212
rect 74442 66172 74448 66184
rect 74500 66172 74506 66224
rect 77478 66212 77484 66224
rect 77439 66184 77484 66212
rect 77478 66172 77484 66184
rect 77536 66172 77542 66224
rect 134886 66172 134892 66224
rect 134944 66212 134950 66224
rect 135070 66212 135076 66224
rect 134944 66184 135076 66212
rect 134944 66172 134950 66184
rect 135070 66172 135076 66184
rect 135128 66172 135134 66224
rect 72418 64852 72424 64864
rect 72379 64824 72424 64852
rect 72418 64812 72424 64824
rect 72476 64812 72482 64864
rect 74810 64852 74816 64864
rect 74771 64824 74816 64852
rect 74810 64812 74816 64824
rect 74868 64812 74874 64864
rect 66438 60664 66444 60716
rect 66496 60704 66502 60716
rect 66622 60704 66628 60716
rect 66496 60676 66628 60704
rect 66496 60664 66502 60676
rect 66622 60664 66628 60676
rect 66680 60664 66686 60716
rect 80238 60664 80244 60716
rect 80296 60704 80302 60716
rect 80422 60704 80428 60716
rect 80296 60676 80428 60704
rect 80296 60664 80302 60676
rect 80422 60664 80428 60676
rect 80480 60664 80486 60716
rect 81710 60664 81716 60716
rect 81768 60704 81774 60716
rect 81894 60704 81900 60716
rect 81768 60676 81900 60704
rect 81768 60664 81774 60676
rect 81894 60664 81900 60676
rect 81952 60664 81958 60716
rect 95510 60664 95516 60716
rect 95568 60704 95574 60716
rect 95694 60704 95700 60716
rect 95568 60676 95700 60704
rect 95568 60664 95574 60676
rect 95694 60664 95700 60676
rect 95752 60664 95758 60716
rect 124398 60596 124404 60648
rect 124456 60636 124462 60648
rect 124582 60636 124588 60648
rect 124456 60608 124588 60636
rect 124456 60596 124462 60608
rect 124582 60596 124588 60608
rect 124640 60596 124646 60648
rect 66533 57919 66591 57925
rect 66533 57885 66545 57919
rect 66579 57916 66591 57919
rect 66622 57916 66628 57928
rect 66579 57888 66628 57916
rect 66579 57885 66591 57888
rect 66533 57879 66591 57885
rect 66622 57876 66628 57888
rect 66680 57876 66686 57928
rect 95605 57919 95663 57925
rect 95605 57885 95617 57919
rect 95651 57916 95663 57919
rect 95694 57916 95700 57928
rect 95651 57888 95700 57916
rect 95651 57885 95663 57888
rect 95605 57879 95663 57885
rect 95694 57876 95700 57888
rect 95752 57876 95758 57928
rect 140869 57919 140927 57925
rect 140869 57885 140881 57919
rect 140915 57916 140927 57919
rect 140958 57916 140964 57928
rect 140915 57888 140964 57916
rect 140915 57885 140927 57888
rect 140869 57879 140927 57885
rect 140958 57876 140964 57888
rect 141016 57876 141022 57928
rect 150253 57919 150311 57925
rect 150253 57885 150265 57919
rect 150299 57916 150311 57919
rect 150342 57916 150348 57928
rect 150299 57888 150348 57916
rect 150299 57885 150311 57888
rect 150253 57879 150311 57885
rect 150342 57876 150348 57888
rect 150400 57876 150406 57928
rect 74442 56624 74448 56636
rect 74403 56596 74448 56624
rect 74442 56584 74448 56596
rect 74500 56584 74506 56636
rect 72418 56556 72424 56568
rect 72379 56528 72424 56556
rect 72418 56516 72424 56528
rect 72476 56516 72482 56568
rect 124398 56556 124404 56568
rect 124359 56528 124404 56556
rect 124398 56516 124404 56528
rect 124456 56516 124462 56568
rect 74813 55267 74871 55273
rect 74813 55233 74825 55267
rect 74859 55264 74871 55267
rect 74902 55264 74908 55276
rect 74859 55236 74908 55264
rect 74859 55233 74871 55236
rect 74813 55227 74871 55233
rect 74902 55224 74908 55236
rect 74960 55224 74966 55276
rect 72329 55199 72387 55205
rect 72329 55165 72341 55199
rect 72375 55196 72387 55199
rect 72418 55196 72424 55208
rect 72375 55168 72424 55196
rect 72375 55165 72387 55168
rect 72329 55159 72387 55165
rect 72418 55156 72424 55168
rect 72476 55156 72482 55208
rect 140866 51048 140872 51060
rect 140827 51020 140872 51048
rect 140866 51008 140872 51020
rect 140924 51008 140930 51060
rect 77478 48396 77484 48408
rect 77439 48368 77484 48396
rect 77478 48356 77484 48368
rect 77536 48356 77542 48408
rect 66530 48328 66536 48340
rect 66491 48300 66536 48328
rect 66530 48288 66536 48300
rect 66588 48288 66594 48340
rect 95602 48328 95608 48340
rect 95563 48300 95608 48328
rect 95602 48288 95608 48300
rect 95660 48288 95666 48340
rect 150250 48328 150256 48340
rect 150211 48300 150256 48328
rect 150250 48288 150256 48300
rect 150308 48288 150314 48340
rect 124401 46971 124459 46977
rect 124401 46937 124413 46971
rect 124447 46968 124459 46971
rect 124490 46968 124496 46980
rect 124447 46940 124496 46968
rect 124447 46937 124459 46940
rect 124401 46931 124459 46937
rect 124490 46928 124496 46940
rect 124548 46928 124554 46980
rect 74442 46900 74448 46912
rect 74403 46872 74448 46900
rect 74442 46860 74448 46872
rect 74500 46860 74506 46912
rect 74902 46860 74908 46912
rect 74960 46900 74966 46912
rect 75086 46900 75092 46912
rect 74960 46872 75092 46900
rect 74960 46860 74966 46872
rect 75086 46860 75092 46872
rect 75144 46860 75150 46912
rect 77478 46860 77484 46912
rect 77536 46900 77542 46912
rect 77754 46900 77760 46912
rect 77536 46872 77760 46900
rect 77536 46860 77542 46872
rect 77754 46860 77760 46872
rect 77812 46860 77818 46912
rect 134886 46860 134892 46912
rect 134944 46900 134950 46912
rect 135070 46900 135076 46912
rect 134944 46872 135076 46900
rect 134944 46860 134950 46872
rect 135070 46860 135076 46872
rect 135128 46860 135134 46912
rect 72326 45676 72332 45688
rect 72287 45648 72332 45676
rect 72326 45636 72332 45648
rect 72384 45636 72390 45688
rect 72326 45540 72332 45552
rect 72287 45512 72332 45540
rect 72326 45500 72332 45512
rect 72384 45500 72390 45552
rect 74997 45543 75055 45549
rect 74997 45509 75009 45543
rect 75043 45540 75055 45543
rect 75086 45540 75092 45552
rect 75043 45512 75092 45540
rect 75043 45509 75055 45512
rect 74997 45503 75055 45509
rect 75086 45500 75092 45512
rect 75144 45500 75150 45552
rect 66438 41352 66444 41404
rect 66496 41392 66502 41404
rect 66622 41392 66628 41404
rect 66496 41364 66628 41392
rect 66496 41352 66502 41364
rect 66622 41352 66628 41364
rect 66680 41352 66686 41404
rect 80238 41352 80244 41404
rect 80296 41392 80302 41404
rect 80422 41392 80428 41404
rect 80296 41364 80428 41392
rect 80296 41352 80302 41364
rect 80422 41352 80428 41364
rect 80480 41352 80486 41404
rect 81710 41352 81716 41404
rect 81768 41392 81774 41404
rect 81894 41392 81900 41404
rect 81768 41364 81900 41392
rect 81768 41352 81774 41364
rect 81894 41352 81900 41364
rect 81952 41352 81958 41404
rect 95510 41352 95516 41404
rect 95568 41392 95574 41404
rect 95694 41392 95700 41404
rect 95568 41364 95700 41392
rect 95568 41352 95574 41364
rect 95694 41352 95700 41364
rect 95752 41352 95758 41404
rect 66533 38607 66591 38613
rect 66533 38573 66545 38607
rect 66579 38604 66591 38607
rect 66622 38604 66628 38616
rect 66579 38576 66628 38604
rect 66579 38573 66591 38576
rect 66533 38567 66591 38573
rect 66622 38564 66628 38576
rect 66680 38564 66686 38616
rect 78858 38604 78864 38616
rect 78819 38576 78864 38604
rect 78858 38564 78864 38576
rect 78916 38564 78922 38616
rect 95605 38607 95663 38613
rect 95605 38573 95617 38607
rect 95651 38604 95663 38607
rect 95694 38604 95700 38616
rect 95651 38576 95700 38604
rect 95651 38573 95663 38576
rect 95605 38567 95663 38573
rect 95694 38564 95700 38576
rect 95752 38564 95758 38616
rect 140869 38607 140927 38613
rect 140869 38573 140881 38607
rect 140915 38604 140927 38607
rect 140958 38604 140964 38616
rect 140915 38576 140964 38604
rect 140915 38573 140927 38576
rect 140869 38567 140927 38573
rect 140958 38564 140964 38576
rect 141016 38564 141022 38616
rect 150253 38607 150311 38613
rect 150253 38573 150265 38607
rect 150299 38604 150311 38607
rect 150342 38604 150348 38616
rect 150299 38576 150348 38604
rect 150299 38573 150311 38576
rect 150253 38567 150311 38573
rect 150342 38564 150348 38576
rect 150400 38564 150406 38616
rect 74442 37312 74448 37324
rect 74403 37284 74448 37312
rect 74442 37272 74448 37284
rect 74500 37272 74506 37324
rect 74997 37247 75055 37253
rect 74997 37213 75009 37247
rect 75043 37244 75055 37247
rect 75086 37244 75092 37256
rect 75043 37216 75092 37244
rect 75043 37213 75055 37216
rect 74997 37207 75055 37213
rect 75086 37204 75092 37216
rect 75144 37204 75150 37256
rect 72142 31696 72148 31748
rect 72200 31736 72206 31748
rect 72329 31739 72387 31745
rect 72329 31736 72341 31739
rect 72200 31708 72341 31736
rect 72200 31696 72206 31708
rect 72329 31705 72341 31708
rect 72375 31705 72387 31739
rect 140866 31736 140872 31748
rect 140827 31708 140872 31736
rect 72329 31699 72387 31705
rect 140866 31696 140872 31708
rect 140924 31696 140930 31748
rect 74810 29724 74816 29776
rect 74868 29764 74874 29776
rect 75086 29764 75092 29776
rect 74868 29736 75092 29764
rect 74868 29724 74874 29736
rect 75086 29724 75092 29736
rect 75144 29724 75150 29776
rect 66530 29016 66536 29028
rect 66491 28988 66536 29016
rect 66530 28976 66536 28988
rect 66588 28976 66594 29028
rect 78858 29016 78864 29028
rect 78819 28988 78864 29016
rect 78858 28976 78864 28988
rect 78916 28976 78922 29028
rect 81802 28976 81808 29028
rect 81860 29016 81866 29028
rect 81894 29016 81900 29028
rect 81860 28988 81900 29016
rect 81860 28976 81866 28988
rect 81894 28976 81900 28988
rect 81952 28976 81958 29028
rect 85850 28976 85856 29028
rect 85908 28976 85914 29028
rect 95602 29016 95608 29028
rect 95563 28988 95608 29016
rect 95602 28976 95608 28988
rect 95660 28976 95666 29028
rect 150250 29016 150256 29028
rect 150211 28988 150256 29016
rect 150250 28976 150256 28988
rect 150308 28976 150314 29028
rect 77202 28840 77208 28892
rect 77260 28880 77266 28892
rect 77754 28880 77760 28892
rect 77260 28852 77760 28880
rect 77260 28840 77266 28852
rect 77754 28840 77760 28852
rect 77812 28840 77818 28892
rect 85868 28880 85896 28976
rect 85942 28880 85948 28892
rect 85868 28852 85948 28880
rect 85942 28840 85948 28852
rect 86000 28840 86006 28892
rect 124398 27616 124404 27668
rect 124456 27656 124462 27668
rect 124582 27656 124588 27668
rect 124456 27628 124588 27656
rect 124456 27616 124462 27628
rect 124582 27616 124588 27628
rect 124640 27616 124646 27668
rect 72142 27548 72148 27600
rect 72200 27548 72206 27600
rect 74261 27591 74319 27597
rect 74261 27557 74273 27591
rect 74307 27588 74319 27591
rect 74442 27588 74448 27600
rect 74307 27560 74448 27588
rect 74307 27557 74319 27560
rect 74261 27551 74319 27557
rect 74442 27548 74448 27560
rect 74500 27548 74506 27600
rect 74810 27548 74816 27600
rect 74868 27588 74874 27600
rect 74905 27591 74963 27597
rect 74905 27588 74917 27591
rect 74868 27560 74917 27588
rect 74868 27548 74874 27560
rect 74905 27557 74917 27560
rect 74951 27557 74963 27591
rect 134886 27588 134892 27600
rect 134847 27560 134892 27588
rect 74905 27551 74963 27557
rect 134886 27548 134892 27560
rect 134944 27548 134950 27600
rect 72160 27520 72188 27548
rect 72326 27520 72332 27532
rect 72160 27492 72332 27520
rect 72326 27480 72332 27492
rect 72384 27480 72390 27532
rect 85942 26188 85948 26240
rect 86000 26228 86006 26240
rect 86034 26228 86040 26240
rect 86000 26200 86040 26228
rect 86000 26188 86006 26200
rect 86034 26188 86040 26200
rect 86092 26188 86098 26240
rect 66438 22040 66444 22092
rect 66496 22080 66502 22092
rect 66622 22080 66628 22092
rect 66496 22052 66628 22080
rect 66496 22040 66502 22052
rect 66622 22040 66628 22052
rect 66680 22040 66686 22092
rect 80238 22040 80244 22092
rect 80296 22080 80302 22092
rect 80422 22080 80428 22092
rect 80296 22052 80428 22080
rect 80296 22040 80302 22052
rect 80422 22040 80428 22052
rect 80480 22040 80486 22092
rect 81710 22040 81716 22092
rect 81768 22080 81774 22092
rect 81894 22080 81900 22092
rect 81768 22052 81900 22080
rect 81768 22040 81774 22052
rect 81894 22040 81900 22052
rect 81952 22040 81958 22092
rect 95510 22040 95516 22092
rect 95568 22080 95574 22092
rect 95694 22080 95700 22092
rect 95568 22052 95700 22080
rect 95568 22040 95574 22052
rect 95694 22040 95700 22052
rect 95752 22040 95758 22092
rect 160646 19320 160652 19372
rect 160704 19360 160710 19372
rect 160738 19360 160744 19372
rect 160704 19332 160744 19360
rect 160704 19320 160710 19332
rect 160738 19320 160744 19332
rect 160796 19320 160802 19372
rect 66622 19292 66628 19304
rect 66583 19264 66628 19292
rect 66622 19252 66628 19264
rect 66680 19252 66686 19304
rect 95694 19292 95700 19304
rect 95655 19264 95700 19292
rect 95694 19252 95700 19264
rect 95752 19252 95758 19304
rect 77202 19184 77208 19236
rect 77260 19224 77266 19236
rect 77754 19224 77760 19236
rect 77260 19196 77760 19224
rect 77260 19184 77266 19196
rect 77754 19184 77760 19196
rect 77812 19184 77818 19236
rect 124398 17960 124404 18012
rect 124456 18000 124462 18012
rect 124582 18000 124588 18012
rect 124456 17972 124588 18000
rect 124456 17960 124462 17972
rect 124582 17960 124588 17972
rect 124640 17960 124646 18012
rect 134889 18003 134947 18009
rect 134889 17969 134901 18003
rect 134935 18000 134947 18003
rect 134978 18000 134984 18012
rect 134935 17972 134984 18000
rect 134935 17969 134947 17972
rect 134889 17963 134947 17969
rect 134978 17960 134984 17972
rect 135036 17960 135042 18012
rect 243998 16532 244004 16584
rect 244056 16572 244062 16584
rect 485774 16572 485780 16584
rect 244056 16544 485780 16572
rect 244056 16532 244062 16544
rect 485774 16532 485780 16544
rect 485832 16532 485838 16584
rect 245378 16464 245384 16516
rect 245436 16504 245442 16516
rect 489914 16504 489920 16516
rect 245436 16476 489920 16504
rect 245436 16464 245442 16476
rect 489914 16464 489920 16476
rect 489972 16464 489978 16516
rect 246850 16396 246856 16448
rect 246908 16436 246914 16448
rect 494054 16436 494060 16448
rect 246908 16408 494060 16436
rect 246908 16396 246914 16408
rect 494054 16396 494060 16408
rect 494112 16396 494118 16448
rect 246758 16328 246764 16380
rect 246816 16368 246822 16380
rect 494146 16368 494152 16380
rect 246816 16340 494152 16368
rect 246816 16328 246822 16340
rect 494146 16328 494152 16340
rect 494204 16328 494210 16380
rect 248138 16260 248144 16312
rect 248196 16300 248202 16312
rect 496814 16300 496820 16312
rect 248196 16272 496820 16300
rect 248196 16260 248202 16272
rect 496814 16260 496820 16272
rect 496872 16260 496878 16312
rect 249518 16192 249524 16244
rect 249576 16232 249582 16244
rect 500954 16232 500960 16244
rect 249576 16204 500960 16232
rect 249576 16192 249582 16204
rect 500954 16192 500960 16204
rect 501012 16192 501018 16244
rect 250898 16124 250904 16176
rect 250956 16164 250962 16176
rect 503714 16164 503720 16176
rect 250956 16136 503720 16164
rect 250956 16124 250962 16136
rect 503714 16124 503720 16136
rect 503772 16124 503778 16176
rect 252278 16056 252284 16108
rect 252336 16096 252342 16108
rect 507854 16096 507860 16108
rect 252336 16068 507860 16096
rect 252336 16056 252342 16068
rect 507854 16056 507860 16068
rect 507912 16056 507918 16108
rect 274358 15988 274364 16040
rect 274416 16028 274422 16040
rect 567194 16028 567200 16040
rect 274416 16000 567200 16028
rect 274416 15988 274422 16000
rect 567194 15988 567200 16000
rect 567252 15988 567258 16040
rect 277118 15920 277124 15972
rect 277176 15960 277182 15972
rect 574094 15960 574100 15972
rect 277176 15932 574100 15960
rect 277176 15920 277182 15932
rect 574094 15920 574100 15932
rect 574152 15920 574158 15972
rect 278498 15852 278504 15904
rect 278556 15892 278562 15904
rect 578234 15892 578240 15904
rect 278556 15864 578240 15892
rect 278556 15852 278562 15864
rect 578234 15852 578240 15864
rect 578292 15852 578298 15904
rect 242526 15784 242532 15836
rect 242584 15824 242590 15836
rect 483014 15824 483020 15836
rect 242584 15796 483020 15824
rect 242584 15784 242590 15796
rect 483014 15784 483020 15796
rect 483072 15784 483078 15836
rect 227438 15716 227444 15768
rect 227496 15756 227502 15768
rect 442994 15756 443000 15768
rect 227496 15728 443000 15756
rect 227496 15716 227502 15728
rect 442994 15716 443000 15728
rect 443052 15716 443058 15768
rect 219158 15648 219164 15700
rect 219216 15688 219222 15700
rect 420914 15688 420920 15700
rect 219216 15660 420920 15688
rect 219216 15648 219222 15660
rect 420914 15648 420920 15660
rect 420972 15648 420978 15700
rect 213638 15580 213644 15632
rect 213696 15620 213702 15632
rect 407114 15620 407120 15632
rect 213696 15592 407120 15620
rect 213696 15580 213702 15592
rect 407114 15580 407120 15592
rect 407172 15580 407178 15632
rect 180518 15512 180524 15564
rect 180576 15552 180582 15564
rect 317414 15552 317420 15564
rect 180576 15524 317420 15552
rect 180576 15512 180582 15524
rect 317414 15512 317420 15524
rect 317472 15512 317478 15564
rect 215018 15104 215024 15156
rect 215076 15144 215082 15156
rect 408494 15144 408500 15156
rect 215076 15116 408500 15144
rect 215076 15104 215082 15116
rect 408494 15104 408500 15116
rect 408552 15104 408558 15156
rect 223298 15036 223304 15088
rect 223356 15076 223362 15088
rect 431954 15076 431960 15088
rect 223356 15048 431960 15076
rect 223356 15036 223362 15048
rect 431954 15036 431960 15048
rect 432012 15036 432018 15088
rect 226058 14968 226064 15020
rect 226116 15008 226122 15020
rect 438854 15008 438860 15020
rect 226116 14980 438860 15008
rect 226116 14968 226122 14980
rect 438854 14968 438860 14980
rect 438912 14968 438918 15020
rect 228818 14900 228824 14952
rect 228876 14940 228882 14952
rect 445754 14940 445760 14952
rect 228876 14912 445760 14940
rect 228876 14900 228882 14912
rect 445754 14900 445760 14912
rect 445812 14900 445818 14952
rect 231578 14832 231584 14884
rect 231636 14872 231642 14884
rect 452654 14872 452660 14884
rect 231636 14844 452660 14872
rect 231636 14832 231642 14844
rect 452654 14832 452660 14844
rect 452712 14832 452718 14884
rect 234338 14764 234344 14816
rect 234396 14804 234402 14816
rect 459554 14804 459560 14816
rect 234396 14776 459560 14804
rect 234396 14764 234402 14776
rect 459554 14764 459560 14776
rect 459612 14764 459618 14816
rect 237098 14696 237104 14748
rect 237156 14736 237162 14748
rect 467834 14736 467840 14748
rect 237156 14708 467840 14736
rect 237156 14696 237162 14708
rect 467834 14696 467840 14708
rect 467892 14696 467898 14748
rect 239858 14628 239864 14680
rect 239916 14668 239922 14680
rect 474734 14668 474740 14680
rect 239916 14640 474740 14668
rect 239916 14628 239922 14640
rect 474734 14628 474740 14640
rect 474792 14628 474798 14680
rect 242618 14560 242624 14612
rect 242676 14600 242682 14612
rect 481634 14600 481640 14612
rect 242676 14572 481640 14600
rect 242676 14560 242682 14572
rect 481634 14560 481640 14572
rect 481692 14560 481698 14612
rect 244090 14492 244096 14544
rect 244148 14532 244154 14544
rect 487154 14532 487160 14544
rect 244148 14504 487160 14532
rect 244148 14492 244154 14504
rect 487154 14492 487160 14504
rect 487212 14492 487218 14544
rect 245470 14424 245476 14476
rect 245528 14464 245534 14476
rect 491294 14464 491300 14476
rect 245528 14436 491300 14464
rect 245528 14424 245534 14436
rect 491294 14424 491300 14436
rect 491352 14424 491358 14476
rect 213730 14356 213736 14408
rect 213788 14396 213794 14408
rect 405734 14396 405740 14408
rect 213788 14368 405740 14396
rect 213788 14356 213794 14368
rect 405734 14356 405740 14368
rect 405792 14356 405798 14408
rect 212258 14288 212264 14340
rect 212316 14328 212322 14340
rect 401594 14328 401600 14340
rect 212316 14300 401600 14328
rect 212316 14288 212322 14300
rect 401594 14288 401600 14300
rect 401652 14288 401658 14340
rect 208118 14220 208124 14272
rect 208176 14260 208182 14272
rect 390554 14260 390560 14272
rect 208176 14232 390560 14260
rect 208176 14220 208182 14232
rect 390554 14220 390560 14232
rect 390612 14220 390618 14272
rect 176470 14152 176476 14204
rect 176528 14192 176534 14204
rect 304994 14192 305000 14204
rect 176528 14164 305000 14192
rect 176528 14152 176534 14164
rect 304994 14152 305000 14164
rect 305052 14152 305058 14204
rect 175090 14084 175096 14136
rect 175148 14124 175154 14136
rect 302234 14124 302240 14136
rect 175148 14096 302240 14124
rect 175148 14084 175154 14096
rect 302234 14084 302240 14096
rect 302292 14084 302298 14136
rect 173710 14016 173716 14068
rect 173768 14056 173774 14068
rect 298094 14056 298100 14068
rect 173768 14028 298100 14056
rect 173768 14016 173774 14028
rect 298094 14016 298100 14028
rect 298152 14016 298158 14068
rect 170950 13948 170956 14000
rect 171008 13988 171014 14000
rect 293954 13988 293960 14000
rect 171008 13960 293960 13988
rect 171008 13948 171014 13960
rect 293954 13948 293960 13960
rect 294012 13948 294018 14000
rect 172330 13880 172336 13932
rect 172388 13920 172394 13932
rect 295334 13920 295340 13932
rect 172388 13892 295340 13920
rect 172388 13880 172394 13892
rect 295334 13880 295340 13892
rect 295392 13880 295398 13932
rect 168098 13812 168104 13864
rect 168156 13852 168162 13864
rect 287054 13852 287060 13864
rect 168156 13824 287060 13852
rect 168156 13812 168162 13824
rect 287054 13812 287060 13824
rect 287112 13812 287118 13864
rect 212350 13744 212356 13796
rect 212408 13784 212414 13796
rect 402974 13784 402980 13796
rect 212408 13756 402980 13784
rect 212408 13744 212414 13756
rect 402974 13744 402980 13756
rect 403032 13744 403038 13796
rect 216398 13676 216404 13728
rect 216456 13716 216462 13728
rect 414014 13716 414020 13728
rect 216456 13688 414020 13716
rect 216456 13676 216462 13688
rect 414014 13676 414020 13688
rect 414072 13676 414078 13728
rect 220538 13608 220544 13660
rect 220596 13648 220602 13660
rect 425054 13648 425060 13660
rect 220596 13620 425060 13648
rect 220596 13608 220602 13620
rect 425054 13608 425060 13620
rect 425112 13608 425118 13660
rect 256418 13540 256424 13592
rect 256476 13580 256482 13592
rect 517514 13580 517520 13592
rect 256476 13552 517520 13580
rect 256476 13540 256482 13552
rect 517514 13540 517520 13552
rect 517572 13540 517578 13592
rect 257798 13472 257804 13524
rect 257856 13512 257862 13524
rect 520274 13512 520280 13524
rect 257856 13484 520280 13512
rect 257856 13472 257862 13484
rect 520274 13472 520280 13484
rect 520332 13472 520338 13524
rect 259178 13404 259184 13456
rect 259236 13444 259242 13456
rect 524414 13444 524420 13456
rect 259236 13416 524420 13444
rect 259236 13404 259242 13416
rect 524414 13404 524420 13416
rect 524472 13404 524478 13456
rect 260558 13336 260564 13388
rect 260616 13376 260622 13388
rect 528554 13376 528560 13388
rect 260616 13348 528560 13376
rect 260616 13336 260622 13348
rect 528554 13336 528560 13348
rect 528612 13336 528618 13388
rect 261938 13268 261944 13320
rect 261996 13308 262002 13320
rect 531314 13308 531320 13320
rect 261996 13280 531320 13308
rect 261996 13268 262002 13280
rect 531314 13268 531320 13280
rect 531372 13268 531378 13320
rect 261846 13200 261852 13252
rect 261904 13240 261910 13252
rect 535454 13240 535460 13252
rect 261904 13212 535460 13240
rect 261904 13200 261910 13212
rect 535454 13200 535460 13212
rect 535512 13200 535518 13252
rect 263318 13132 263324 13184
rect 263376 13172 263382 13184
rect 538214 13172 538220 13184
rect 263376 13144 538220 13172
rect 263376 13132 263382 13144
rect 538214 13132 538220 13144
rect 538272 13132 538278 13184
rect 124398 13064 124404 13116
rect 124456 13104 124462 13116
rect 125318 13104 125324 13116
rect 124456 13076 125324 13104
rect 124456 13064 124462 13076
rect 125318 13064 125324 13076
rect 125376 13064 125382 13116
rect 264698 13064 264704 13116
rect 264756 13104 264762 13116
rect 542354 13104 542360 13116
rect 264756 13076 542360 13104
rect 264756 13064 264762 13076
rect 542354 13064 542360 13076
rect 542412 13064 542418 13116
rect 208210 12996 208216 13048
rect 208268 13036 208274 13048
rect 391934 13036 391940 13048
rect 208268 13008 391940 13036
rect 208268 12996 208274 13008
rect 391934 12996 391940 13008
rect 391992 12996 391998 13048
rect 205358 12928 205364 12980
rect 205416 12968 205422 12980
rect 385034 12968 385040 12980
rect 205416 12940 385040 12968
rect 205416 12928 205422 12940
rect 385034 12928 385040 12940
rect 385092 12928 385098 12980
rect 203978 12860 203984 12912
rect 204036 12900 204042 12912
rect 378134 12900 378140 12912
rect 204036 12872 378140 12900
rect 204036 12860 204042 12872
rect 378134 12860 378140 12872
rect 378192 12860 378198 12912
rect 202598 12792 202604 12844
rect 202656 12832 202662 12844
rect 373994 12832 374000 12844
rect 202656 12804 374000 12832
rect 202656 12792 202662 12804
rect 373994 12792 374000 12804
rect 374052 12792 374058 12844
rect 201218 12724 201224 12776
rect 201276 12764 201282 12776
rect 371234 12764 371240 12776
rect 201276 12736 371240 12764
rect 201276 12724 201282 12736
rect 371234 12724 371240 12736
rect 371292 12724 371298 12776
rect 198458 12656 198464 12708
rect 198516 12696 198522 12708
rect 364334 12696 364340 12708
rect 198516 12668 364340 12696
rect 198516 12656 198522 12668
rect 364334 12656 364340 12668
rect 364392 12656 364398 12708
rect 195698 12588 195704 12640
rect 195756 12628 195762 12640
rect 356054 12628 356060 12640
rect 195756 12600 356060 12628
rect 195756 12588 195762 12600
rect 356054 12588 356060 12600
rect 356112 12588 356118 12640
rect 192938 12520 192944 12572
rect 192996 12560 193002 12572
rect 349154 12560 349160 12572
rect 192996 12532 349160 12560
rect 192996 12520 193002 12532
rect 349154 12520 349160 12532
rect 349212 12520 349218 12572
rect 134978 12492 134984 12504
rect 134904 12464 134984 12492
rect 134904 12436 134932 12464
rect 134978 12452 134984 12464
rect 135036 12452 135042 12504
rect 190178 12452 190184 12504
rect 190236 12492 190242 12504
rect 342254 12492 342260 12504
rect 190236 12464 342260 12492
rect 190236 12452 190242 12464
rect 342254 12452 342260 12464
rect 342312 12452 342318 12504
rect 134886 12384 134892 12436
rect 134944 12384 134950 12436
rect 160370 12384 160376 12436
rect 160428 12424 160434 12436
rect 161106 12424 161112 12436
rect 160428 12396 161112 12424
rect 160428 12384 160434 12396
rect 161106 12384 161112 12396
rect 161164 12384 161170 12436
rect 228910 12384 228916 12436
rect 228968 12424 228974 12436
rect 444374 12424 444380 12436
rect 228968 12396 444380 12424
rect 228968 12384 228974 12396
rect 444374 12384 444380 12396
rect 444432 12384 444438 12436
rect 230198 12316 230204 12368
rect 230256 12356 230262 12368
rect 448514 12356 448520 12368
rect 230256 12328 448520 12356
rect 230256 12316 230262 12328
rect 448514 12316 448520 12328
rect 448572 12316 448578 12368
rect 231670 12248 231676 12300
rect 231728 12288 231734 12300
rect 451274 12288 451280 12300
rect 231728 12260 451280 12288
rect 231728 12248 231734 12260
rect 451274 12248 451280 12260
rect 451332 12248 451338 12300
rect 232958 12180 232964 12232
rect 233016 12220 233022 12232
rect 455414 12220 455420 12232
rect 233016 12192 455420 12220
rect 233016 12180 233022 12192
rect 455414 12180 455420 12192
rect 455472 12180 455478 12232
rect 234430 12112 234436 12164
rect 234488 12152 234494 12164
rect 459646 12152 459652 12164
rect 234488 12124 459652 12152
rect 234488 12112 234494 12124
rect 459646 12112 459652 12124
rect 459704 12112 459710 12164
rect 235718 12044 235724 12096
rect 235776 12084 235782 12096
rect 462314 12084 462320 12096
rect 235776 12056 462320 12084
rect 235776 12044 235782 12056
rect 462314 12044 462320 12056
rect 462372 12044 462378 12096
rect 237190 11976 237196 12028
rect 237248 12016 237254 12028
rect 466454 12016 466460 12028
rect 237248 11988 466460 12016
rect 237248 11976 237254 11988
rect 466454 11976 466460 11988
rect 466512 11976 466518 12028
rect 238478 11908 238484 11960
rect 238536 11948 238542 11960
rect 469214 11948 469220 11960
rect 238536 11920 469220 11948
rect 238536 11908 238542 11920
rect 469214 11908 469220 11920
rect 469272 11908 469278 11960
rect 239950 11840 239956 11892
rect 240008 11880 240014 11892
rect 473354 11880 473360 11892
rect 240008 11852 473360 11880
rect 240008 11840 240014 11852
rect 473354 11840 473360 11852
rect 473412 11840 473418 11892
rect 241238 11772 241244 11824
rect 241296 11812 241302 11824
rect 477494 11812 477500 11824
rect 241296 11784 477500 11812
rect 241296 11772 241302 11784
rect 477494 11772 477500 11784
rect 477552 11772 477558 11824
rect 242710 11704 242716 11756
rect 242768 11744 242774 11756
rect 480254 11744 480260 11756
rect 242768 11716 480260 11744
rect 242768 11704 242774 11716
rect 480254 11704 480260 11716
rect 480312 11704 480318 11756
rect 227530 11636 227536 11688
rect 227588 11676 227594 11688
rect 441614 11676 441620 11688
rect 227588 11648 441620 11676
rect 227588 11636 227594 11648
rect 441614 11636 441620 11648
rect 441672 11636 441678 11688
rect 226150 11568 226156 11620
rect 226208 11608 226214 11620
rect 437474 11608 437480 11620
rect 226208 11580 437480 11608
rect 226208 11568 226214 11580
rect 437474 11568 437480 11580
rect 437532 11568 437538 11620
rect 224678 11500 224684 11552
rect 224736 11540 224742 11552
rect 433334 11540 433340 11552
rect 224736 11512 433340 11540
rect 224736 11500 224742 11512
rect 433334 11500 433340 11512
rect 433392 11500 433398 11552
rect 223390 11432 223396 11484
rect 223448 11472 223454 11484
rect 430574 11472 430580 11484
rect 223448 11444 430580 11472
rect 223448 11432 223454 11444
rect 430574 11432 430580 11444
rect 430632 11432 430638 11484
rect 221918 11364 221924 11416
rect 221976 11404 221982 11416
rect 426434 11404 426440 11416
rect 221976 11376 426440 11404
rect 221976 11364 221982 11376
rect 426434 11364 426440 11376
rect 426492 11364 426498 11416
rect 220630 11296 220636 11348
rect 220688 11336 220694 11348
rect 423674 11336 423680 11348
rect 220688 11308 423680 11336
rect 220688 11296 220694 11308
rect 423674 11296 423680 11308
rect 423732 11296 423738 11348
rect 219250 11228 219256 11280
rect 219308 11268 219314 11280
rect 419534 11268 419540 11280
rect 219308 11240 419540 11268
rect 219308 11228 219314 11240
rect 419534 11228 419540 11240
rect 419592 11228 419598 11280
rect 217870 11160 217876 11212
rect 217928 11200 217934 11212
rect 416866 11200 416872 11212
rect 217928 11172 416872 11200
rect 217928 11160 217934 11172
rect 416866 11160 416872 11172
rect 416924 11160 416930 11212
rect 216490 11092 216496 11144
rect 216548 11132 216554 11144
rect 412634 11132 412640 11144
rect 216548 11104 412640 11132
rect 216548 11092 216554 11104
rect 412634 11092 412640 11104
rect 412692 11092 412698 11144
rect 188890 10956 188896 11008
rect 188948 10996 188954 11008
rect 340874 10996 340880 11008
rect 188948 10968 340880 10996
rect 188948 10956 188954 10968
rect 340874 10956 340880 10968
rect 340932 10956 340938 11008
rect 190270 10888 190276 10940
rect 190328 10928 190334 10940
rect 345014 10928 345020 10940
rect 190328 10900 345020 10928
rect 190328 10888 190334 10900
rect 345014 10888 345020 10900
rect 345072 10888 345078 10940
rect 191558 10820 191564 10872
rect 191616 10860 191622 10872
rect 347774 10860 347780 10872
rect 191616 10832 347780 10860
rect 191616 10820 191622 10832
rect 347774 10820 347780 10832
rect 347832 10820 347838 10872
rect 193030 10752 193036 10804
rect 193088 10792 193094 10804
rect 351914 10792 351920 10804
rect 193088 10764 351920 10792
rect 193088 10752 193094 10764
rect 351914 10752 351920 10764
rect 351972 10752 351978 10804
rect 194410 10684 194416 10736
rect 194468 10724 194474 10736
rect 356146 10724 356152 10736
rect 194468 10696 356152 10724
rect 194468 10684 194474 10696
rect 356146 10684 356152 10696
rect 356204 10684 356210 10736
rect 195790 10616 195796 10668
rect 195848 10656 195854 10668
rect 358814 10656 358820 10668
rect 195848 10628 358820 10656
rect 195848 10616 195854 10628
rect 358814 10616 358820 10628
rect 358872 10616 358878 10668
rect 197078 10548 197084 10600
rect 197136 10588 197142 10600
rect 362954 10588 362960 10600
rect 197136 10560 362960 10588
rect 197136 10548 197142 10560
rect 362954 10548 362960 10560
rect 363012 10548 363018 10600
rect 198550 10480 198556 10532
rect 198608 10520 198614 10532
rect 365714 10520 365720 10532
rect 198608 10492 365720 10520
rect 198608 10480 198614 10492
rect 365714 10480 365720 10492
rect 365772 10480 365778 10532
rect 199930 10412 199936 10464
rect 199988 10452 199994 10464
rect 369854 10452 369860 10464
rect 199988 10424 369860 10452
rect 199988 10412 199994 10424
rect 369854 10412 369860 10424
rect 369912 10412 369918 10464
rect 201310 10344 201316 10396
rect 201368 10384 201374 10396
rect 374086 10384 374092 10396
rect 201368 10356 374092 10384
rect 201368 10344 201374 10356
rect 374086 10344 374092 10356
rect 374144 10344 374150 10396
rect 202690 10276 202696 10328
rect 202748 10316 202754 10328
rect 376754 10316 376760 10328
rect 202748 10288 376760 10316
rect 202748 10276 202754 10288
rect 376754 10276 376760 10288
rect 376812 10276 376818 10328
rect 187510 10208 187516 10260
rect 187568 10248 187574 10260
rect 338114 10248 338120 10260
rect 187568 10220 338120 10248
rect 187568 10208 187574 10220
rect 338114 10208 338120 10220
rect 338172 10208 338178 10260
rect 187418 10140 187424 10192
rect 187476 10180 187482 10192
rect 333974 10180 333980 10192
rect 187476 10152 333980 10180
rect 187476 10140 187482 10152
rect 333974 10140 333980 10152
rect 334032 10140 334038 10192
rect 186130 10072 186136 10124
rect 186188 10112 186194 10124
rect 331306 10112 331312 10124
rect 186188 10084 331312 10112
rect 186188 10072 186194 10084
rect 331306 10072 331312 10084
rect 331364 10072 331370 10124
rect 184750 10004 184756 10056
rect 184808 10044 184814 10056
rect 327074 10044 327080 10056
rect 184808 10016 327080 10044
rect 184808 10004 184814 10016
rect 327074 10004 327080 10016
rect 327132 10004 327138 10056
rect 183370 9936 183376 9988
rect 183428 9976 183434 9988
rect 322934 9976 322940 9988
rect 183428 9948 322940 9976
rect 183428 9936 183434 9948
rect 322934 9936 322940 9948
rect 322992 9936 322998 9988
rect 181990 9868 181996 9920
rect 182048 9908 182054 9920
rect 320174 9908 320180 9920
rect 182048 9880 320180 9908
rect 182048 9868 182054 9880
rect 320174 9868 320180 9880
rect 320232 9868 320238 9920
rect 180610 9800 180616 9852
rect 180668 9840 180674 9852
rect 316034 9840 316040 9852
rect 180668 9812 316040 9840
rect 180668 9800 180674 9812
rect 316034 9800 316040 9812
rect 316092 9800 316098 9852
rect 179230 9732 179236 9784
rect 179288 9772 179294 9784
rect 313274 9772 313280 9784
rect 179288 9744 313280 9772
rect 179288 9732 179294 9744
rect 313274 9732 313280 9744
rect 313332 9732 313338 9784
rect 66622 9704 66628 9716
rect 66583 9676 66628 9704
rect 66622 9664 66628 9676
rect 66680 9664 66686 9716
rect 72050 9664 72056 9716
rect 72108 9704 72114 9716
rect 72326 9704 72332 9716
rect 72108 9676 72332 9704
rect 72108 9664 72114 9676
rect 72326 9664 72332 9676
rect 72384 9664 72390 9716
rect 74258 9704 74264 9716
rect 74219 9676 74264 9704
rect 74258 9664 74264 9676
rect 74316 9664 74322 9716
rect 74902 9704 74908 9716
rect 74863 9676 74908 9704
rect 74902 9664 74908 9676
rect 74960 9664 74966 9716
rect 77478 9664 77484 9716
rect 77536 9704 77542 9716
rect 77754 9704 77760 9716
rect 77536 9676 77760 9704
rect 77536 9664 77542 9676
rect 77754 9664 77760 9676
rect 77812 9664 77818 9716
rect 95694 9704 95700 9716
rect 95655 9676 95700 9704
rect 95694 9664 95700 9676
rect 95752 9664 95758 9716
rect 177850 9664 177856 9716
rect 177908 9704 177914 9716
rect 309134 9704 309140 9716
rect 177908 9676 309140 9704
rect 177908 9664 177914 9676
rect 309134 9664 309140 9676
rect 309192 9664 309198 9716
rect 140774 9596 140780 9648
rect 140832 9636 140838 9648
rect 140869 9639 140927 9645
rect 140869 9636 140881 9639
rect 140832 9608 140881 9636
rect 140832 9596 140838 9608
rect 140869 9605 140881 9608
rect 140915 9605 140927 9639
rect 140869 9599 140927 9605
rect 154298 9596 154304 9648
rect 154356 9636 154362 9648
rect 249150 9636 249156 9648
rect 154356 9608 249156 9636
rect 154356 9596 154362 9608
rect 249150 9596 249156 9608
rect 249208 9596 249214 9648
rect 253750 9596 253756 9648
rect 253808 9636 253814 9648
rect 513190 9636 513196 9648
rect 253808 9608 513196 9636
rect 253808 9596 253814 9608
rect 513190 9596 513196 9608
rect 513248 9596 513254 9648
rect 154390 9528 154396 9580
rect 154448 9568 154454 9580
rect 250346 9568 250352 9580
rect 154448 9540 250352 9568
rect 154448 9528 154454 9540
rect 250346 9528 250352 9540
rect 250404 9528 250410 9580
rect 255130 9528 255136 9580
rect 255188 9568 255194 9580
rect 516778 9568 516784 9580
rect 255188 9540 516784 9568
rect 255188 9528 255194 9540
rect 516778 9528 516784 9540
rect 516836 9528 516842 9580
rect 155770 9460 155776 9512
rect 155828 9500 155834 9512
rect 252646 9500 252652 9512
rect 155828 9472 252652 9500
rect 155828 9460 155834 9472
rect 252646 9460 252652 9472
rect 252704 9460 252710 9512
rect 256510 9460 256516 9512
rect 256568 9500 256574 9512
rect 520366 9500 520372 9512
rect 256568 9472 520372 9500
rect 256568 9460 256574 9472
rect 520366 9460 520372 9472
rect 520424 9460 520430 9512
rect 157058 9392 157064 9444
rect 157116 9432 157122 9444
rect 256234 9432 256240 9444
rect 157116 9404 256240 9432
rect 157116 9392 157122 9404
rect 256234 9392 256240 9404
rect 256292 9392 256298 9444
rect 257890 9392 257896 9444
rect 257948 9432 257954 9444
rect 523862 9432 523868 9444
rect 257948 9404 523868 9432
rect 257948 9392 257954 9404
rect 523862 9392 523868 9404
rect 523920 9392 523926 9444
rect 157150 9324 157156 9376
rect 157208 9364 157214 9376
rect 257430 9364 257436 9376
rect 157208 9336 257436 9364
rect 157208 9324 157214 9336
rect 257430 9324 257436 9336
rect 257488 9324 257494 9376
rect 259270 9324 259276 9376
rect 259328 9364 259334 9376
rect 527450 9364 527456 9376
rect 259328 9336 527456 9364
rect 259328 9324 259334 9336
rect 527450 9324 527456 9336
rect 527508 9324 527514 9376
rect 158438 9256 158444 9308
rect 158496 9296 158502 9308
rect 261018 9296 261024 9308
rect 158496 9268 261024 9296
rect 158496 9256 158502 9268
rect 261018 9256 261024 9268
rect 261076 9256 261082 9308
rect 262030 9256 262036 9308
rect 262088 9296 262094 9308
rect 534534 9296 534540 9308
rect 262088 9268 534540 9296
rect 262088 9256 262094 9268
rect 534534 9256 534540 9268
rect 534592 9256 534598 9308
rect 159818 9188 159824 9240
rect 159876 9228 159882 9240
rect 264606 9228 264612 9240
rect 159876 9200 264612 9228
rect 159876 9188 159882 9200
rect 264606 9188 264612 9200
rect 264664 9188 264670 9240
rect 264790 9188 264796 9240
rect 264848 9228 264854 9240
rect 541710 9228 541716 9240
rect 264848 9200 541716 9228
rect 264848 9188 264854 9200
rect 541710 9188 541716 9200
rect 541768 9188 541774 9240
rect 161198 9120 161204 9172
rect 161256 9160 161262 9172
rect 268102 9160 268108 9172
rect 161256 9132 268108 9160
rect 161256 9120 161262 9132
rect 268102 9120 268108 9132
rect 268160 9120 268166 9172
rect 268930 9120 268936 9172
rect 268988 9160 268994 9172
rect 552382 9160 552388 9172
rect 268988 9132 552388 9160
rect 268988 9120 268994 9132
rect 552382 9120 552388 9132
rect 552440 9120 552446 9172
rect 162670 9052 162676 9104
rect 162728 9092 162734 9104
rect 270494 9092 270500 9104
rect 162728 9064 270500 9092
rect 162728 9052 162734 9064
rect 270494 9052 270500 9064
rect 270552 9052 270558 9104
rect 271690 9052 271696 9104
rect 271748 9092 271754 9104
rect 559558 9092 559564 9104
rect 271748 9064 559564 9092
rect 271748 9052 271754 9064
rect 559558 9052 559564 9064
rect 559616 9052 559622 9104
rect 164050 8984 164056 9036
rect 164108 9024 164114 9036
rect 274082 9024 274088 9036
rect 164108 8996 274088 9024
rect 164108 8984 164114 8996
rect 274082 8984 274088 8996
rect 274140 8984 274146 9036
rect 274450 8984 274456 9036
rect 274508 9024 274514 9036
rect 566734 9024 566740 9036
rect 274508 8996 566740 9024
rect 274508 8984 274514 8996
rect 566734 8984 566740 8996
rect 566792 8984 566798 9036
rect 165430 8916 165436 8968
rect 165488 8956 165494 8968
rect 277670 8956 277676 8968
rect 165488 8928 277676 8956
rect 165488 8916 165494 8928
rect 277670 8916 277676 8928
rect 277728 8916 277734 8968
rect 278590 8916 278596 8968
rect 278648 8956 278654 8968
rect 577406 8956 577412 8968
rect 278648 8928 577412 8956
rect 278648 8916 278654 8928
rect 577406 8916 577412 8928
rect 577464 8916 577470 8968
rect 151630 8848 151636 8900
rect 151688 8888 151694 8900
rect 243170 8888 243176 8900
rect 151688 8860 243176 8888
rect 151688 8848 151694 8860
rect 243170 8848 243176 8860
rect 243228 8848 243234 8900
rect 252462 8848 252468 8900
rect 252520 8888 252526 8900
rect 509602 8888 509608 8900
rect 252520 8860 509608 8888
rect 252520 8848 252526 8860
rect 509602 8848 509608 8860
rect 509660 8848 509666 8900
rect 153010 8780 153016 8832
rect 153068 8820 153074 8832
rect 245562 8820 245568 8832
rect 153068 8792 245568 8820
rect 153068 8780 153074 8792
rect 245562 8780 245568 8792
rect 245620 8780 245626 8832
rect 251082 8780 251088 8832
rect 251140 8820 251146 8832
rect 506014 8820 506020 8832
rect 251140 8792 506020 8820
rect 251140 8780 251146 8792
rect 506014 8780 506020 8792
rect 506072 8780 506078 8832
rect 151538 8712 151544 8764
rect 151596 8752 151602 8764
rect 241974 8752 241980 8764
rect 151596 8724 241980 8752
rect 151596 8712 151602 8724
rect 241974 8712 241980 8724
rect 242032 8712 242038 8764
rect 249702 8712 249708 8764
rect 249760 8752 249766 8764
rect 502426 8752 502432 8764
rect 249760 8724 502432 8752
rect 249760 8712 249766 8724
rect 502426 8712 502432 8724
rect 502484 8712 502490 8764
rect 248322 8644 248328 8696
rect 248380 8684 248386 8696
rect 498930 8684 498936 8696
rect 248380 8656 498936 8684
rect 248380 8644 248386 8656
rect 498930 8644 498936 8656
rect 498988 8644 498994 8696
rect 206738 8576 206744 8628
rect 206796 8616 206802 8628
rect 388254 8616 388260 8628
rect 206796 8588 388260 8616
rect 206796 8576 206802 8588
rect 388254 8576 388260 8588
rect 388312 8576 388318 8628
rect 171042 8508 171048 8560
rect 171100 8548 171106 8560
rect 291930 8548 291936 8560
rect 171100 8520 291936 8548
rect 171100 8508 171106 8520
rect 291930 8508 291936 8520
rect 291988 8508 291994 8560
rect 169570 8440 169576 8492
rect 169628 8480 169634 8492
rect 288342 8480 288348 8492
rect 169628 8452 288348 8480
rect 169628 8440 169634 8452
rect 288342 8440 288348 8452
rect 288400 8440 288406 8492
rect 168190 8372 168196 8424
rect 168248 8412 168254 8424
rect 284754 8412 284760 8424
rect 168248 8384 284760 8412
rect 168248 8372 168254 8384
rect 284754 8372 284760 8384
rect 284812 8372 284818 8424
rect 166810 8304 166816 8356
rect 166868 8344 166874 8356
rect 281258 8344 281264 8356
rect 166868 8316 281264 8344
rect 166868 8304 166874 8316
rect 281258 8304 281264 8316
rect 281316 8304 281322 8356
rect 222010 8236 222016 8288
rect 222068 8276 222074 8288
rect 426342 8276 426348 8288
rect 222068 8248 426348 8276
rect 222068 8236 222074 8248
rect 426342 8236 426348 8248
rect 426400 8236 426406 8288
rect 137738 8168 137744 8220
rect 137796 8208 137802 8220
rect 206278 8208 206284 8220
rect 137796 8180 206284 8208
rect 137796 8168 137802 8180
rect 206278 8168 206284 8180
rect 206336 8168 206342 8220
rect 223482 8168 223488 8220
rect 223540 8208 223546 8220
rect 429930 8208 429936 8220
rect 223540 8180 429936 8208
rect 223540 8168 223546 8180
rect 429930 8168 429936 8180
rect 429988 8168 429994 8220
rect 139118 8100 139124 8152
rect 139176 8140 139182 8152
rect 209866 8140 209872 8152
rect 139176 8112 209872 8140
rect 139176 8100 139182 8112
rect 209866 8100 209872 8112
rect 209924 8100 209930 8152
rect 224862 8100 224868 8152
rect 224920 8140 224926 8152
rect 433518 8140 433524 8152
rect 224920 8112 433524 8140
rect 224920 8100 224926 8112
rect 433518 8100 433524 8112
rect 433576 8100 433582 8152
rect 140498 8032 140504 8084
rect 140556 8072 140562 8084
rect 213454 8072 213460 8084
rect 140556 8044 213460 8072
rect 140556 8032 140562 8044
rect 213454 8032 213460 8044
rect 213512 8032 213518 8084
rect 224770 8032 224776 8084
rect 224828 8072 224834 8084
rect 437014 8072 437020 8084
rect 224828 8044 437020 8072
rect 224828 8032 224834 8044
rect 437014 8032 437020 8044
rect 437072 8032 437078 8084
rect 141878 7964 141884 8016
rect 141936 8004 141942 8016
rect 217042 8004 217048 8016
rect 141936 7976 217048 8004
rect 141936 7964 141942 7976
rect 217042 7964 217048 7976
rect 217100 7964 217106 8016
rect 226242 7964 226248 8016
rect 226300 8004 226306 8016
rect 440602 8004 440608 8016
rect 226300 7976 440608 8004
rect 226300 7964 226306 7976
rect 440602 7964 440608 7976
rect 440660 7964 440666 8016
rect 143258 7896 143264 7948
rect 143316 7936 143322 7948
rect 220538 7936 220544 7948
rect 143316 7908 220544 7936
rect 143316 7896 143322 7908
rect 220538 7896 220544 7908
rect 220596 7896 220602 7948
rect 227622 7896 227628 7948
rect 227680 7936 227686 7948
rect 444190 7936 444196 7948
rect 227680 7908 444196 7936
rect 227680 7896 227686 7908
rect 444190 7896 444196 7908
rect 444248 7896 444254 7948
rect 144638 7828 144644 7880
rect 144696 7868 144702 7880
rect 224126 7868 224132 7880
rect 144696 7840 224132 7868
rect 144696 7828 144702 7840
rect 224126 7828 224132 7840
rect 224184 7828 224190 7880
rect 229002 7828 229008 7880
rect 229060 7868 229066 7880
rect 447778 7868 447784 7880
rect 229060 7840 447784 7868
rect 229060 7828 229066 7840
rect 447778 7828 447784 7840
rect 447836 7828 447842 7880
rect 147490 7760 147496 7812
rect 147548 7800 147554 7812
rect 228910 7800 228916 7812
rect 147548 7772 228916 7800
rect 147548 7760 147554 7772
rect 228910 7760 228916 7772
rect 228968 7760 228974 7812
rect 230290 7760 230296 7812
rect 230348 7800 230354 7812
rect 451366 7800 451372 7812
rect 230348 7772 451372 7800
rect 230348 7760 230354 7772
rect 451366 7760 451372 7772
rect 451424 7760 451430 7812
rect 146110 7692 146116 7744
rect 146168 7732 146174 7744
rect 227714 7732 227720 7744
rect 146168 7704 227720 7732
rect 146168 7692 146174 7704
rect 227714 7692 227720 7704
rect 227772 7692 227778 7744
rect 231762 7692 231768 7744
rect 231820 7732 231826 7744
rect 454862 7732 454868 7744
rect 231820 7704 454868 7732
rect 231820 7692 231826 7704
rect 454862 7692 454868 7704
rect 454920 7692 454926 7744
rect 148870 7624 148876 7676
rect 148928 7664 148934 7676
rect 232498 7664 232504 7676
rect 148928 7636 232504 7664
rect 148928 7624 148934 7636
rect 232498 7624 232504 7636
rect 232556 7624 232562 7676
rect 233050 7624 233056 7676
rect 233108 7664 233114 7676
rect 458450 7664 458456 7676
rect 233108 7636 458456 7664
rect 233108 7624 233114 7636
rect 458450 7624 458456 7636
rect 458508 7624 458514 7676
rect 147398 7556 147404 7608
rect 147456 7596 147462 7608
rect 231302 7596 231308 7608
rect 147456 7568 231308 7596
rect 147456 7556 147462 7568
rect 231302 7556 231308 7568
rect 231360 7556 231366 7608
rect 234522 7556 234528 7608
rect 234580 7596 234586 7608
rect 462038 7596 462044 7608
rect 234580 7568 462044 7596
rect 234580 7556 234586 7568
rect 462038 7556 462044 7568
rect 462096 7556 462102 7608
rect 220722 7488 220728 7540
rect 220780 7528 220786 7540
rect 422754 7528 422760 7540
rect 220780 7500 422760 7528
rect 220780 7488 220786 7500
rect 422754 7488 422760 7500
rect 422812 7488 422818 7540
rect 219342 7420 219348 7472
rect 219400 7460 219406 7472
rect 419166 7460 419172 7472
rect 219400 7432 419172 7460
rect 219400 7420 219406 7432
rect 419166 7420 419172 7432
rect 419224 7420 419230 7472
rect 217962 7352 217968 7404
rect 218020 7392 218026 7404
rect 415670 7392 415676 7404
rect 218020 7364 415676 7392
rect 218020 7352 218026 7364
rect 415670 7352 415676 7364
rect 415728 7352 415734 7404
rect 216582 7284 216588 7336
rect 216640 7324 216646 7336
rect 412082 7324 412088 7336
rect 216640 7296 412088 7324
rect 216640 7284 216646 7296
rect 412082 7284 412088 7296
rect 412140 7284 412146 7336
rect 215110 7216 215116 7268
rect 215168 7256 215174 7268
rect 408586 7256 408592 7268
rect 215168 7228 408592 7256
rect 215168 7216 215174 7228
rect 408586 7216 408592 7228
rect 408644 7216 408650 7268
rect 213822 7148 213828 7200
rect 213880 7188 213886 7200
rect 404906 7188 404912 7200
rect 213880 7160 404912 7188
rect 213880 7148 213886 7160
rect 404906 7148 404912 7160
rect 404964 7148 404970 7200
rect 212442 7080 212448 7132
rect 212500 7120 212506 7132
rect 401318 7120 401324 7132
rect 212500 7092 401324 7120
rect 212500 7080 212506 7092
rect 401318 7080 401324 7092
rect 401376 7080 401382 7132
rect 211062 7012 211068 7064
rect 211120 7052 211126 7064
rect 397822 7052 397828 7064
rect 211120 7024 397828 7052
rect 211120 7012 211126 7024
rect 397822 7012 397828 7024
rect 397880 7012 397886 7064
rect 161290 6944 161296 6996
rect 161348 6984 161354 6996
rect 266998 6984 267004 6996
rect 161348 6956 267004 6984
rect 161348 6944 161354 6956
rect 266998 6944 267004 6956
rect 267056 6944 267062 6996
rect 202782 6916 202788 6928
rect 202743 6888 202788 6916
rect 202782 6876 202788 6888
rect 202840 6876 202846 6928
rect 125410 6808 125416 6860
rect 125468 6848 125474 6860
rect 170582 6848 170588 6860
rect 125468 6820 170588 6848
rect 125468 6808 125474 6820
rect 170582 6808 170588 6820
rect 170640 6808 170646 6860
rect 184842 6808 184848 6860
rect 184900 6848 184906 6860
rect 330018 6848 330024 6860
rect 184900 6820 330024 6848
rect 184900 6808 184906 6820
rect 330018 6808 330024 6820
rect 330076 6808 330082 6860
rect 126882 6740 126888 6792
rect 126940 6780 126946 6792
rect 174170 6780 174176 6792
rect 126940 6752 174176 6780
rect 126940 6740 126946 6752
rect 174170 6740 174176 6752
rect 174228 6740 174234 6792
rect 186222 6740 186228 6792
rect 186280 6780 186286 6792
rect 333606 6780 333612 6792
rect 186280 6752 333612 6780
rect 186280 6740 186286 6752
rect 333606 6740 333612 6752
rect 333664 6740 333670 6792
rect 128262 6672 128268 6724
rect 128320 6712 128326 6724
rect 177758 6712 177764 6724
rect 128320 6684 177764 6712
rect 128320 6672 128326 6684
rect 177758 6672 177764 6684
rect 177816 6672 177822 6724
rect 187602 6672 187608 6724
rect 187660 6712 187666 6724
rect 337102 6712 337108 6724
rect 187660 6684 337108 6712
rect 187660 6672 187666 6684
rect 337102 6672 337108 6684
rect 337160 6672 337166 6724
rect 129550 6604 129556 6656
rect 129608 6644 129614 6656
rect 181346 6644 181352 6656
rect 129608 6616 181352 6644
rect 129608 6604 129614 6616
rect 181346 6604 181352 6616
rect 181404 6604 181410 6656
rect 188982 6604 188988 6656
rect 189040 6644 189046 6656
rect 340690 6644 340696 6656
rect 189040 6616 340696 6644
rect 189040 6604 189046 6616
rect 340690 6604 340696 6616
rect 340748 6604 340754 6656
rect 131022 6536 131028 6588
rect 131080 6576 131086 6588
rect 184842 6576 184848 6588
rect 131080 6548 184848 6576
rect 131080 6536 131086 6548
rect 184842 6536 184848 6548
rect 184900 6536 184906 6588
rect 190362 6536 190368 6588
rect 190420 6576 190426 6588
rect 344278 6576 344284 6588
rect 190420 6548 344284 6576
rect 190420 6536 190426 6548
rect 344278 6536 344284 6548
rect 344336 6536 344342 6588
rect 130930 6468 130936 6520
rect 130988 6508 130994 6520
rect 188430 6508 188436 6520
rect 130988 6480 188436 6508
rect 130988 6468 130994 6480
rect 188430 6468 188436 6480
rect 188488 6468 188494 6520
rect 193122 6468 193128 6520
rect 193180 6508 193186 6520
rect 351362 6508 351368 6520
rect 193180 6480 351368 6508
rect 193180 6468 193186 6480
rect 351362 6468 351368 6480
rect 351420 6468 351426 6520
rect 132310 6400 132316 6452
rect 132368 6440 132374 6452
rect 192018 6440 192024 6452
rect 132368 6412 192024 6440
rect 132368 6400 132374 6412
rect 192018 6400 192024 6412
rect 192076 6400 192082 6452
rect 194502 6400 194508 6452
rect 194560 6440 194566 6452
rect 354950 6440 354956 6452
rect 194560 6412 354956 6440
rect 194560 6400 194566 6412
rect 354950 6400 354956 6412
rect 355008 6400 355014 6452
rect 133690 6332 133696 6384
rect 133748 6372 133754 6384
rect 195606 6372 195612 6384
rect 133748 6344 195612 6372
rect 133748 6332 133754 6344
rect 195606 6332 195612 6344
rect 195664 6332 195670 6384
rect 195882 6332 195888 6384
rect 195940 6372 195946 6384
rect 358538 6372 358544 6384
rect 195940 6344 358544 6372
rect 195940 6332 195946 6344
rect 358538 6332 358544 6344
rect 358596 6332 358602 6384
rect 134886 6264 134892 6316
rect 134944 6304 134950 6316
rect 199194 6304 199200 6316
rect 134944 6276 199200 6304
rect 134944 6264 134950 6276
rect 199194 6264 199200 6276
rect 199252 6264 199258 6316
rect 200022 6264 200028 6316
rect 200080 6304 200086 6316
rect 369210 6304 369216 6316
rect 200080 6276 369216 6304
rect 200080 6264 200086 6276
rect 369210 6264 369216 6276
rect 369268 6264 369274 6316
rect 158530 6196 158536 6248
rect 158588 6236 158594 6248
rect 259822 6236 259828 6248
rect 158588 6208 259828 6236
rect 158588 6196 158594 6208
rect 259822 6196 259828 6208
rect 259880 6196 259886 6248
rect 273070 6196 273076 6248
rect 273128 6236 273134 6248
rect 563146 6236 563152 6248
rect 273128 6208 563152 6236
rect 273128 6196 273134 6208
rect 563146 6196 563152 6208
rect 563204 6196 563210 6248
rect 159910 6128 159916 6180
rect 159968 6168 159974 6180
rect 263410 6168 263416 6180
rect 159968 6140 263416 6168
rect 159968 6128 159974 6140
rect 263410 6128 263416 6140
rect 263468 6128 263474 6180
rect 277210 6128 277216 6180
rect 277268 6168 277274 6180
rect 573818 6168 573824 6180
rect 277268 6140 573824 6168
rect 277268 6128 277274 6140
rect 573818 6128 573824 6140
rect 573876 6128 573882 6180
rect 123938 6060 123944 6112
rect 123996 6100 124002 6112
rect 167086 6100 167092 6112
rect 123996 6072 167092 6100
rect 123996 6060 124002 6072
rect 167086 6060 167092 6072
rect 167144 6060 167150 6112
rect 175918 6060 175924 6112
rect 175976 6100 175982 6112
rect 181533 6103 181591 6109
rect 181533 6100 181545 6103
rect 175976 6072 181545 6100
rect 175976 6060 175982 6072
rect 181533 6069 181545 6072
rect 181579 6069 181591 6103
rect 181533 6063 181591 6069
rect 183462 6060 183468 6112
rect 183520 6100 183526 6112
rect 326430 6100 326436 6112
rect 183520 6072 326436 6100
rect 183520 6060 183526 6072
rect 326430 6060 326436 6072
rect 326488 6060 326494 6112
rect 122650 5992 122656 6044
rect 122708 6032 122714 6044
rect 163498 6032 163504 6044
rect 122708 6004 163504 6032
rect 122708 5992 122714 6004
rect 163498 5992 163504 6004
rect 163556 5992 163562 6044
rect 182082 5992 182088 6044
rect 182140 6032 182146 6044
rect 322842 6032 322848 6044
rect 182140 6004 322848 6032
rect 182140 5992 182146 6004
rect 322842 5992 322848 6004
rect 322900 5992 322906 6044
rect 180702 5924 180708 5976
rect 180760 5964 180766 5976
rect 319254 5964 319260 5976
rect 180760 5936 319260 5964
rect 180760 5924 180766 5936
rect 319254 5924 319260 5936
rect 319312 5924 319318 5976
rect 179322 5856 179328 5908
rect 179380 5896 179386 5908
rect 315758 5896 315764 5908
rect 179380 5868 315764 5896
rect 179380 5856 179386 5868
rect 315758 5856 315764 5868
rect 315816 5856 315822 5908
rect 177942 5788 177948 5840
rect 178000 5828 178006 5840
rect 312170 5828 312176 5840
rect 178000 5800 312176 5828
rect 178000 5788 178006 5800
rect 312170 5788 312176 5800
rect 312228 5788 312234 5840
rect 176562 5720 176568 5772
rect 176620 5760 176626 5772
rect 308582 5760 308588 5772
rect 176620 5732 308588 5760
rect 176620 5720 176626 5732
rect 308582 5720 308588 5732
rect 308640 5720 308646 5772
rect 175182 5652 175188 5704
rect 175240 5692 175246 5704
rect 305086 5692 305092 5704
rect 175240 5664 305092 5692
rect 175240 5652 175246 5664
rect 305086 5652 305092 5664
rect 305144 5652 305150 5704
rect 173802 5584 173808 5636
rect 173860 5624 173866 5636
rect 301406 5624 301412 5636
rect 173860 5596 301412 5624
rect 173860 5584 173866 5596
rect 301406 5584 301412 5596
rect 301464 5584 301470 5636
rect 172422 5516 172428 5568
rect 172480 5556 172486 5568
rect 297910 5556 297916 5568
rect 172480 5528 297916 5556
rect 172480 5516 172486 5528
rect 297910 5516 297916 5528
rect 297968 5516 297974 5568
rect 148962 5448 148968 5500
rect 149020 5488 149026 5500
rect 233694 5488 233700 5500
rect 149020 5460 233700 5488
rect 149020 5448 149026 5460
rect 233694 5448 233700 5460
rect 233752 5448 233758 5500
rect 262122 5448 262128 5500
rect 262180 5488 262186 5500
rect 533430 5488 533436 5500
rect 262180 5460 533436 5488
rect 262180 5448 262186 5460
rect 533430 5448 533436 5460
rect 533488 5448 533494 5500
rect 150158 5380 150164 5432
rect 150216 5420 150222 5432
rect 237190 5420 237196 5432
rect 150216 5392 237196 5420
rect 150216 5380 150222 5392
rect 237190 5380 237196 5392
rect 237248 5380 237254 5432
rect 263502 5380 263508 5432
rect 263560 5420 263566 5432
rect 536926 5420 536932 5432
rect 263560 5392 536932 5420
rect 263560 5380 263566 5392
rect 536926 5380 536932 5392
rect 536984 5380 536990 5432
rect 151722 5312 151728 5364
rect 151780 5352 151786 5364
rect 240778 5352 240784 5364
rect 151780 5324 240784 5352
rect 151780 5312 151786 5324
rect 240778 5312 240784 5324
rect 240836 5312 240842 5364
rect 264882 5312 264888 5364
rect 264940 5352 264946 5364
rect 540514 5352 540520 5364
rect 264940 5324 540520 5352
rect 264940 5312 264946 5324
rect 540514 5312 540520 5324
rect 540572 5312 540578 5364
rect 153102 5244 153108 5296
rect 153160 5284 153166 5296
rect 244366 5284 244372 5296
rect 153160 5256 244372 5284
rect 153160 5244 153166 5256
rect 244366 5244 244372 5256
rect 244424 5244 244430 5296
rect 266262 5244 266268 5296
rect 266320 5284 266326 5296
rect 544102 5284 544108 5296
rect 266320 5256 544108 5284
rect 266320 5244 266326 5256
rect 544102 5244 544108 5256
rect 544160 5244 544166 5296
rect 66257 5219 66315 5225
rect 66257 5185 66269 5219
rect 66303 5216 66315 5219
rect 71866 5216 71872 5228
rect 66303 5188 71872 5216
rect 66303 5185 66315 5188
rect 66257 5179 66315 5185
rect 71866 5176 71872 5188
rect 71924 5176 71930 5228
rect 154482 5176 154488 5228
rect 154540 5216 154546 5228
rect 247954 5216 247960 5228
rect 154540 5188 247960 5216
rect 154540 5176 154546 5188
rect 247954 5176 247960 5188
rect 248012 5176 248018 5228
rect 267642 5176 267648 5228
rect 267700 5216 267706 5228
rect 547690 5216 547696 5228
rect 267700 5188 547696 5216
rect 267700 5176 267706 5188
rect 547690 5176 547696 5188
rect 547748 5176 547754 5228
rect 155862 5108 155868 5160
rect 155920 5148 155926 5160
rect 251450 5148 251456 5160
rect 155920 5120 251456 5148
rect 155920 5108 155926 5120
rect 251450 5108 251456 5120
rect 251508 5108 251514 5160
rect 269022 5108 269028 5160
rect 269080 5148 269086 5160
rect 551186 5148 551192 5160
rect 269080 5120 551192 5148
rect 269080 5108 269086 5120
rect 551186 5108 551192 5120
rect 551244 5108 551250 5160
rect 157242 5040 157248 5092
rect 157300 5080 157306 5092
rect 255038 5080 255044 5092
rect 157300 5052 255044 5080
rect 157300 5040 157306 5052
rect 255038 5040 255044 5052
rect 255096 5040 255102 5092
rect 270402 5040 270408 5092
rect 270460 5080 270466 5092
rect 554774 5080 554780 5092
rect 270460 5052 554780 5080
rect 270460 5040 270466 5052
rect 554774 5040 554780 5052
rect 554832 5040 554838 5092
rect 158622 4972 158628 5024
rect 158680 5012 158686 5024
rect 258626 5012 258632 5024
rect 158680 4984 258632 5012
rect 158680 4972 158686 4984
rect 258626 4972 258632 4984
rect 258684 4972 258690 5024
rect 271782 4972 271788 5024
rect 271840 5012 271846 5024
rect 558362 5012 558368 5024
rect 271840 4984 558368 5012
rect 271840 4972 271846 4984
rect 558362 4972 558368 4984
rect 558420 4972 558426 5024
rect 160002 4904 160008 4956
rect 160060 4944 160066 4956
rect 262214 4944 262220 4956
rect 160060 4916 262220 4944
rect 160060 4904 160066 4916
rect 262214 4904 262220 4916
rect 262272 4904 262278 4956
rect 273162 4904 273168 4956
rect 273220 4944 273226 4956
rect 561950 4944 561956 4956
rect 273220 4916 561956 4944
rect 273220 4904 273226 4916
rect 561950 4904 561956 4916
rect 562008 4904 562014 4956
rect 161382 4836 161388 4888
rect 161440 4876 161446 4888
rect 265802 4876 265808 4888
rect 161440 4848 265808 4876
rect 161440 4836 161446 4848
rect 265802 4836 265808 4848
rect 265860 4836 265866 4888
rect 274542 4836 274548 4888
rect 274600 4876 274606 4888
rect 565538 4876 565544 4888
rect 274600 4848 565544 4876
rect 274600 4836 274606 4848
rect 565538 4836 565544 4848
rect 565596 4836 565602 4888
rect 55214 4768 55220 4820
rect 55272 4808 55278 4820
rect 80422 4808 80428 4820
rect 55272 4780 80428 4808
rect 55272 4768 55278 4780
rect 80422 4768 80428 4780
rect 80480 4768 80486 4820
rect 86957 4811 87015 4817
rect 86957 4777 86969 4811
rect 87003 4808 87015 4811
rect 90358 4808 90364 4820
rect 87003 4780 90364 4808
rect 87003 4777 87015 4780
rect 86957 4771 87015 4777
rect 90358 4768 90364 4780
rect 90416 4768 90422 4820
rect 162762 4768 162768 4820
rect 162820 4808 162826 4820
rect 269298 4808 269304 4820
rect 162820 4780 269304 4808
rect 162820 4768 162826 4780
rect 269298 4768 269304 4780
rect 269356 4768 269362 4820
rect 275922 4768 275928 4820
rect 275980 4808 275986 4820
rect 569034 4808 569040 4820
rect 275980 4780 569040 4808
rect 275980 4768 275986 4780
rect 569034 4768 569040 4780
rect 569092 4768 569098 4820
rect 147582 4700 147588 4752
rect 147640 4740 147646 4752
rect 230106 4740 230112 4752
rect 147640 4712 230112 4740
rect 147640 4700 147646 4712
rect 230106 4700 230112 4712
rect 230164 4700 230170 4752
rect 260742 4700 260748 4752
rect 260800 4740 260806 4752
rect 529842 4740 529848 4752
rect 260800 4712 529848 4740
rect 260800 4700 260806 4712
rect 529842 4700 529848 4712
rect 529900 4700 529906 4752
rect 146202 4632 146208 4684
rect 146260 4672 146266 4684
rect 226518 4672 226524 4684
rect 146260 4644 226524 4672
rect 146260 4632 146266 4644
rect 226518 4632 226524 4644
rect 226576 4632 226582 4684
rect 259362 4632 259368 4684
rect 259420 4672 259426 4684
rect 526254 4672 526260 4684
rect 259420 4644 526260 4672
rect 259420 4632 259426 4644
rect 526254 4632 526260 4644
rect 526312 4632 526318 4684
rect 144730 4564 144736 4616
rect 144788 4604 144794 4616
rect 222930 4604 222936 4616
rect 144788 4576 222936 4604
rect 144788 4564 144794 4576
rect 222930 4564 222936 4576
rect 222988 4564 222994 4616
rect 257982 4564 257988 4616
rect 258040 4604 258046 4616
rect 522666 4604 522672 4616
rect 258040 4576 522672 4604
rect 258040 4564 258046 4576
rect 522666 4564 522672 4576
rect 522724 4564 522730 4616
rect 143350 4496 143356 4548
rect 143408 4536 143414 4548
rect 219342 4536 219348 4548
rect 143408 4508 219348 4536
rect 143408 4496 143414 4508
rect 219342 4496 219348 4508
rect 219400 4496 219406 4548
rect 256602 4496 256608 4548
rect 256660 4536 256666 4548
rect 519078 4536 519084 4548
rect 256660 4508 519084 4536
rect 256660 4496 256666 4508
rect 519078 4496 519084 4508
rect 519136 4496 519142 4548
rect 141970 4428 141976 4480
rect 142028 4468 142034 4480
rect 215846 4468 215852 4480
rect 142028 4440 215852 4468
rect 142028 4428 142034 4440
rect 215846 4428 215852 4440
rect 215904 4428 215910 4480
rect 255222 4428 255228 4480
rect 255280 4468 255286 4480
rect 515582 4468 515588 4480
rect 255280 4440 515588 4468
rect 255280 4428 255286 4440
rect 515582 4428 515588 4440
rect 515640 4428 515646 4480
rect 140590 4360 140596 4412
rect 140648 4400 140654 4412
rect 212258 4400 212264 4412
rect 140648 4372 212264 4400
rect 140648 4360 140654 4372
rect 212258 4360 212264 4372
rect 212316 4360 212322 4412
rect 253842 4360 253848 4412
rect 253900 4400 253906 4412
rect 511994 4400 512000 4412
rect 253900 4372 512000 4400
rect 253900 4360 253906 4372
rect 511994 4360 512000 4372
rect 512052 4360 512058 4412
rect 139210 4292 139216 4344
rect 139268 4332 139274 4344
rect 208670 4332 208676 4344
rect 139268 4304 208676 4332
rect 139268 4292 139274 4304
rect 208670 4292 208676 4304
rect 208728 4292 208734 4344
rect 209590 4292 209596 4344
rect 209648 4332 209654 4344
rect 394234 4332 394240 4344
rect 209648 4304 394240 4332
rect 209648 4292 209654 4304
rect 394234 4292 394240 4304
rect 394292 4292 394298 4344
rect 66625 4267 66683 4273
rect 66625 4233 66637 4267
rect 66671 4264 66683 4267
rect 70578 4264 70584 4276
rect 66671 4236 70584 4264
rect 66671 4233 66683 4236
rect 66625 4227 66683 4233
rect 70578 4224 70584 4236
rect 70636 4224 70642 4276
rect 137830 4224 137836 4276
rect 137888 4264 137894 4276
rect 205082 4264 205088 4276
rect 137888 4236 205088 4264
rect 137888 4224 137894 4236
rect 205082 4224 205088 4236
rect 205140 4224 205146 4276
rect 205542 4224 205548 4276
rect 205600 4264 205606 4276
rect 383562 4264 383568 4276
rect 205600 4236 383568 4264
rect 205600 4224 205606 4236
rect 383562 4224 383568 4236
rect 383620 4224 383626 4276
rect 55217 4199 55275 4205
rect 55217 4165 55229 4199
rect 55263 4196 55275 4199
rect 60921 4199 60979 4205
rect 55263 4168 60872 4196
rect 55263 4165 55275 4168
rect 55217 4159 55275 4165
rect 37366 4088 37372 4140
rect 37424 4128 37430 4140
rect 38562 4128 38568 4140
rect 37424 4100 38568 4128
rect 37424 4088 37430 4100
rect 38562 4088 38568 4100
rect 38620 4088 38626 4140
rect 40681 4131 40739 4137
rect 40681 4097 40693 4131
rect 40727 4128 40739 4131
rect 60737 4131 60795 4137
rect 60737 4128 60749 4131
rect 40727 4100 60749 4128
rect 40727 4097 40739 4100
rect 40681 4091 40739 4097
rect 60737 4097 60749 4100
rect 60783 4097 60795 4131
rect 60844 4128 60872 4168
rect 60921 4165 60933 4199
rect 60967 4196 60979 4199
rect 66257 4199 66315 4205
rect 66257 4196 66269 4199
rect 60967 4168 66269 4196
rect 60967 4165 60979 4168
rect 60921 4159 60979 4165
rect 66257 4165 66269 4168
rect 66303 4165 66315 4199
rect 75365 4199 75423 4205
rect 75365 4196 75377 4199
rect 66257 4159 66315 4165
rect 70412 4168 75377 4196
rect 70412 4137 70440 4168
rect 75365 4165 75377 4168
rect 75411 4165 75423 4199
rect 75365 4159 75423 4165
rect 119890 4156 119896 4208
rect 119948 4196 119954 4208
rect 122009 4199 122067 4205
rect 122009 4196 122021 4199
rect 119948 4168 122021 4196
rect 119948 4156 119954 4168
rect 122009 4165 122021 4168
rect 122055 4165 122067 4199
rect 122009 4159 122067 4165
rect 136542 4156 136548 4208
rect 136600 4196 136606 4208
rect 201494 4196 201500 4208
rect 136600 4168 201500 4196
rect 136600 4156 136606 4168
rect 201494 4156 201500 4168
rect 201552 4156 201558 4208
rect 202785 4199 202843 4205
rect 202785 4165 202797 4199
rect 202831 4196 202843 4199
rect 376386 4196 376392 4208
rect 202831 4168 376392 4196
rect 202831 4165 202843 4168
rect 202785 4159 202843 4165
rect 376386 4156 376392 4168
rect 376444 4156 376450 4208
rect 66625 4131 66683 4137
rect 66625 4128 66637 4131
rect 60844 4100 66637 4128
rect 60737 4091 60795 4097
rect 66625 4097 66637 4100
rect 66671 4097 66683 4131
rect 66625 4091 66683 4097
rect 70397 4131 70455 4137
rect 70397 4097 70409 4131
rect 70443 4097 70455 4131
rect 70397 4091 70455 4097
rect 72142 4088 72148 4140
rect 72200 4128 72206 4140
rect 75178 4128 75184 4140
rect 72200 4100 75184 4128
rect 72200 4088 72206 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 75288 4100 80192 4128
rect 29086 4020 29092 4072
rect 29144 4060 29150 4072
rect 30282 4060 30288 4072
rect 29144 4032 30288 4060
rect 29144 4020 29150 4032
rect 30282 4020 30288 4032
rect 30340 4020 30346 4072
rect 30377 4063 30435 4069
rect 30377 4029 30389 4063
rect 30423 4060 30435 4063
rect 35897 4063 35955 4069
rect 35897 4060 35909 4063
rect 30423 4032 35909 4060
rect 30423 4029 30435 4032
rect 30377 4023 30435 4029
rect 35897 4029 35909 4032
rect 35943 4029 35955 4063
rect 35897 4023 35955 4029
rect 45465 4063 45523 4069
rect 45465 4029 45477 4063
rect 45511 4060 45523 4063
rect 55217 4063 55275 4069
rect 55217 4060 55229 4063
rect 45511 4032 55229 4060
rect 45511 4029 45523 4032
rect 45465 4023 45523 4029
rect 55217 4029 55229 4032
rect 55263 4029 55275 4063
rect 55217 4023 55275 4029
rect 75089 4063 75147 4069
rect 75089 4029 75101 4063
rect 75135 4060 75147 4063
rect 75288 4060 75316 4100
rect 75135 4032 75316 4060
rect 75365 4063 75423 4069
rect 75135 4029 75147 4032
rect 75089 4023 75147 4029
rect 75365 4029 75377 4063
rect 75411 4060 75423 4063
rect 78766 4060 78772 4072
rect 75411 4032 78772 4060
rect 75411 4029 75423 4032
rect 75365 4023 75423 4029
rect 78766 4020 78772 4032
rect 78824 4020 78830 4072
rect 79042 4020 79048 4072
rect 79100 4060 79106 4072
rect 80057 4063 80115 4069
rect 80057 4060 80069 4063
rect 79100 4032 80069 4060
rect 79100 4020 79106 4032
rect 80057 4029 80069 4032
rect 80103 4029 80115 4063
rect 80164 4060 80192 4100
rect 80238 4088 80244 4140
rect 80296 4128 80302 4140
rect 82078 4128 82084 4140
rect 80296 4100 82084 4128
rect 80296 4088 80302 4100
rect 82078 4088 82084 4100
rect 82136 4088 82142 4140
rect 83826 4088 83832 4140
rect 83884 4128 83890 4140
rect 84838 4128 84844 4140
rect 83884 4100 84844 4128
rect 83884 4088 83890 4100
rect 84838 4088 84844 4100
rect 84896 4088 84902 4140
rect 84930 4088 84936 4140
rect 84988 4128 84994 4140
rect 85482 4128 85488 4140
rect 84988 4100 85488 4128
rect 84988 4088 84994 4100
rect 85482 4088 85488 4100
rect 85540 4088 85546 4140
rect 88518 4088 88524 4140
rect 88576 4128 88582 4140
rect 89622 4128 89628 4140
rect 88576 4100 89628 4128
rect 88576 4088 88582 4100
rect 89622 4088 89628 4100
rect 89680 4088 89686 4140
rect 93302 4088 93308 4140
rect 93360 4128 93366 4140
rect 93762 4128 93768 4140
rect 93360 4100 93768 4128
rect 93360 4088 93366 4100
rect 93762 4088 93768 4100
rect 93820 4088 93826 4140
rect 96522 4088 96528 4140
rect 96580 4128 96586 4140
rect 96890 4128 96896 4140
rect 96580 4100 96896 4128
rect 96580 4088 96586 4100
rect 96890 4088 96896 4100
rect 96948 4088 96954 4140
rect 97902 4088 97908 4140
rect 97960 4128 97966 4140
rect 99282 4128 99288 4140
rect 97960 4100 99288 4128
rect 97960 4088 97966 4100
rect 99282 4088 99288 4100
rect 99340 4088 99346 4140
rect 100018 4088 100024 4140
rect 100076 4128 100082 4140
rect 103974 4128 103980 4140
rect 100076 4100 103980 4128
rect 100076 4088 100082 4100
rect 103974 4088 103980 4100
rect 104032 4088 104038 4140
rect 104618 4088 104624 4140
rect 104676 4128 104682 4140
rect 117130 4128 117136 4140
rect 104676 4100 117136 4128
rect 104676 4088 104682 4100
rect 117130 4088 117136 4100
rect 117188 4088 117194 4140
rect 117222 4088 117228 4140
rect 117280 4128 117286 4140
rect 148229 4131 148287 4137
rect 148229 4128 148241 4131
rect 117280 4100 148241 4128
rect 117280 4088 117286 4100
rect 148229 4097 148241 4100
rect 148275 4097 148287 4131
rect 148229 4091 148287 4097
rect 148318 4088 148324 4140
rect 148376 4128 148382 4140
rect 151538 4128 151544 4140
rect 148376 4100 151544 4128
rect 148376 4088 148382 4100
rect 151538 4088 151544 4100
rect 151596 4088 151602 4140
rect 152458 4088 152464 4140
rect 152516 4128 152522 4140
rect 155126 4128 155132 4140
rect 152516 4100 155132 4128
rect 152516 4088 152522 4100
rect 155126 4088 155132 4100
rect 155184 4088 155190 4140
rect 155218 4088 155224 4140
rect 155276 4128 155282 4140
rect 162029 4131 162087 4137
rect 155276 4100 161980 4128
rect 155276 4088 155282 4100
rect 82906 4060 82912 4072
rect 80164 4032 82912 4060
rect 80057 4023 80115 4029
rect 82906 4020 82912 4032
rect 82964 4020 82970 4072
rect 104802 4020 104808 4072
rect 104860 4060 104866 4072
rect 118234 4060 118240 4072
rect 104860 4032 118240 4060
rect 104860 4020 104866 4032
rect 118234 4020 118240 4032
rect 118292 4020 118298 4072
rect 118510 4020 118516 4072
rect 118568 4060 118574 4072
rect 143445 4063 143503 4069
rect 143445 4060 143457 4063
rect 118568 4032 143457 4060
rect 118568 4020 118574 4032
rect 143445 4029 143457 4032
rect 143491 4029 143503 4063
rect 143445 4023 143503 4029
rect 153838 4020 153844 4072
rect 153896 4060 153902 4072
rect 161952 4069 161980 4100
rect 162029 4097 162041 4131
rect 162075 4128 162087 4131
rect 187053 4131 187111 4137
rect 162075 4100 187004 4128
rect 162075 4097 162087 4100
rect 162029 4091 162087 4097
rect 161845 4063 161903 4069
rect 161845 4060 161857 4063
rect 153896 4032 161857 4060
rect 153896 4020 153902 4032
rect 161845 4029 161857 4032
rect 161891 4029 161903 4063
rect 161845 4023 161903 4029
rect 161937 4063 161995 4069
rect 161937 4029 161949 4063
rect 161983 4029 161995 4063
rect 161937 4023 161995 4029
rect 162121 4063 162179 4069
rect 162121 4029 162133 4063
rect 162167 4060 162179 4063
rect 162167 4032 186544 4060
rect 162167 4029 162179 4032
rect 162121 4023 162179 4029
rect 25498 3952 25504 4004
rect 25556 3992 25562 4004
rect 69106 3992 69112 4004
rect 25556 3964 69112 3992
rect 25556 3952 25562 3964
rect 69106 3952 69112 3964
rect 69164 3952 69170 4004
rect 69201 3995 69259 4001
rect 69201 3961 69213 3995
rect 69247 3992 69259 3995
rect 72050 3992 72056 4004
rect 69247 3964 72056 3992
rect 69247 3961 69259 3964
rect 69201 3955 69259 3961
rect 72050 3952 72056 3964
rect 72108 3952 72114 4004
rect 73062 3952 73068 4004
rect 73120 3992 73126 4004
rect 79318 3992 79324 4004
rect 73120 3964 79324 3992
rect 73120 3952 73126 3964
rect 79318 3952 79324 3964
rect 79376 3952 79382 4004
rect 79413 3995 79471 4001
rect 79413 3961 79425 3995
rect 79459 3992 79471 3995
rect 85574 3992 85580 4004
rect 79459 3964 85580 3992
rect 79459 3961 79471 3964
rect 79413 3955 79471 3961
rect 85574 3952 85580 3964
rect 85632 3952 85638 4004
rect 106090 3952 106096 4004
rect 106148 3992 106154 4004
rect 120626 3992 120632 4004
rect 106148 3964 120632 3992
rect 106148 3952 106154 3964
rect 120626 3952 120632 3964
rect 120684 3952 120690 4004
rect 121270 3952 121276 4004
rect 121328 3992 121334 4004
rect 159910 3992 159916 4004
rect 121328 3964 159916 3992
rect 121328 3952 121334 3964
rect 159910 3952 159916 3964
rect 159968 3952 159974 4004
rect 167638 3952 167644 4004
rect 167696 3992 167702 4004
rect 167696 3964 168328 3992
rect 167696 3952 167702 3964
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 66622 3924 66628 3936
rect 18380 3896 66628 3924
rect 18380 3884 18386 3896
rect 66622 3884 66628 3896
rect 66680 3884 66686 3936
rect 67174 3884 67180 3936
rect 67232 3924 67238 3936
rect 74169 3927 74227 3933
rect 74169 3924 74181 3927
rect 67232 3896 74181 3924
rect 67232 3884 67238 3896
rect 74169 3893 74181 3896
rect 74215 3893 74227 3927
rect 75273 3927 75331 3933
rect 75273 3924 75285 3927
rect 74169 3887 74227 3893
rect 74276 3896 75285 3924
rect 16022 3816 16028 3868
rect 16080 3856 16086 3868
rect 64874 3856 64880 3868
rect 16080 3828 64880 3856
rect 16080 3816 16086 3828
rect 64874 3816 64880 3828
rect 64932 3816 64938 3868
rect 74276 3856 74304 3896
rect 75273 3893 75285 3896
rect 75319 3893 75331 3927
rect 75273 3887 75331 3893
rect 75454 3884 75460 3936
rect 75512 3924 75518 3936
rect 81253 3927 81311 3933
rect 81253 3924 81265 3927
rect 75512 3896 81265 3924
rect 75512 3884 75518 3896
rect 81253 3893 81265 3896
rect 81299 3893 81311 3927
rect 81253 3887 81311 3893
rect 81345 3927 81403 3933
rect 81345 3893 81357 3927
rect 81391 3924 81403 3927
rect 85758 3924 85764 3936
rect 81391 3896 85764 3924
rect 81391 3893 81403 3896
rect 81345 3887 81403 3893
rect 85758 3884 85764 3896
rect 85816 3884 85822 3936
rect 107562 3884 107568 3936
rect 107620 3924 107626 3936
rect 120813 3927 120871 3933
rect 120813 3924 120825 3927
rect 107620 3896 120825 3924
rect 107620 3884 107626 3896
rect 120813 3893 120825 3896
rect 120859 3893 120871 3927
rect 124214 3924 124220 3936
rect 120813 3887 120871 3893
rect 121932 3896 124220 3924
rect 65076 3828 74304 3856
rect 74353 3859 74411 3865
rect 14826 3748 14832 3800
rect 14884 3788 14890 3800
rect 64966 3788 64972 3800
rect 14884 3760 64972 3788
rect 14884 3748 14890 3760
rect 64966 3748 64972 3760
rect 65024 3748 65030 3800
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 63586 3720 63592 3732
rect 10100 3692 63592 3720
rect 10100 3680 10106 3692
rect 63586 3680 63592 3692
rect 63644 3680 63650 3732
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 62206 3652 62212 3664
rect 7708 3624 62212 3652
rect 7708 3612 7714 3624
rect 62206 3612 62212 3624
rect 62264 3612 62270 3664
rect 62390 3612 62396 3664
rect 62448 3652 62454 3664
rect 65076 3652 65104 3828
rect 74353 3825 74365 3859
rect 74399 3856 74411 3859
rect 77938 3856 77944 3868
rect 74399 3828 77944 3856
rect 74399 3825 74411 3828
rect 74353 3819 74411 3825
rect 77938 3816 77944 3828
rect 77996 3816 78002 3868
rect 80057 3859 80115 3865
rect 80057 3825 80069 3859
rect 80103 3856 80115 3859
rect 87598 3856 87604 3868
rect 80103 3828 87604 3856
rect 80103 3825 80115 3828
rect 80057 3819 80115 3825
rect 87598 3816 87604 3828
rect 87656 3816 87662 3868
rect 89714 3816 89720 3868
rect 89772 3856 89778 3868
rect 92566 3856 92572 3868
rect 89772 3828 92572 3856
rect 89772 3816 89778 3828
rect 92566 3816 92572 3828
rect 92624 3816 92630 3868
rect 94498 3816 94504 3868
rect 94556 3856 94562 3868
rect 95326 3856 95332 3868
rect 94556 3828 95332 3856
rect 94556 3816 94562 3828
rect 95326 3816 95332 3828
rect 95384 3816 95390 3868
rect 106182 3816 106188 3868
rect 106240 3856 106246 3868
rect 121822 3856 121828 3868
rect 106240 3828 121828 3856
rect 106240 3816 106246 3828
rect 121822 3816 121828 3828
rect 121880 3816 121886 3868
rect 68278 3748 68284 3800
rect 68336 3788 68342 3800
rect 75273 3791 75331 3797
rect 68336 3760 75224 3788
rect 68336 3748 68342 3760
rect 65153 3723 65211 3729
rect 65153 3689 65165 3723
rect 65199 3720 65211 3723
rect 75089 3723 75147 3729
rect 75089 3720 75101 3723
rect 65199 3692 75101 3720
rect 65199 3689 65211 3692
rect 65153 3683 65211 3689
rect 75089 3689 75101 3692
rect 75135 3689 75147 3723
rect 75196 3720 75224 3760
rect 75273 3757 75285 3791
rect 75319 3788 75331 3791
rect 79410 3788 79416 3800
rect 75319 3760 79416 3788
rect 75319 3757 75331 3760
rect 75273 3751 75331 3757
rect 79410 3748 79416 3760
rect 79468 3748 79474 3800
rect 79505 3791 79563 3797
rect 79505 3757 79517 3791
rect 79551 3788 79563 3791
rect 81894 3788 81900 3800
rect 79551 3760 81900 3788
rect 79551 3757 79563 3760
rect 79505 3751 79563 3757
rect 81894 3748 81900 3760
rect 81952 3748 81958 3800
rect 107470 3748 107476 3800
rect 107528 3788 107534 3800
rect 121932 3788 121960 3896
rect 124214 3884 124220 3896
rect 124272 3884 124278 3936
rect 125502 3884 125508 3936
rect 125560 3924 125566 3936
rect 133141 3927 133199 3933
rect 133141 3924 133153 3927
rect 125560 3896 133153 3924
rect 125560 3884 125566 3896
rect 133141 3893 133153 3896
rect 133187 3893 133199 3927
rect 133141 3887 133199 3893
rect 133233 3927 133291 3933
rect 133233 3893 133245 3927
rect 133279 3924 133291 3927
rect 137465 3927 137523 3933
rect 137465 3924 137477 3927
rect 133279 3896 137477 3924
rect 133279 3893 133291 3896
rect 133233 3887 133291 3893
rect 137465 3893 137477 3896
rect 137511 3893 137523 3927
rect 137465 3887 137523 3893
rect 137557 3927 137615 3933
rect 137557 3893 137569 3927
rect 137603 3924 137615 3927
rect 168190 3924 168196 3936
rect 137603 3896 168196 3924
rect 137603 3893 137615 3896
rect 137557 3887 137615 3893
rect 168190 3884 168196 3896
rect 168248 3884 168254 3936
rect 168300 3924 168328 3964
rect 169018 3952 169024 4004
rect 169076 3992 169082 4004
rect 176470 3992 176476 4004
rect 169076 3964 176476 3992
rect 169076 3952 169082 3964
rect 176470 3952 176476 3964
rect 176528 3952 176534 4004
rect 176565 3995 176623 4001
rect 176565 3961 176577 3995
rect 176611 3992 176623 3995
rect 176657 3995 176715 4001
rect 176657 3992 176669 3995
rect 176611 3964 176669 3992
rect 176611 3961 176623 3964
rect 176565 3955 176623 3961
rect 176657 3961 176669 3964
rect 176703 3961 176715 3995
rect 182542 3992 182548 4004
rect 176657 3955 176715 3961
rect 176764 3964 182548 3992
rect 169849 3927 169907 3933
rect 169849 3924 169861 3927
rect 168300 3896 169861 3924
rect 169849 3893 169861 3896
rect 169895 3893 169907 3927
rect 169849 3887 169907 3893
rect 169938 3884 169944 3936
rect 169996 3924 170002 3936
rect 172974 3924 172980 3936
rect 169996 3896 172980 3924
rect 169996 3884 170002 3896
rect 172974 3884 172980 3896
rect 173032 3884 173038 3936
rect 176764 3924 176792 3964
rect 182542 3952 182548 3964
rect 182600 3952 182606 4004
rect 182637 3995 182695 4001
rect 182637 3961 182649 3995
rect 182683 3992 182695 3995
rect 186225 3995 186283 4001
rect 186225 3992 186237 3995
rect 182683 3964 186237 3992
rect 182683 3961 182695 3964
rect 182637 3955 182695 3961
rect 186225 3961 186237 3964
rect 186271 3961 186283 3995
rect 186516 3992 186544 4032
rect 186777 3995 186835 4001
rect 186777 3992 186789 3995
rect 186516 3964 186789 3992
rect 186225 3955 186283 3961
rect 186777 3961 186789 3964
rect 186823 3961 186835 3995
rect 186976 3992 187004 4100
rect 187053 4097 187065 4131
rect 187099 4128 187111 4131
rect 300302 4128 300308 4140
rect 187099 4100 300308 4128
rect 187099 4097 187111 4100
rect 187053 4091 187111 4097
rect 300302 4088 300308 4100
rect 300360 4088 300366 4140
rect 304258 4088 304264 4140
rect 304316 4128 304322 4140
rect 307386 4128 307392 4140
rect 304316 4100 307392 4128
rect 304316 4088 304322 4100
rect 307386 4088 307392 4100
rect 307444 4088 307450 4140
rect 187237 4063 187295 4069
rect 187237 4029 187249 4063
rect 187283 4060 187295 4063
rect 193214 4060 193220 4072
rect 187283 4032 193220 4060
rect 187283 4029 187295 4032
rect 187237 4023 187295 4029
rect 193214 4020 193220 4032
rect 193272 4020 193278 4072
rect 310974 4060 310980 4072
rect 193324 4032 310980 4060
rect 190822 3992 190828 4004
rect 186976 3964 190828 3992
rect 186777 3955 186835 3961
rect 190822 3952 190828 3964
rect 190880 3952 190886 4004
rect 190917 3995 190975 4001
rect 190917 3961 190929 3995
rect 190963 3992 190975 3995
rect 193125 3995 193183 4001
rect 193125 3992 193137 3995
rect 190963 3964 193137 3992
rect 190963 3961 190975 3964
rect 190917 3955 190975 3961
rect 193125 3961 193137 3964
rect 193171 3961 193183 3995
rect 193125 3955 193183 3961
rect 176672 3896 176792 3924
rect 122742 3816 122748 3868
rect 122800 3856 122806 3868
rect 159361 3859 159419 3865
rect 159361 3856 159373 3859
rect 122800 3828 159373 3856
rect 122800 3816 122806 3828
rect 159361 3825 159373 3828
rect 159407 3825 159419 3859
rect 159361 3819 159419 3825
rect 159450 3816 159456 3868
rect 159508 3856 159514 3868
rect 164694 3856 164700 3868
rect 159508 3828 164700 3856
rect 159508 3816 159514 3828
rect 164694 3816 164700 3828
rect 164752 3816 164758 3868
rect 166258 3816 166264 3868
rect 166316 3856 166322 3868
rect 176562 3856 176568 3868
rect 166316 3828 176568 3856
rect 166316 3816 166322 3828
rect 176562 3816 176568 3828
rect 176620 3816 176626 3868
rect 107528 3760 121960 3788
rect 122009 3791 122067 3797
rect 107528 3748 107534 3760
rect 122009 3757 122021 3791
rect 122055 3788 122067 3791
rect 123297 3791 123355 3797
rect 123297 3788 123309 3791
rect 122055 3760 123309 3788
rect 122055 3757 122067 3760
rect 122009 3751 122067 3757
rect 123297 3757 123309 3760
rect 123343 3757 123355 3791
rect 131390 3788 131396 3800
rect 123297 3751 123355 3757
rect 123404 3760 131396 3788
rect 81345 3723 81403 3729
rect 81345 3720 81357 3723
rect 75196 3692 81357 3720
rect 75089 3683 75147 3689
rect 81345 3689 81357 3692
rect 81391 3689 81403 3723
rect 81345 3683 81403 3689
rect 81434 3680 81440 3732
rect 81492 3720 81498 3732
rect 82722 3720 82728 3732
rect 81492 3692 82728 3720
rect 81492 3680 81498 3692
rect 82722 3680 82728 3692
rect 82780 3680 82786 3732
rect 104710 3680 104716 3732
rect 104768 3720 104774 3732
rect 104768 3692 108896 3720
rect 104768 3680 104774 3692
rect 62448 3624 65104 3652
rect 62448 3612 62454 3624
rect 65978 3612 65984 3664
rect 66036 3652 66042 3664
rect 84286 3652 84292 3664
rect 66036 3624 84292 3652
rect 66036 3612 66042 3624
rect 84286 3612 84292 3624
rect 84344 3612 84350 3664
rect 102778 3612 102784 3664
rect 102836 3652 102842 3664
rect 108758 3652 108764 3664
rect 102836 3624 108764 3652
rect 102836 3612 102842 3624
rect 108758 3612 108764 3624
rect 108816 3612 108822 3664
rect 108868 3652 108896 3692
rect 108942 3680 108948 3732
rect 109000 3720 109006 3732
rect 120721 3723 120779 3729
rect 120721 3720 120733 3723
rect 109000 3692 120733 3720
rect 109000 3680 109006 3692
rect 120721 3689 120733 3692
rect 120767 3689 120779 3723
rect 120721 3683 120779 3689
rect 120813 3723 120871 3729
rect 120813 3689 120825 3723
rect 120859 3720 120871 3723
rect 123018 3720 123024 3732
rect 120859 3692 123024 3720
rect 120859 3689 120871 3692
rect 120813 3683 120871 3689
rect 123018 3680 123024 3692
rect 123076 3680 123082 3732
rect 108868 3624 110092 3652
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 62114 3584 62120 3596
rect 6512 3556 62120 3584
rect 6512 3544 6518 3556
rect 62114 3544 62120 3556
rect 62172 3544 62178 3596
rect 63586 3544 63592 3596
rect 63644 3584 63650 3596
rect 64693 3587 64751 3593
rect 64693 3584 64705 3587
rect 63644 3556 64705 3584
rect 63644 3544 63650 3556
rect 64693 3553 64705 3556
rect 64739 3553 64751 3587
rect 64693 3547 64751 3553
rect 64782 3544 64788 3596
rect 64840 3584 64846 3596
rect 84378 3584 84384 3596
rect 64840 3556 84384 3584
rect 64840 3544 64846 3556
rect 84378 3544 84384 3556
rect 84436 3544 84442 3596
rect 87322 3544 87328 3596
rect 87380 3584 87386 3596
rect 88242 3584 88248 3596
rect 87380 3556 88248 3584
rect 87380 3544 87386 3556
rect 88242 3544 88248 3556
rect 88300 3544 88306 3596
rect 100662 3544 100668 3596
rect 100720 3584 100726 3596
rect 106366 3584 106372 3596
rect 100720 3556 106372 3584
rect 100720 3544 100726 3556
rect 106366 3544 106372 3556
rect 106424 3544 106430 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 59354 3516 59360 3528
rect 1728 3488 59360 3516
rect 1728 3476 1734 3488
rect 59354 3476 59360 3488
rect 59412 3476 59418 3528
rect 59998 3476 60004 3528
rect 60056 3516 60062 3528
rect 60056 3488 75224 3516
rect 60056 3476 60062 3488
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 59906 3448 59912 3460
rect 624 3420 59912 3448
rect 624 3408 630 3420
rect 59906 3408 59912 3420
rect 59964 3408 59970 3460
rect 61194 3408 61200 3460
rect 61252 3448 61258 3460
rect 75089 3451 75147 3457
rect 75089 3448 75101 3451
rect 61252 3420 75101 3448
rect 61252 3408 61258 3420
rect 75089 3417 75101 3420
rect 75135 3417 75147 3451
rect 75196 3448 75224 3488
rect 76650 3476 76656 3528
rect 76708 3516 76714 3528
rect 82170 3516 82176 3528
rect 76708 3488 82176 3516
rect 76708 3476 76714 3488
rect 82170 3476 82176 3488
rect 82228 3476 82234 3528
rect 100110 3476 100116 3528
rect 100168 3516 100174 3528
rect 101582 3516 101588 3528
rect 100168 3488 101588 3516
rect 100168 3476 100174 3488
rect 101582 3476 101588 3488
rect 101640 3476 101646 3528
rect 101950 3476 101956 3528
rect 102008 3516 102014 3528
rect 109954 3516 109960 3528
rect 102008 3488 109960 3516
rect 102008 3476 102014 3488
rect 109954 3476 109960 3488
rect 110012 3476 110018 3528
rect 110064 3516 110092 3624
rect 110138 3612 110144 3664
rect 110196 3652 110202 3664
rect 123404 3652 123432 3760
rect 131390 3748 131396 3760
rect 131448 3748 131454 3800
rect 133049 3791 133107 3797
rect 133049 3788 133061 3791
rect 131500 3760 133061 3788
rect 124122 3680 124128 3732
rect 124180 3720 124186 3732
rect 126701 3723 126759 3729
rect 126701 3720 126713 3723
rect 124180 3692 126713 3720
rect 124180 3680 124186 3692
rect 126701 3689 126713 3692
rect 126747 3689 126759 3723
rect 126701 3683 126759 3689
rect 127618 3680 127624 3732
rect 127676 3720 127682 3732
rect 131301 3723 131359 3729
rect 131301 3720 131313 3723
rect 127676 3692 131313 3720
rect 127676 3680 127682 3692
rect 131301 3689 131313 3692
rect 131347 3689 131359 3723
rect 131301 3683 131359 3689
rect 110196 3624 123432 3652
rect 123481 3655 123539 3661
rect 110196 3612 110202 3624
rect 123481 3621 123493 3655
rect 123527 3652 123539 3655
rect 127897 3655 127955 3661
rect 127897 3652 127909 3655
rect 123527 3624 127909 3652
rect 123527 3621 123539 3624
rect 123481 3615 123539 3621
rect 127897 3621 127909 3624
rect 127943 3621 127955 3655
rect 127897 3615 127955 3621
rect 130378 3612 130384 3664
rect 130436 3652 130442 3664
rect 131500 3652 131528 3760
rect 133049 3757 133061 3760
rect 133095 3757 133107 3791
rect 133049 3751 133107 3757
rect 133141 3791 133199 3797
rect 133141 3757 133153 3791
rect 133187 3788 133199 3791
rect 169938 3788 169944 3800
rect 133187 3760 169944 3788
rect 133187 3757 133199 3760
rect 133141 3751 133199 3757
rect 169938 3748 169944 3760
rect 169996 3748 170002 3800
rect 170033 3791 170091 3797
rect 170033 3757 170045 3791
rect 170079 3788 170091 3791
rect 171689 3791 171747 3797
rect 171689 3788 171701 3791
rect 170079 3760 171701 3788
rect 170079 3757 170091 3760
rect 170033 3751 170091 3757
rect 171689 3757 171701 3760
rect 171735 3757 171747 3791
rect 176672 3788 176700 3896
rect 176838 3884 176844 3936
rect 176896 3924 176902 3936
rect 189353 3927 189411 3933
rect 189353 3924 189365 3927
rect 176896 3896 189365 3924
rect 176896 3884 176902 3896
rect 189353 3893 189365 3896
rect 189399 3893 189411 3927
rect 189353 3887 189411 3893
rect 189810 3884 189816 3936
rect 189868 3924 189874 3936
rect 193324 3924 193352 4032
rect 310974 4020 310980 4032
rect 311032 4020 311038 4072
rect 193401 3995 193459 4001
rect 193401 3961 193413 3995
rect 193447 3992 193459 3995
rect 289538 3992 289544 4004
rect 193447 3964 289544 3992
rect 193447 3961 193459 3964
rect 193401 3955 193459 3961
rect 289538 3952 289544 3964
rect 289596 3952 289602 4004
rect 295978 3952 295984 4004
rect 296036 3992 296042 4004
rect 417970 3992 417976 4004
rect 296036 3964 417976 3992
rect 296036 3952 296042 3964
rect 417970 3952 417976 3964
rect 418028 3952 418034 4004
rect 332410 3924 332416 3936
rect 189868 3896 193352 3924
rect 193416 3896 332416 3924
rect 189868 3884 189874 3896
rect 176746 3816 176752 3868
rect 176804 3856 176810 3868
rect 190917 3859 190975 3865
rect 190917 3856 190929 3859
rect 176804 3828 190929 3856
rect 176804 3816 176810 3828
rect 190917 3825 190929 3828
rect 190963 3825 190975 3859
rect 193416 3856 193444 3896
rect 332410 3884 332416 3896
rect 332468 3884 332474 3936
rect 190917 3819 190975 3825
rect 191024 3828 193444 3856
rect 181441 3791 181499 3797
rect 181441 3788 181453 3791
rect 171689 3751 171747 3757
rect 171796 3760 176700 3788
rect 176764 3760 181453 3788
rect 131577 3723 131635 3729
rect 131577 3689 131589 3723
rect 131623 3720 131635 3723
rect 133782 3720 133788 3732
rect 131623 3692 133788 3720
rect 131623 3689 131635 3692
rect 131577 3683 131635 3689
rect 133782 3680 133788 3692
rect 133840 3680 133846 3732
rect 133877 3723 133935 3729
rect 133877 3689 133889 3723
rect 133923 3720 133935 3723
rect 148229 3723 148287 3729
rect 148229 3720 148241 3723
rect 133923 3692 148241 3720
rect 133923 3689 133935 3692
rect 133877 3683 133935 3689
rect 148229 3689 148241 3692
rect 148275 3689 148287 3723
rect 148229 3683 148287 3689
rect 148321 3723 148379 3729
rect 148321 3689 148333 3723
rect 148367 3720 148379 3723
rect 150434 3720 150440 3732
rect 148367 3692 150440 3720
rect 148367 3689 148379 3692
rect 148321 3683 148379 3689
rect 150434 3680 150440 3692
rect 150492 3680 150498 3732
rect 151078 3680 151084 3732
rect 151136 3720 151142 3732
rect 156509 3723 156567 3729
rect 156509 3720 156521 3723
rect 151136 3692 156521 3720
rect 151136 3680 151142 3692
rect 156509 3689 156521 3692
rect 156555 3689 156567 3723
rect 156509 3683 156567 3689
rect 157978 3680 157984 3732
rect 158036 3720 158042 3732
rect 162029 3723 162087 3729
rect 162029 3720 162041 3723
rect 158036 3692 162041 3720
rect 158036 3680 158042 3692
rect 162029 3689 162041 3692
rect 162075 3689 162087 3723
rect 162029 3683 162087 3689
rect 162121 3723 162179 3729
rect 162121 3689 162133 3723
rect 162167 3720 162179 3723
rect 171796 3720 171824 3760
rect 162167 3692 171824 3720
rect 171873 3723 171931 3729
rect 162167 3689 162179 3692
rect 162121 3683 162179 3689
rect 171873 3689 171885 3723
rect 171919 3720 171931 3723
rect 175921 3723 175979 3729
rect 175921 3720 175933 3723
rect 171919 3692 175933 3720
rect 171919 3689 171931 3692
rect 171873 3683 171931 3689
rect 175921 3689 175933 3692
rect 175967 3689 175979 3723
rect 175921 3683 175979 3689
rect 176010 3680 176016 3732
rect 176068 3720 176074 3732
rect 176764 3720 176792 3760
rect 181441 3757 181453 3760
rect 181487 3757 181499 3791
rect 181441 3751 181499 3757
rect 181530 3748 181536 3800
rect 181588 3788 181594 3800
rect 185489 3791 185547 3797
rect 185489 3788 185501 3791
rect 181588 3760 185501 3788
rect 181588 3748 181594 3760
rect 185489 3757 185501 3760
rect 185535 3757 185547 3791
rect 185489 3751 185547 3757
rect 185578 3748 185584 3800
rect 185636 3788 185642 3800
rect 187053 3791 187111 3797
rect 187053 3788 187065 3791
rect 185636 3760 187065 3788
rect 185636 3748 185642 3760
rect 187053 3757 187065 3760
rect 187099 3757 187111 3791
rect 187053 3751 187111 3757
rect 187145 3791 187203 3797
rect 187145 3757 187157 3791
rect 187191 3788 187203 3791
rect 190365 3791 190423 3797
rect 190365 3788 190377 3791
rect 187191 3760 190377 3788
rect 187191 3757 187203 3760
rect 187145 3751 187203 3757
rect 190365 3757 190377 3760
rect 190411 3757 190423 3791
rect 190365 3751 190423 3757
rect 190454 3748 190460 3800
rect 190512 3788 190518 3800
rect 191024 3788 191052 3828
rect 193858 3816 193864 3868
rect 193916 3856 193922 3868
rect 335906 3856 335912 3868
rect 193916 3828 335912 3856
rect 193916 3816 193922 3828
rect 335906 3816 335912 3828
rect 335964 3816 335970 3868
rect 190512 3760 191052 3788
rect 190512 3748 190518 3760
rect 191742 3748 191748 3800
rect 191800 3788 191806 3800
rect 346670 3788 346676 3800
rect 191800 3760 346676 3788
rect 191800 3748 191806 3760
rect 346670 3748 346676 3760
rect 346728 3748 346734 3800
rect 360930 3788 360936 3800
rect 355980 3760 360936 3788
rect 176068 3692 176792 3720
rect 176068 3680 176074 3692
rect 176930 3680 176936 3732
rect 176988 3720 176994 3732
rect 183738 3720 183744 3732
rect 176988 3692 183744 3720
rect 176988 3680 176994 3692
rect 183738 3680 183744 3692
rect 183796 3680 183802 3732
rect 184198 3680 184204 3732
rect 184256 3720 184262 3732
rect 190825 3723 190883 3729
rect 190825 3720 190837 3723
rect 184256 3692 190837 3720
rect 184256 3680 184262 3692
rect 190825 3689 190837 3692
rect 190871 3689 190883 3723
rect 190825 3683 190883 3689
rect 191101 3723 191159 3729
rect 191101 3689 191113 3723
rect 191147 3720 191159 3723
rect 200390 3720 200396 3732
rect 191147 3692 200396 3720
rect 191147 3689 191159 3692
rect 191101 3683 191159 3689
rect 200390 3680 200396 3692
rect 200448 3680 200454 3732
rect 355980 3720 356008 3760
rect 360930 3748 360936 3760
rect 360988 3748 360994 3800
rect 201144 3692 356008 3720
rect 130436 3624 131528 3652
rect 130436 3612 130442 3624
rect 132402 3612 132408 3664
rect 132460 3652 132466 3664
rect 132460 3624 132724 3652
rect 132460 3612 132466 3624
rect 110230 3544 110236 3596
rect 110288 3584 110294 3596
rect 132586 3584 132592 3596
rect 110288 3556 132592 3584
rect 110288 3544 110294 3556
rect 132586 3544 132592 3556
rect 132644 3544 132650 3596
rect 132696 3584 132724 3624
rect 133138 3612 133144 3664
rect 133196 3652 133202 3664
rect 137278 3652 137284 3664
rect 133196 3624 137284 3652
rect 133196 3612 133202 3624
rect 137278 3612 137284 3624
rect 137336 3612 137342 3664
rect 189626 3652 189632 3664
rect 137388 3624 189632 3652
rect 137388 3584 137416 3624
rect 189626 3612 189632 3624
rect 189684 3612 189690 3664
rect 189718 3612 189724 3664
rect 189776 3652 189782 3664
rect 190270 3652 190276 3664
rect 189776 3624 190276 3652
rect 189776 3612 189782 3624
rect 190270 3612 190276 3624
rect 190328 3612 190334 3664
rect 190365 3655 190423 3661
rect 190365 3621 190377 3655
rect 190411 3652 190423 3655
rect 194410 3652 194416 3664
rect 190411 3624 194416 3652
rect 190411 3621 190423 3624
rect 190365 3615 190423 3621
rect 194410 3612 194416 3624
rect 194468 3612 194474 3664
rect 197262 3612 197268 3664
rect 197320 3652 197326 3664
rect 201144 3652 201172 3692
rect 356054 3680 356060 3732
rect 356112 3720 356118 3732
rect 357342 3720 357348 3732
rect 356112 3692 357348 3720
rect 356112 3680 356118 3692
rect 357342 3680 357348 3692
rect 357400 3680 357406 3732
rect 373994 3680 374000 3732
rect 374052 3720 374058 3732
rect 375190 3720 375196 3732
rect 374052 3692 375196 3720
rect 374052 3680 374058 3692
rect 375190 3680 375196 3692
rect 375248 3680 375254 3732
rect 197320 3624 201172 3652
rect 197320 3612 197326 3624
rect 206922 3612 206928 3664
rect 206980 3652 206986 3664
rect 389450 3652 389456 3664
rect 206980 3624 389456 3652
rect 206980 3612 206986 3624
rect 389450 3612 389456 3624
rect 389508 3612 389514 3664
rect 132696 3556 137416 3584
rect 137465 3587 137523 3593
rect 137465 3553 137477 3587
rect 137511 3584 137523 3587
rect 141789 3587 141847 3593
rect 141789 3584 141801 3587
rect 137511 3556 141801 3584
rect 137511 3553 137523 3556
rect 137465 3547 137523 3553
rect 141789 3553 141801 3556
rect 141835 3553 141847 3587
rect 141789 3547 141847 3553
rect 141881 3587 141939 3593
rect 141881 3553 141893 3587
rect 141927 3584 141939 3587
rect 186317 3587 186375 3593
rect 186317 3584 186329 3587
rect 141927 3556 186329 3584
rect 141927 3553 141939 3556
rect 141881 3547 141939 3553
rect 186317 3553 186329 3556
rect 186363 3553 186375 3587
rect 186317 3547 186375 3553
rect 186406 3544 186412 3596
rect 186464 3584 186470 3596
rect 187234 3584 187240 3596
rect 186464 3556 187240 3584
rect 186464 3544 186470 3556
rect 187234 3544 187240 3556
rect 187292 3544 187298 3596
rect 189353 3587 189411 3593
rect 189353 3553 189365 3587
rect 189399 3584 189411 3587
rect 196802 3584 196808 3596
rect 189399 3556 196808 3584
rect 189399 3553 189411 3556
rect 189353 3547 189411 3553
rect 196802 3544 196808 3556
rect 196860 3544 196866 3596
rect 209682 3544 209688 3596
rect 209740 3584 209746 3596
rect 396626 3584 396632 3596
rect 209740 3556 396632 3584
rect 209740 3544 209746 3556
rect 396626 3544 396632 3556
rect 396684 3544 396690 3596
rect 408494 3544 408500 3596
rect 408552 3584 408558 3596
rect 409690 3584 409696 3596
rect 408552 3556 409696 3584
rect 408552 3544 408558 3556
rect 409690 3544 409696 3556
rect 409748 3544 409754 3596
rect 485774 3544 485780 3596
rect 485832 3584 485838 3596
rect 486970 3584 486976 3596
rect 485832 3556 486976 3584
rect 485832 3544 485838 3556
rect 486970 3544 486976 3556
rect 487028 3544 487034 3596
rect 110064 3488 111288 3516
rect 81526 3448 81532 3460
rect 75196 3420 81532 3448
rect 75089 3411 75147 3417
rect 81526 3408 81532 3420
rect 81584 3408 81590 3460
rect 82630 3408 82636 3460
rect 82688 3448 82694 3460
rect 86957 3451 87015 3457
rect 86957 3448 86969 3451
rect 82688 3420 86969 3448
rect 82688 3408 82694 3420
rect 86957 3417 86969 3420
rect 87003 3417 87015 3451
rect 86957 3411 87015 3417
rect 97810 3408 97816 3460
rect 97868 3448 97874 3460
rect 100478 3448 100484 3460
rect 97868 3420 100484 3448
rect 97868 3408 97874 3420
rect 100478 3408 100484 3420
rect 100536 3408 100542 3460
rect 102042 3408 102048 3460
rect 102100 3448 102106 3460
rect 111150 3448 111156 3460
rect 102100 3420 111156 3448
rect 102100 3408 102106 3420
rect 111150 3408 111156 3420
rect 111208 3408 111214 3460
rect 111260 3448 111288 3488
rect 111702 3476 111708 3528
rect 111760 3516 111766 3528
rect 136082 3516 136088 3528
rect 111760 3488 136088 3516
rect 111760 3476 111766 3488
rect 136082 3476 136088 3488
rect 136140 3476 136146 3528
rect 137922 3476 137928 3528
rect 137980 3516 137986 3528
rect 203886 3516 203892 3528
rect 137980 3488 203892 3516
rect 137980 3476 137986 3488
rect 203886 3476 203892 3488
rect 203944 3476 203950 3528
rect 215202 3476 215208 3528
rect 215260 3516 215266 3528
rect 410886 3516 410892 3528
rect 215260 3488 410892 3516
rect 215260 3476 215266 3488
rect 410886 3476 410892 3488
rect 410944 3476 410950 3528
rect 433334 3476 433340 3528
rect 433392 3516 433398 3528
rect 434622 3516 434628 3528
rect 433392 3488 434628 3516
rect 433392 3476 433398 3488
rect 434622 3476 434628 3488
rect 434680 3476 434686 3528
rect 451274 3476 451280 3528
rect 451332 3516 451338 3528
rect 452470 3516 452476 3528
rect 451332 3488 452476 3516
rect 451332 3476 451338 3488
rect 452470 3476 452476 3488
rect 452528 3476 452534 3528
rect 459554 3476 459560 3528
rect 459612 3516 459618 3528
rect 460842 3516 460848 3528
rect 459612 3488 460848 3516
rect 459612 3476 459618 3488
rect 460842 3476 460848 3488
rect 460900 3476 460906 3528
rect 502334 3476 502340 3528
rect 502392 3516 502398 3528
rect 503622 3516 503628 3528
rect 502392 3488 503628 3516
rect 502392 3476 502398 3488
rect 503622 3476 503628 3488
rect 503680 3476 503686 3528
rect 520274 3476 520280 3528
rect 520332 3516 520338 3528
rect 521470 3516 521476 3528
rect 520332 3488 521476 3516
rect 520332 3476 520338 3488
rect 521470 3476 521476 3488
rect 521528 3476 521534 3528
rect 529474 3476 529480 3528
rect 529532 3516 529538 3528
rect 564342 3516 564348 3528
rect 529532 3488 564348 3516
rect 529532 3476 529538 3488
rect 564342 3476 564348 3488
rect 564400 3476 564406 3528
rect 111260 3420 112576 3448
rect 11238 3340 11244 3392
rect 11296 3380 11302 3392
rect 12342 3380 12348 3392
rect 11296 3352 12348 3380
rect 11296 3340 11302 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 17862 3380 17868 3392
rect 17276 3352 17868 3380
rect 17276 3340 17282 3352
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 20622 3380 20628 3392
rect 19576 3352 20628 3380
rect 19576 3340 19582 3352
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 26694 3340 26700 3392
rect 26752 3380 26758 3392
rect 27522 3380 27528 3392
rect 26752 3352 27528 3380
rect 26752 3340 26758 3352
rect 27522 3340 27528 3352
rect 27580 3340 27586 3392
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 30377 3383 30435 3389
rect 30377 3380 30389 3383
rect 27948 3352 30389 3380
rect 27948 3340 27954 3352
rect 30377 3349 30389 3352
rect 30423 3349 30435 3383
rect 30377 3343 30435 3349
rect 33870 3340 33876 3392
rect 33928 3380 33934 3392
rect 65705 3383 65763 3389
rect 33928 3352 65656 3380
rect 33928 3340 33934 3352
rect 32674 3272 32680 3324
rect 32732 3312 32738 3324
rect 32732 3284 36124 3312
rect 32732 3272 32738 3284
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 13722 3176 13728 3188
rect 12492 3148 13728 3176
rect 12492 3136 12498 3148
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 36096 3176 36124 3284
rect 36170 3272 36176 3324
rect 36228 3312 36234 3324
rect 37182 3312 37188 3324
rect 36228 3284 37188 3312
rect 36228 3272 36234 3284
rect 37182 3272 37188 3284
rect 37240 3272 37246 3324
rect 43346 3272 43352 3324
rect 43404 3312 43410 3324
rect 44082 3312 44088 3324
rect 43404 3284 44088 3312
rect 43404 3272 43410 3284
rect 44082 3272 44088 3284
rect 44140 3272 44146 3324
rect 44542 3272 44548 3324
rect 44600 3312 44606 3324
rect 45462 3312 45468 3324
rect 44600 3284 45468 3312
rect 44600 3272 44606 3284
rect 45462 3272 45468 3284
rect 45520 3272 45526 3324
rect 45738 3272 45744 3324
rect 45796 3312 45802 3324
rect 46842 3312 46848 3324
rect 45796 3284 46848 3312
rect 45796 3272 45802 3284
rect 46842 3272 46848 3284
rect 46900 3272 46906 3324
rect 50522 3272 50528 3324
rect 50580 3312 50586 3324
rect 50982 3312 50988 3324
rect 50580 3284 50988 3312
rect 50580 3272 50586 3284
rect 50982 3272 50988 3284
rect 51040 3272 51046 3324
rect 52822 3272 52828 3324
rect 52880 3312 52886 3324
rect 53742 3312 53748 3324
rect 52880 3284 53748 3312
rect 52880 3272 52886 3284
rect 53742 3272 53748 3284
rect 53800 3272 53806 3324
rect 65521 3315 65579 3321
rect 65521 3312 65533 3315
rect 53852 3284 65533 3312
rect 42150 3204 42156 3256
rect 42208 3244 42214 3256
rect 53852 3244 53880 3284
rect 65521 3281 65533 3284
rect 65567 3281 65579 3315
rect 65628 3312 65656 3352
rect 65705 3349 65717 3383
rect 65751 3380 65763 3383
rect 70581 3383 70639 3389
rect 70581 3380 70593 3383
rect 65751 3352 70593 3380
rect 65751 3349 65763 3352
rect 65705 3343 65763 3349
rect 70581 3349 70593 3352
rect 70627 3349 70639 3383
rect 70581 3343 70639 3349
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 79413 3383 79471 3389
rect 79413 3380 79425 3383
rect 70728 3352 79425 3380
rect 70728 3340 70734 3352
rect 79413 3349 79425 3352
rect 79459 3349 79471 3383
rect 79413 3343 79471 3349
rect 81253 3383 81311 3389
rect 81253 3349 81265 3383
rect 81299 3380 81311 3383
rect 86218 3380 86224 3392
rect 81299 3352 86224 3380
rect 81299 3349 81311 3352
rect 81253 3343 81311 3349
rect 86218 3340 86224 3352
rect 86276 3340 86282 3392
rect 104250 3340 104256 3392
rect 104308 3380 104314 3392
rect 112346 3380 112352 3392
rect 104308 3352 112352 3380
rect 104308 3340 104314 3352
rect 112346 3340 112352 3352
rect 112404 3340 112410 3392
rect 69201 3315 69259 3321
rect 69201 3312 69213 3315
rect 65628 3284 69213 3312
rect 65521 3275 65579 3281
rect 69201 3281 69213 3284
rect 69247 3281 69259 3315
rect 69201 3275 69259 3281
rect 69474 3272 69480 3324
rect 69532 3312 69538 3324
rect 86034 3312 86040 3324
rect 69532 3284 86040 3312
rect 69532 3272 69538 3284
rect 86034 3272 86040 3284
rect 86092 3272 86098 3324
rect 105998 3272 106004 3324
rect 106056 3312 106062 3324
rect 112441 3315 112499 3321
rect 112441 3312 112453 3315
rect 106056 3284 112453 3312
rect 106056 3272 106062 3284
rect 112441 3281 112453 3284
rect 112487 3281 112499 3315
rect 112548 3312 112576 3420
rect 112990 3408 112996 3460
rect 113048 3448 113054 3460
rect 133141 3451 133199 3457
rect 133141 3448 133153 3451
rect 113048 3420 133153 3448
rect 113048 3408 113054 3420
rect 133141 3417 133153 3420
rect 133187 3417 133199 3451
rect 133141 3411 133199 3417
rect 133690 3408 133696 3460
rect 133748 3448 133754 3460
rect 141881 3451 141939 3457
rect 141881 3448 141893 3451
rect 133748 3420 141893 3448
rect 133748 3408 133754 3420
rect 141881 3417 141893 3420
rect 141927 3417 141939 3451
rect 141881 3411 141939 3417
rect 141973 3451 142031 3457
rect 141973 3417 141985 3451
rect 142019 3448 142031 3451
rect 207474 3448 207480 3460
rect 142019 3420 207480 3448
rect 142019 3417 142031 3420
rect 141973 3411 142031 3417
rect 207474 3408 207480 3420
rect 207532 3408 207538 3460
rect 222102 3408 222108 3460
rect 222160 3448 222166 3460
rect 428734 3448 428740 3460
rect 222160 3420 428740 3448
rect 222160 3408 222166 3420
rect 428734 3408 428740 3420
rect 428792 3408 428798 3460
rect 494054 3408 494060 3460
rect 494112 3448 494118 3460
rect 495342 3448 495348 3460
rect 494112 3420 495348 3448
rect 494112 3408 494118 3420
rect 495342 3408 495348 3420
rect 495400 3408 495406 3460
rect 529382 3408 529388 3460
rect 529440 3448 529446 3460
rect 571426 3448 571432 3460
rect 529440 3420 571432 3448
rect 529440 3408 529446 3420
rect 571426 3408 571432 3420
rect 571484 3408 571490 3460
rect 112625 3383 112683 3389
rect 112625 3349 112637 3383
rect 112671 3380 112683 3383
rect 119430 3380 119436 3392
rect 112671 3352 119436 3380
rect 112671 3349 112683 3352
rect 112625 3343 112683 3349
rect 119430 3340 119436 3352
rect 119488 3340 119494 3392
rect 120721 3383 120779 3389
rect 120721 3349 120733 3383
rect 120767 3380 120779 3383
rect 127802 3380 127808 3392
rect 120767 3352 127808 3380
rect 120767 3349 120779 3352
rect 120721 3343 120779 3349
rect 127802 3340 127808 3352
rect 127860 3340 127866 3392
rect 127897 3383 127955 3389
rect 127897 3349 127909 3383
rect 127943 3380 127955 3383
rect 148229 3383 148287 3389
rect 127943 3352 148180 3380
rect 127943 3349 127955 3352
rect 127897 3343 127955 3349
rect 115934 3312 115940 3324
rect 112548 3284 115940 3312
rect 112441 3275 112499 3281
rect 115934 3272 115940 3284
rect 115992 3272 115998 3324
rect 116946 3272 116952 3324
rect 117004 3312 117010 3324
rect 142801 3315 142859 3321
rect 142801 3312 142813 3315
rect 117004 3284 142813 3312
rect 117004 3272 117010 3284
rect 142801 3281 142813 3284
rect 142847 3281 142859 3315
rect 142801 3275 142859 3281
rect 145834 3272 145840 3324
rect 145892 3312 145898 3324
rect 148042 3312 148048 3324
rect 145892 3284 148048 3312
rect 145892 3272 145898 3284
rect 148042 3272 148048 3284
rect 148100 3272 148106 3324
rect 148152 3312 148180 3352
rect 148229 3349 148241 3383
rect 148275 3380 148287 3383
rect 162121 3383 162179 3389
rect 162121 3380 162133 3383
rect 148275 3352 162133 3380
rect 148275 3349 148287 3352
rect 148229 3343 148287 3349
rect 162121 3349 162133 3352
rect 162167 3349 162179 3383
rect 162121 3343 162179 3349
rect 162213 3383 162271 3389
rect 162213 3349 162225 3383
rect 162259 3380 162271 3383
rect 165985 3383 166043 3389
rect 165985 3380 165997 3383
rect 162259 3352 165997 3380
rect 162259 3349 162271 3352
rect 162213 3343 162271 3349
rect 165985 3349 165997 3352
rect 166031 3349 166043 3383
rect 165985 3343 166043 3349
rect 166350 3340 166356 3392
rect 166408 3380 166414 3392
rect 178954 3380 178960 3392
rect 166408 3352 178960 3380
rect 166408 3340 166414 3352
rect 178954 3340 178960 3352
rect 179012 3340 179018 3392
rect 180058 3340 180064 3392
rect 180116 3380 180122 3392
rect 182637 3383 182695 3389
rect 182637 3380 182649 3383
rect 180116 3352 182649 3380
rect 180116 3340 180122 3352
rect 182637 3349 182649 3352
rect 182683 3349 182695 3383
rect 182637 3343 182695 3349
rect 182818 3340 182824 3392
rect 182876 3380 182882 3392
rect 186130 3380 186136 3392
rect 182876 3352 186136 3380
rect 182876 3340 182882 3352
rect 186130 3340 186136 3352
rect 186188 3340 186194 3392
rect 186225 3383 186283 3389
rect 186225 3349 186237 3383
rect 186271 3380 186283 3383
rect 271690 3380 271696 3392
rect 186271 3352 271696 3380
rect 186271 3349 186283 3352
rect 186225 3343 186283 3349
rect 271690 3340 271696 3352
rect 271748 3340 271754 3392
rect 275278 3340 275284 3392
rect 275336 3380 275342 3392
rect 277949 3383 278007 3389
rect 277949 3380 277961 3383
rect 275336 3352 277961 3380
rect 275336 3340 275342 3352
rect 277949 3349 277961 3352
rect 277995 3349 278007 3383
rect 277949 3343 278007 3349
rect 278041 3383 278099 3389
rect 278041 3349 278053 3383
rect 278087 3380 278099 3383
rect 382366 3380 382372 3392
rect 278087 3352 382372 3380
rect 278087 3349 278099 3352
rect 278041 3343 278099 3349
rect 382366 3340 382372 3352
rect 382424 3340 382430 3392
rect 390646 3340 390652 3392
rect 390704 3380 390710 3392
rect 391842 3380 391848 3392
rect 390704 3352 391848 3380
rect 390704 3340 390710 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 156322 3312 156328 3324
rect 148152 3284 156328 3312
rect 156322 3272 156328 3284
rect 156380 3272 156386 3324
rect 186314 3312 186320 3324
rect 156432 3284 186320 3312
rect 70489 3247 70547 3253
rect 70489 3244 70501 3247
rect 42208 3216 53880 3244
rect 53944 3216 70501 3244
rect 42208 3204 42214 3216
rect 40681 3179 40739 3185
rect 40681 3176 40693 3179
rect 36096 3148 40693 3176
rect 40681 3145 40693 3148
rect 40727 3145 40739 3179
rect 40681 3139 40739 3145
rect 48130 3136 48136 3188
rect 48188 3176 48194 3188
rect 53944 3176 53972 3216
rect 70489 3213 70501 3216
rect 70535 3213 70547 3247
rect 70489 3207 70547 3213
rect 70581 3247 70639 3253
rect 70581 3213 70593 3247
rect 70627 3244 70639 3247
rect 74902 3244 74908 3256
rect 70627 3216 74908 3244
rect 70627 3213 70639 3216
rect 70581 3207 70639 3213
rect 74902 3204 74908 3216
rect 74960 3204 74966 3256
rect 74997 3247 75055 3253
rect 74997 3213 75009 3247
rect 75043 3244 75055 3247
rect 77478 3244 77484 3256
rect 75043 3216 77484 3244
rect 75043 3213 75055 3216
rect 74997 3207 75055 3213
rect 77478 3204 77484 3216
rect 77536 3204 77542 3256
rect 77846 3204 77852 3256
rect 77904 3244 77910 3256
rect 88426 3244 88432 3256
rect 77904 3216 88432 3244
rect 77904 3204 77910 3216
rect 88426 3204 88432 3216
rect 88484 3204 88490 3256
rect 103422 3204 103428 3256
rect 103480 3244 103486 3256
rect 114738 3244 114744 3256
rect 103480 3216 114744 3244
rect 103480 3204 103486 3216
rect 114738 3204 114744 3216
rect 114796 3204 114802 3256
rect 115842 3204 115848 3256
rect 115900 3244 115906 3256
rect 145650 3244 145656 3256
rect 115900 3216 145656 3244
rect 115900 3204 115906 3216
rect 145650 3204 145656 3216
rect 145708 3204 145714 3256
rect 147677 3247 147735 3253
rect 147677 3213 147689 3247
rect 147723 3244 147735 3247
rect 152461 3247 152519 3253
rect 152461 3244 152473 3247
rect 147723 3216 152473 3244
rect 147723 3213 147735 3216
rect 147677 3207 147735 3213
rect 152461 3213 152473 3216
rect 152507 3213 152519 3247
rect 152461 3207 152519 3213
rect 152550 3204 152556 3256
rect 152608 3244 152614 3256
rect 156432 3244 156460 3284
rect 186314 3272 186320 3284
rect 186372 3272 186378 3324
rect 186406 3272 186412 3324
rect 186464 3312 186470 3324
rect 282454 3312 282460 3324
rect 186464 3284 282460 3312
rect 186464 3272 186470 3284
rect 282454 3272 282460 3284
rect 282512 3272 282518 3324
rect 282549 3315 282607 3321
rect 282549 3281 282561 3315
rect 282595 3312 282607 3315
rect 293126 3312 293132 3324
rect 282595 3284 293132 3312
rect 282595 3281 282607 3284
rect 282549 3275 282607 3281
rect 293126 3272 293132 3284
rect 293184 3272 293190 3324
rect 293218 3272 293224 3324
rect 293276 3312 293282 3324
rect 400214 3312 400220 3324
rect 293276 3284 400220 3312
rect 293276 3272 293282 3284
rect 400214 3272 400220 3284
rect 400272 3272 400278 3324
rect 152608 3216 156460 3244
rect 156509 3247 156567 3253
rect 152608 3204 152614 3216
rect 156509 3213 156521 3247
rect 156555 3244 156567 3247
rect 176654 3244 176660 3256
rect 156555 3216 176660 3244
rect 156555 3213 156567 3216
rect 156509 3207 156567 3213
rect 176654 3204 176660 3216
rect 176712 3204 176718 3256
rect 181349 3247 181407 3253
rect 181349 3213 181361 3247
rect 181395 3244 181407 3247
rect 186038 3244 186044 3256
rect 181395 3216 186044 3244
rect 181395 3213 181407 3216
rect 181349 3207 181407 3213
rect 186038 3204 186044 3216
rect 186096 3204 186102 3256
rect 186133 3247 186191 3253
rect 186133 3213 186145 3247
rect 186179 3244 186191 3247
rect 253842 3244 253848 3256
rect 186179 3216 253848 3244
rect 186179 3213 186191 3216
rect 186133 3207 186191 3213
rect 253842 3204 253848 3216
rect 253900 3204 253906 3256
rect 255958 3204 255964 3256
rect 256016 3244 256022 3256
rect 339494 3244 339500 3256
rect 256016 3216 339500 3244
rect 256016 3204 256022 3216
rect 339494 3204 339500 3216
rect 339552 3204 339558 3256
rect 347774 3204 347780 3256
rect 347832 3244 347838 3256
rect 349062 3244 349068 3256
rect 347832 3216 349068 3244
rect 347832 3204 347838 3216
rect 349062 3204 349068 3216
rect 349120 3204 349126 3256
rect 48188 3148 53972 3176
rect 54113 3179 54171 3185
rect 48188 3136 48194 3148
rect 54113 3145 54125 3179
rect 54159 3176 54171 3179
rect 77294 3176 77300 3188
rect 54159 3148 77300 3176
rect 54159 3145 54171 3148
rect 54113 3139 54171 3145
rect 77294 3136 77300 3148
rect 77352 3136 77358 3188
rect 103330 3136 103336 3188
rect 103388 3176 103394 3188
rect 113542 3176 113548 3188
rect 103388 3148 113548 3176
rect 103388 3136 103394 3148
rect 113542 3136 113548 3148
rect 113600 3136 113606 3188
rect 114278 3136 114284 3188
rect 114336 3176 114342 3188
rect 143258 3176 143264 3188
rect 114336 3148 143264 3176
rect 114336 3136 114342 3148
rect 143258 3136 143264 3148
rect 143316 3136 143322 3188
rect 143445 3179 143503 3185
rect 143445 3145 143457 3179
rect 143491 3176 143503 3179
rect 152734 3176 152740 3188
rect 143491 3148 152740 3176
rect 143491 3145 143503 3148
rect 143445 3139 143503 3145
rect 152734 3136 152740 3148
rect 152792 3136 152798 3188
rect 152829 3179 152887 3185
rect 152829 3145 152841 3179
rect 152875 3176 152887 3179
rect 157518 3176 157524 3188
rect 152875 3148 157524 3176
rect 152875 3145 152887 3148
rect 152829 3139 152887 3145
rect 157518 3136 157524 3148
rect 157576 3136 157582 3188
rect 157981 3179 158039 3185
rect 157981 3145 157993 3179
rect 158027 3176 158039 3179
rect 173161 3179 173219 3185
rect 173161 3176 173173 3179
rect 158027 3148 173173 3176
rect 158027 3145 158039 3148
rect 157981 3139 158039 3145
rect 173161 3145 173173 3148
rect 173207 3145 173219 3179
rect 173161 3139 173219 3145
rect 181441 3179 181499 3185
rect 181441 3145 181453 3179
rect 181487 3176 181499 3179
rect 246758 3176 246764 3188
rect 181487 3148 246764 3176
rect 181487 3145 181499 3148
rect 181441 3139 181499 3145
rect 246758 3136 246764 3148
rect 246816 3136 246822 3188
rect 253198 3136 253204 3188
rect 253256 3176 253262 3188
rect 328822 3176 328828 3188
rect 253256 3148 328828 3176
rect 253256 3136 253262 3148
rect 328822 3136 328828 3148
rect 328880 3136 328886 3188
rect 8846 3068 8852 3120
rect 8904 3108 8910 3120
rect 9582 3108 9588 3120
rect 8904 3080 9588 3108
rect 8904 3068 8910 3080
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 35897 3111 35955 3117
rect 35897 3077 35909 3111
rect 35943 3108 35955 3111
rect 45465 3111 45523 3117
rect 45465 3108 45477 3111
rect 35943 3080 45477 3108
rect 35943 3077 35955 3080
rect 35897 3071 35955 3077
rect 45465 3077 45477 3080
rect 45511 3077 45523 3111
rect 45465 3071 45523 3077
rect 49326 3068 49332 3120
rect 49384 3108 49390 3120
rect 74905 3111 74963 3117
rect 74905 3108 74917 3111
rect 49384 3080 74917 3108
rect 49384 3068 49390 3080
rect 74905 3077 74917 3080
rect 74951 3077 74963 3111
rect 74905 3071 74963 3077
rect 74997 3111 75055 3117
rect 74997 3077 75009 3111
rect 75043 3108 75055 3111
rect 79505 3111 79563 3117
rect 79505 3108 79517 3111
rect 75043 3080 79517 3108
rect 75043 3077 75055 3080
rect 74997 3071 75055 3077
rect 79505 3077 79517 3080
rect 79551 3077 79563 3111
rect 79505 3071 79563 3077
rect 104158 3068 104164 3120
rect 104216 3108 104222 3120
rect 107562 3108 107568 3120
rect 104216 3080 107568 3108
rect 104216 3068 104222 3080
rect 107562 3068 107568 3080
rect 107620 3068 107626 3120
rect 110322 3068 110328 3120
rect 110380 3108 110386 3120
rect 130194 3108 130200 3120
rect 110380 3080 130200 3108
rect 110380 3068 110386 3080
rect 130194 3068 130200 3080
rect 130252 3068 130258 3120
rect 133141 3111 133199 3117
rect 133141 3077 133153 3111
rect 133187 3108 133199 3111
rect 138474 3108 138480 3120
rect 133187 3080 138480 3108
rect 133187 3077 133199 3080
rect 133141 3071 133199 3077
rect 138474 3068 138480 3080
rect 138532 3068 138538 3120
rect 141789 3111 141847 3117
rect 141789 3077 141801 3111
rect 141835 3108 141847 3111
rect 147677 3111 147735 3117
rect 147677 3108 147689 3111
rect 141835 3080 147689 3108
rect 141835 3077 141847 3080
rect 141789 3071 141847 3077
rect 147677 3077 147689 3080
rect 147723 3077 147735 3111
rect 147677 3071 147735 3077
rect 160738 3068 160744 3120
rect 160796 3108 160802 3120
rect 162029 3111 162087 3117
rect 162029 3108 162041 3111
rect 160796 3080 162041 3108
rect 160796 3068 160802 3080
rect 162029 3077 162041 3080
rect 162075 3077 162087 3111
rect 162029 3071 162087 3077
rect 164878 3068 164884 3120
rect 164936 3108 164942 3120
rect 175366 3108 175372 3120
rect 164936 3080 175372 3108
rect 164936 3068 164942 3080
rect 175366 3068 175372 3080
rect 175424 3068 175430 3120
rect 235994 3108 236000 3120
rect 176764 3080 236000 3108
rect 51626 3000 51632 3052
rect 51684 3040 51690 3052
rect 70397 3043 70455 3049
rect 70397 3040 70409 3043
rect 51684 3012 70409 3040
rect 51684 3000 51690 3012
rect 70397 3009 70409 3012
rect 70443 3009 70455 3043
rect 70397 3003 70455 3009
rect 70489 3043 70547 3049
rect 70489 3009 70501 3043
rect 70535 3040 70547 3043
rect 77386 3040 77392 3052
rect 70535 3012 77392 3040
rect 70535 3009 70547 3012
rect 70489 3003 70547 3009
rect 77386 3000 77392 3012
rect 77444 3000 77450 3052
rect 86126 3000 86132 3052
rect 86184 3040 86190 3052
rect 92658 3040 92664 3052
rect 86184 3012 92664 3040
rect 86184 3000 86190 3012
rect 92658 3000 92664 3012
rect 92716 3000 92722 3052
rect 114370 3000 114376 3052
rect 114428 3040 114434 3052
rect 142062 3040 142068 3052
rect 114428 3012 142068 3040
rect 114428 3000 114434 3012
rect 142062 3000 142068 3012
rect 142120 3000 142126 3052
rect 142801 3043 142859 3049
rect 142801 3009 142813 3043
rect 142847 3040 142859 3043
rect 149238 3040 149244 3052
rect 142847 3012 149244 3040
rect 142847 3009 142859 3012
rect 142801 3003 142859 3009
rect 149238 3000 149244 3012
rect 149296 3000 149302 3052
rect 160465 3043 160523 3049
rect 160465 3040 160477 3043
rect 152476 3012 160477 3040
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 22002 2972 22008 2984
rect 20772 2944 22008 2972
rect 20772 2932 20778 2944
rect 22002 2932 22008 2944
rect 22060 2932 22066 2984
rect 54018 2932 54024 2984
rect 54076 2972 54082 2984
rect 80054 2972 80060 2984
rect 54076 2944 80060 2972
rect 54076 2932 54082 2944
rect 80054 2932 80060 2944
rect 80112 2932 80118 2984
rect 113082 2932 113088 2984
rect 113140 2972 113146 2984
rect 139670 2972 139676 2984
rect 113140 2944 139676 2972
rect 113140 2932 113146 2944
rect 139670 2932 139676 2944
rect 139728 2932 139734 2984
rect 46934 2864 46940 2916
rect 46992 2904 46998 2916
rect 54113 2907 54171 2913
rect 54113 2904 54125 2907
rect 46992 2876 54125 2904
rect 46992 2864 46998 2876
rect 54113 2873 54125 2876
rect 54159 2873 54171 2907
rect 54113 2867 54171 2873
rect 56410 2864 56416 2916
rect 56468 2904 56474 2916
rect 80146 2904 80152 2916
rect 56468 2876 80152 2904
rect 56468 2864 56474 2876
rect 80146 2864 80152 2876
rect 80204 2864 80210 2916
rect 111610 2864 111616 2916
rect 111668 2904 111674 2916
rect 134886 2904 134892 2916
rect 111668 2876 134892 2904
rect 111668 2864 111674 2876
rect 134886 2864 134892 2876
rect 134944 2864 134950 2916
rect 139302 2864 139308 2916
rect 139360 2904 139366 2916
rect 141973 2907 142031 2913
rect 141973 2904 141985 2907
rect 139360 2876 141985 2904
rect 139360 2864 139366 2876
rect 141973 2873 141985 2876
rect 142019 2873 142031 2907
rect 141973 2867 142031 2873
rect 145558 2864 145564 2916
rect 145616 2904 145622 2916
rect 152476 2904 152504 3012
rect 160465 3009 160477 3012
rect 160511 3009 160523 3043
rect 160465 3003 160523 3009
rect 160649 3043 160707 3049
rect 160649 3009 160661 3043
rect 160695 3040 160707 3043
rect 176562 3040 176568 3052
rect 160695 3012 176568 3040
rect 160695 3009 160707 3012
rect 160649 3003 160707 3009
rect 176562 3000 176568 3012
rect 176620 3000 176626 3052
rect 176764 3040 176792 3080
rect 235994 3068 236000 3080
rect 236052 3068 236058 3120
rect 271230 3068 271236 3120
rect 271288 3108 271294 3120
rect 278041 3111 278099 3117
rect 278041 3108 278053 3111
rect 271288 3080 278053 3108
rect 271288 3068 271294 3080
rect 278041 3077 278053 3080
rect 278087 3077 278099 3111
rect 278041 3071 278099 3077
rect 278133 3111 278191 3117
rect 278133 3077 278145 3111
rect 278179 3108 278191 3111
rect 282549 3111 282607 3117
rect 282549 3108 282561 3111
rect 278179 3080 282561 3108
rect 278179 3077 278191 3080
rect 278133 3071 278191 3077
rect 282549 3077 282561 3080
rect 282595 3077 282607 3111
rect 282549 3071 282607 3077
rect 291838 3068 291844 3120
rect 291896 3108 291902 3120
rect 368014 3108 368020 3120
rect 291896 3080 368020 3108
rect 291896 3068 291902 3080
rect 368014 3068 368020 3080
rect 368072 3068 368078 3120
rect 176672 3012 176792 3040
rect 176841 3043 176899 3049
rect 157981 2975 158039 2981
rect 157981 2972 157993 2975
rect 145616 2876 152504 2904
rect 152568 2944 157993 2972
rect 145616 2864 145622 2876
rect 58802 2796 58808 2848
rect 58860 2836 58866 2848
rect 74997 2839 75055 2845
rect 74997 2836 75009 2839
rect 58860 2808 75009 2836
rect 58860 2796 58866 2808
rect 74997 2805 75009 2808
rect 75043 2805 75055 2839
rect 74997 2799 75055 2805
rect 75089 2839 75147 2845
rect 75089 2805 75101 2839
rect 75135 2836 75147 2839
rect 83090 2836 83096 2848
rect 75135 2808 83096 2836
rect 75135 2805 75147 2808
rect 75089 2799 75147 2805
rect 83090 2796 83096 2808
rect 83148 2796 83154 2848
rect 95418 2796 95424 2848
rect 95476 2836 95482 2848
rect 95694 2836 95700 2848
rect 95476 2808 95700 2836
rect 95476 2796 95482 2808
rect 95694 2796 95700 2808
rect 95752 2796 95758 2848
rect 108850 2796 108856 2848
rect 108908 2836 108914 2848
rect 126606 2836 126612 2848
rect 108908 2808 126612 2836
rect 108908 2796 108914 2808
rect 126606 2796 126612 2808
rect 126664 2796 126670 2848
rect 126701 2839 126759 2845
rect 126701 2805 126713 2839
rect 126747 2836 126759 2839
rect 129550 2836 129556 2848
rect 126747 2808 129556 2836
rect 126747 2805 126759 2808
rect 126701 2799 126759 2805
rect 129550 2796 129556 2808
rect 129608 2796 129614 2848
rect 129642 2796 129648 2848
rect 129700 2836 129706 2848
rect 133877 2839 133935 2845
rect 133877 2836 133889 2839
rect 129700 2808 133889 2836
rect 129700 2796 129706 2808
rect 133877 2805 133889 2808
rect 133923 2805 133935 2839
rect 133877 2799 133935 2805
rect 133966 2796 133972 2848
rect 134024 2836 134030 2848
rect 137557 2839 137615 2845
rect 137557 2836 137569 2839
rect 134024 2808 137569 2836
rect 134024 2796 134030 2808
rect 137557 2805 137569 2808
rect 137603 2805 137615 2839
rect 137557 2799 137615 2805
rect 148410 2796 148416 2848
rect 148468 2836 148474 2848
rect 152568 2836 152596 2944
rect 157981 2941 157993 2944
rect 158027 2941 158039 2975
rect 157981 2935 158039 2941
rect 162213 2975 162271 2981
rect 162213 2941 162225 2975
rect 162259 2972 162271 2975
rect 171778 2972 171784 2984
rect 162259 2944 171784 2972
rect 162259 2941 162271 2944
rect 162213 2935 162271 2941
rect 171778 2932 171784 2944
rect 171836 2932 171842 2984
rect 173158 2932 173164 2984
rect 173216 2972 173222 2984
rect 176672 2972 176700 3012
rect 176841 3009 176853 3043
rect 176887 3040 176899 3043
rect 181349 3043 181407 3049
rect 181349 3040 181361 3043
rect 176887 3012 181361 3040
rect 176887 3009 176899 3012
rect 176841 3003 176899 3009
rect 181349 3009 181361 3012
rect 181395 3009 181407 3043
rect 181349 3003 181407 3009
rect 181533 3043 181591 3049
rect 181533 3009 181545 3043
rect 181579 3040 181591 3043
rect 239582 3040 239588 3052
rect 181579 3012 239588 3040
rect 181579 3009 181591 3012
rect 181533 3003 181591 3009
rect 239582 3000 239588 3012
rect 239640 3000 239646 3052
rect 250438 3000 250444 3052
rect 250496 3040 250502 3052
rect 325234 3040 325240 3052
rect 250496 3012 325240 3040
rect 250496 3000 250502 3012
rect 325234 3000 325240 3012
rect 325292 3000 325298 3052
rect 173216 2944 176700 2972
rect 173216 2932 173222 2944
rect 176746 2932 176752 2984
rect 176804 2972 176810 2984
rect 225322 2972 225328 2984
rect 176804 2944 225328 2972
rect 176804 2932 176810 2944
rect 225322 2932 225328 2944
rect 225380 2932 225386 2984
rect 253290 2932 253296 2984
rect 253348 2972 253354 2984
rect 278866 2972 278872 2984
rect 253348 2944 278872 2972
rect 253348 2932 253354 2944
rect 278866 2932 278872 2944
rect 278924 2932 278930 2984
rect 289078 2932 289084 2984
rect 289136 2972 289142 2984
rect 353754 2972 353760 2984
rect 289136 2944 353760 2972
rect 289136 2932 289142 2944
rect 353754 2932 353760 2944
rect 353812 2932 353818 2984
rect 159361 2907 159419 2913
rect 159361 2873 159373 2907
rect 159407 2904 159419 2907
rect 165890 2904 165896 2916
rect 159407 2876 165896 2904
rect 159407 2873 159419 2876
rect 159361 2867 159419 2873
rect 165890 2864 165896 2876
rect 165948 2864 165954 2916
rect 165985 2907 166043 2913
rect 165985 2873 165997 2907
rect 166031 2904 166043 2907
rect 202690 2904 202696 2916
rect 166031 2876 202696 2904
rect 166031 2873 166043 2876
rect 165985 2867 166043 2873
rect 202690 2864 202696 2876
rect 202748 2864 202754 2916
rect 246298 2864 246304 2916
rect 246356 2904 246362 2916
rect 275278 2904 275284 2916
rect 246356 2876 275284 2904
rect 246356 2864 246362 2876
rect 275278 2864 275284 2876
rect 275336 2864 275342 2916
rect 285950 2904 285956 2916
rect 277504 2876 285956 2904
rect 148468 2808 152596 2836
rect 148468 2796 148474 2808
rect 156598 2796 156604 2848
rect 156656 2836 156662 2848
rect 197998 2836 198004 2848
rect 156656 2808 198004 2836
rect 156656 2796 156662 2808
rect 197998 2796 198004 2808
rect 198056 2796 198062 2848
rect 271138 2796 271144 2848
rect 271196 2836 271202 2848
rect 277504 2836 277532 2876
rect 285950 2864 285956 2876
rect 286008 2864 286014 2916
rect 286318 2864 286324 2916
rect 286376 2904 286382 2916
rect 303798 2904 303804 2916
rect 286376 2876 303804 2904
rect 286376 2864 286382 2876
rect 303798 2864 303804 2876
rect 303856 2864 303862 2916
rect 304994 2864 305000 2916
rect 305052 2904 305058 2916
rect 306190 2904 306196 2916
rect 305052 2876 306196 2904
rect 305052 2864 305058 2876
rect 306190 2864 306196 2876
rect 306248 2864 306254 2916
rect 271196 2808 277532 2836
rect 271196 2796 271202 2808
rect 279418 2796 279424 2848
rect 279476 2836 279482 2848
rect 296714 2836 296720 2848
rect 279476 2808 296720 2836
rect 279476 2796 279482 2808
rect 296714 2796 296720 2808
rect 296772 2796 296778 2848
rect 173161 2771 173219 2777
rect 173161 2737 173173 2771
rect 173207 2768 173219 2771
rect 180150 2768 180156 2780
rect 173207 2740 180156 2768
rect 173207 2737 173219 2740
rect 173161 2731 173219 2737
rect 180150 2728 180156 2740
rect 180208 2728 180214 2780
rect 273438 2320 273444 2372
rect 273496 2360 273502 2372
rect 280062 2360 280068 2372
rect 273496 2332 280068 2360
rect 273496 2320 273502 2332
rect 280062 2320 280068 2332
rect 280120 2320 280126 2372
rect 365714 1368 365720 1420
rect 365772 1408 365778 1420
rect 366910 1408 366916 1420
rect 365772 1380 366916 1408
rect 365772 1368 365778 1380
rect 366910 1368 366916 1380
rect 366968 1368 366974 1420
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 5442 592 5448 604
rect 5316 564 5448 592
rect 5316 552 5322 564
rect 5442 552 5448 564
rect 5500 552 5506 604
rect 23106 552 23112 604
rect 23164 592 23170 604
rect 23382 592 23388 604
rect 23164 564 23388 592
rect 23164 552 23170 564
rect 23382 552 23388 564
rect 23440 552 23446 604
rect 92106 552 92112 604
rect 92164 592 92170 604
rect 92382 592 92388 604
rect 92164 564 92388 592
rect 92164 552 92170 564
rect 92382 552 92388 564
rect 92440 552 92446 604
rect 95418 552 95424 604
rect 95476 592 95482 604
rect 95694 592 95700 604
rect 95476 564 95700 592
rect 95476 552 95482 564
rect 95694 552 95700 564
rect 95752 552 95758 604
rect 128630 552 128636 604
rect 128688 592 128694 604
rect 128998 592 129004 604
rect 128688 564 129004 592
rect 128688 552 128694 564
rect 128998 552 129004 564
rect 129056 552 129062 604
rect 140866 592 140872 604
rect 140827 564 140872 592
rect 140866 552 140872 564
rect 140924 552 140930 604
rect 295334 552 295340 604
rect 295392 592 295398 604
rect 295518 592 295524 604
rect 295392 564 295524 592
rect 295392 552 295398 564
rect 295518 552 295524 564
rect 295576 552 295582 604
rect 298094 552 298100 604
rect 298152 592 298158 604
rect 299106 592 299112 604
rect 298152 564 299112 592
rect 298152 552 298158 564
rect 299106 552 299112 564
rect 299164 552 299170 604
rect 309134 552 309140 604
rect 309192 592 309198 604
rect 309778 592 309784 604
rect 309192 564 309784 592
rect 309192 552 309198 564
rect 309778 552 309784 564
rect 309836 552 309842 604
rect 316034 552 316040 604
rect 316092 592 316098 604
rect 316954 592 316960 604
rect 316092 564 316960 592
rect 316092 552 316098 564
rect 316954 552 316960 564
rect 317012 552 317018 604
rect 317414 552 317420 604
rect 317472 592 317478 604
rect 318058 592 318064 604
rect 317472 564 318064 592
rect 317472 552 317478 564
rect 318058 552 318064 564
rect 318116 552 318122 604
rect 322934 552 322940 604
rect 322992 592 322998 604
rect 324038 592 324044 604
rect 322992 564 324044 592
rect 322992 552 322998 564
rect 324038 552 324044 564
rect 324096 552 324102 604
rect 327074 552 327080 604
rect 327132 592 327138 604
rect 327626 592 327632 604
rect 327132 564 327632 592
rect 327132 552 327138 564
rect 327626 552 327632 564
rect 327684 552 327690 604
rect 333974 552 333980 604
rect 334032 592 334038 604
rect 334710 592 334716 604
rect 334032 564 334716 592
rect 334032 552 334038 564
rect 334710 552 334716 564
rect 334768 552 334774 604
rect 340874 552 340880 604
rect 340932 592 340938 604
rect 341886 592 341892 604
rect 340932 564 341892 592
rect 340932 552 340938 564
rect 341886 552 341892 564
rect 341944 552 341950 604
rect 342254 552 342260 604
rect 342312 592 342318 604
rect 343082 592 343088 604
rect 342312 564 343088 592
rect 342312 552 342318 564
rect 343082 552 343088 564
rect 343140 552 343146 604
rect 364334 552 364340 604
rect 364392 592 364398 604
rect 364518 592 364524 604
rect 364392 564 364524 592
rect 364392 552 364398 564
rect 364518 552 364524 564
rect 364576 552 364582 604
rect 369854 552 369860 604
rect 369912 592 369918 604
rect 370406 592 370412 604
rect 369912 564 370412 592
rect 369912 552 369918 564
rect 370406 552 370412 564
rect 370464 552 370470 604
rect 376754 552 376760 604
rect 376812 592 376818 604
rect 377582 592 377588 604
rect 376812 564 377588 592
rect 376812 552 376818 564
rect 377582 552 377588 564
rect 377640 552 377646 604
rect 378134 552 378140 604
rect 378192 592 378198 604
rect 378778 592 378784 604
rect 378192 564 378784 592
rect 378192 552 378198 564
rect 378778 552 378784 564
rect 378836 552 378842 604
rect 412634 552 412640 604
rect 412692 592 412698 604
rect 413278 592 413284 604
rect 412692 564 413284 592
rect 412692 552 412698 564
rect 413278 552 413284 564
rect 413336 552 413342 604
rect 419534 552 419540 604
rect 419592 592 419598 604
rect 420362 592 420368 604
rect 419592 564 420368 592
rect 419592 552 419598 564
rect 420362 552 420368 564
rect 420420 552 420426 604
rect 420914 552 420920 604
rect 420972 592 420978 604
rect 421558 592 421564 604
rect 420972 564 421564 592
rect 420972 552 420978 564
rect 421558 552 421564 564
rect 421616 552 421622 604
rect 423674 552 423680 604
rect 423732 592 423738 604
rect 423950 592 423956 604
rect 423732 564 423956 592
rect 423732 552 423738 564
rect 423950 552 423956 564
rect 424008 552 424014 604
rect 426434 552 426440 604
rect 426492 592 426498 604
rect 427538 592 427544 604
rect 426492 564 427544 592
rect 426492 552 426498 564
rect 427538 552 427544 564
rect 427596 552 427602 604
rect 430574 552 430580 604
rect 430632 592 430638 604
rect 431126 592 431132 604
rect 430632 564 431132 592
rect 430632 552 430638 564
rect 431126 552 431132 564
rect 431184 552 431190 604
rect 438854 552 438860 604
rect 438912 592 438918 604
rect 439406 592 439412 604
rect 438912 564 439412 592
rect 438912 552 438918 564
rect 439406 552 439412 564
rect 439464 552 439470 604
rect 441614 552 441620 604
rect 441672 592 441678 604
rect 441798 592 441804 604
rect 441672 564 441804 592
rect 441672 552 441678 564
rect 441798 552 441804 564
rect 441856 552 441862 604
rect 444374 552 444380 604
rect 444432 592 444438 604
rect 445386 592 445392 604
rect 444432 564 445392 592
rect 444432 552 444438 564
rect 445386 552 445392 564
rect 445444 552 445450 604
rect 445754 552 445760 604
rect 445812 592 445818 604
rect 446582 592 446588 604
rect 445812 564 446588 592
rect 445812 552 445818 564
rect 446582 552 446588 564
rect 446640 552 446646 604
rect 448514 552 448520 604
rect 448572 592 448578 604
rect 448974 592 448980 604
rect 448572 564 448980 592
rect 448572 552 448578 564
rect 448974 552 448980 564
rect 449032 552 449038 604
rect 452654 552 452660 604
rect 452712 592 452718 604
rect 453666 592 453672 604
rect 452712 564 453672 592
rect 452712 552 452718 564
rect 453666 552 453672 564
rect 453724 552 453730 604
rect 455414 552 455420 604
rect 455472 592 455478 604
rect 456058 592 456064 604
rect 455472 564 456064 592
rect 455472 552 455478 564
rect 456058 552 456064 564
rect 456116 552 456122 604
rect 462314 552 462320 604
rect 462372 592 462378 604
rect 463234 592 463240 604
rect 462372 564 463240 592
rect 462372 552 462378 564
rect 463234 552 463240 564
rect 463292 552 463298 604
rect 466454 552 466460 604
rect 466512 592 466518 604
rect 466822 592 466828 604
rect 466512 564 466828 592
rect 466512 552 466518 564
rect 466822 552 466828 564
rect 466880 552 466886 604
rect 469214 552 469220 604
rect 469272 592 469278 604
rect 470318 592 470324 604
rect 469272 564 470324 592
rect 469272 552 469278 564
rect 470318 552 470324 564
rect 470376 552 470382 604
rect 489914 552 489920 604
rect 489972 592 489978 604
rect 490558 592 490564 604
rect 489972 564 490564 592
rect 489972 552 489978 564
rect 490558 552 490564 564
rect 490616 552 490622 604
rect 495434 552 495440 604
rect 495492 592 495498 604
rect 496538 592 496544 604
rect 495492 564 496544 592
rect 495492 552 495498 564
rect 496538 552 496544 564
rect 496596 552 496602 604
rect 496814 552 496820 604
rect 496872 592 496878 604
rect 497734 592 497740 604
rect 496872 564 497740 592
rect 496872 552 496878 564
rect 497734 552 497740 564
rect 497792 552 497798 604
rect 499574 552 499580 604
rect 499632 592 499638 604
rect 500126 592 500132 604
rect 499632 564 500132 592
rect 499632 552 499638 564
rect 500126 552 500132 564
rect 500184 552 500190 604
rect 500954 552 500960 604
rect 501012 592 501018 604
rect 501230 592 501236 604
rect 501012 564 501236 592
rect 501012 552 501018 564
rect 501230 552 501236 564
rect 501288 552 501294 604
rect 503714 552 503720 604
rect 503772 592 503778 604
rect 504818 592 504824 604
rect 503772 564 504824 592
rect 503772 552 503778 564
rect 504818 552 504824 564
rect 504876 552 504882 604
rect 506474 552 506480 604
rect 506532 592 506538 604
rect 507210 592 507216 604
rect 506532 564 507216 592
rect 506532 552 506538 564
rect 507210 552 507216 564
rect 507268 552 507274 604
rect 507854 552 507860 604
rect 507912 592 507918 604
rect 508406 592 508412 604
rect 507912 564 508412 592
rect 507912 552 507918 564
rect 508406 552 508412 564
rect 508464 552 508470 604
rect 510614 552 510620 604
rect 510672 592 510678 604
rect 510798 592 510804 604
rect 510672 564 510804 592
rect 510672 552 510678 564
rect 510798 552 510804 564
rect 510856 552 510862 604
rect 513374 552 513380 604
rect 513432 592 513438 604
rect 514386 592 514392 604
rect 513432 564 514392 592
rect 513432 552 513438 564
rect 514386 552 514392 564
rect 514444 552 514450 604
rect 524414 552 524420 604
rect 524472 592 524478 604
rect 525058 592 525064 604
rect 524472 564 525064 592
rect 524472 552 524478 564
rect 525058 552 525064 564
rect 525116 552 525122 604
rect 538214 552 538220 604
rect 538272 592 538278 604
rect 539318 592 539324 604
rect 538272 564 539324 592
rect 538272 552 538278 564
rect 539318 552 539324 564
rect 539376 552 539382 604
rect 542354 552 542360 604
rect 542412 592 542418 604
rect 542906 592 542912 604
rect 542412 564 542912 592
rect 542412 552 542418 564
rect 542906 552 542912 564
rect 542964 552 542970 604
rect 549254 552 549260 604
rect 549312 592 549318 604
rect 550082 592 550088 604
rect 549312 564 550088 592
rect 549312 552 549318 564
rect 550082 552 550088 564
rect 550140 552 550146 604
rect 556154 552 556160 604
rect 556212 592 556218 604
rect 557166 592 557172 604
rect 556212 564 557172 592
rect 556212 552 556218 564
rect 557166 552 557172 564
rect 557224 552 557230 604
<< via1 >>
rect 264888 653352 264940 653404
rect 378140 653352 378192 653404
rect 383568 653352 383620 653404
rect 508412 653352 508464 653404
rect 259184 652876 259236 652928
rect 263600 652876 263652 652928
rect 264888 652876 264940 652928
rect 378140 652876 378192 652928
rect 383568 652876 383620 652928
rect 508412 652808 508464 652860
rect 513380 652808 513432 652860
rect 129280 652740 129332 652792
rect 133696 652740 133748 652792
rect 139400 652740 139452 652792
rect 518900 652740 518952 652792
rect 137652 650428 137704 650480
rect 266452 650496 266504 650548
rect 282828 650428 282880 650480
rect 516416 650428 516468 650480
rect 266452 650224 266504 650276
rect 387156 650224 387208 650276
rect 282276 650156 282328 650208
rect 282828 650156 282880 650208
rect 294696 645872 294748 645924
rect 307392 645872 307444 645924
rect 291844 644444 291896 644496
rect 307116 644444 307168 644496
rect 290464 643084 290516 643136
rect 307116 643084 307168 643136
rect 287704 641724 287756 641776
rect 307668 641724 307720 641776
rect 286324 640296 286376 640348
rect 307668 640296 307720 640348
rect 284944 638936 284996 638988
rect 306656 638936 306708 638988
rect 294604 637576 294656 637628
rect 306840 637576 306892 637628
rect 389180 580252 389232 580304
rect 437848 580252 437900 580304
rect 302884 579640 302936 579692
rect 306932 579640 306984 579692
rect 139400 579572 139452 579624
rect 187700 579572 187752 579624
rect 282184 578892 282236 578944
rect 307668 578892 307720 578944
rect 66168 558832 66220 558884
rect 200212 558832 200264 558884
rect 282092 558832 282144 558884
rect 67456 558764 67508 558816
rect 201500 558764 201552 558816
rect 220084 558764 220136 558816
rect 229376 558764 229428 558816
rect 79508 558696 79560 558748
rect 88892 558696 88944 558748
rect 98552 558696 98604 558748
rect 104900 558696 104952 558748
rect 125508 558696 125560 558748
rect 208492 558696 208544 558748
rect 211160 558696 211212 558748
rect 217968 558696 218020 558748
rect 225972 558696 226024 558748
rect 234620 558696 234672 558748
rect 78496 558628 78548 558680
rect 87880 558628 87932 558680
rect 97080 558628 97132 558680
rect 77392 558560 77444 558612
rect 86684 558560 86736 558612
rect 75920 558492 75972 558544
rect 85396 558492 85448 558544
rect 94872 558560 94924 558612
rect 102048 558628 102100 558680
rect 140044 558628 140096 558680
rect 220728 558671 220780 558680
rect 220728 558637 220737 558671
rect 220737 558637 220771 558671
rect 220771 558637 220780 558671
rect 220728 558628 220780 558637
rect 227260 558628 227312 558680
rect 236000 558628 236052 558680
rect 283932 558832 283984 558884
rect 317420 558832 317472 558884
rect 326344 558832 326396 558884
rect 334256 558832 334308 558884
rect 343640 558832 343692 558884
rect 344744 558832 344796 558884
rect 344836 558832 344888 558884
rect 353300 558832 353352 558884
rect 446404 558832 446456 558884
rect 480536 558832 480588 558884
rect 284208 558764 284260 558816
rect 320272 558764 320324 558816
rect 332508 558764 332560 558816
rect 341248 558764 341300 558816
rect 350540 558764 350592 558816
rect 441620 558764 441672 558816
rect 457352 558764 457404 558816
rect 466552 558764 466604 558816
rect 475476 558764 475528 558816
rect 483020 558764 483072 558816
rect 284116 558696 284168 558748
rect 320180 558696 320232 558748
rect 324964 558696 325016 558748
rect 334256 558696 334308 558748
rect 336280 558696 336332 558748
rect 345756 558696 345808 558748
rect 349344 558696 349396 558748
rect 453672 558696 453724 558748
rect 462596 558696 462648 558748
rect 472164 558696 472216 558748
rect 481640 558696 481692 558748
rect 322848 558628 322900 558680
rect 327724 558628 327776 558680
rect 80796 558424 80848 558476
rect 86684 558424 86736 558476
rect 95700 558492 95752 558544
rect 102784 558560 102836 558612
rect 104808 558560 104860 558612
rect 144184 558560 144236 558612
rect 212540 558560 212592 558612
rect 213092 558560 213144 558612
rect 222292 558560 222344 558612
rect 231860 558560 231912 558612
rect 292580 558560 292632 558612
rect 323492 558560 323544 558612
rect 333152 558560 333204 558612
rect 333888 558560 333940 558612
rect 335912 558628 335964 558680
rect 344836 558628 344888 558680
rect 336280 558560 336332 558612
rect 336740 558560 336792 558612
rect 337752 558560 337804 558612
rect 346492 558628 346544 558680
rect 356060 558628 356112 558680
rect 418252 558628 418304 558680
rect 454040 558628 454092 558680
rect 454684 558628 454736 558680
rect 354680 558560 354732 558612
rect 455972 558560 456024 558612
rect 465264 558628 465316 558680
rect 474832 558628 474884 558680
rect 462964 558560 463016 558612
rect 468668 558560 468720 558612
rect 475476 558560 475528 558612
rect 484400 558560 484452 558612
rect 104164 558492 104216 558544
rect 108488 558492 108540 558544
rect 148324 558492 148376 558544
rect 218796 558492 218848 558544
rect 228088 558492 228140 558544
rect 237380 558492 237432 558544
rect 284024 558492 284076 558544
rect 302148 558492 302200 558544
rect 318800 558492 318852 558544
rect 383568 558492 383620 558544
rect 443092 558492 443144 558544
rect 451740 558492 451792 558544
rect 452384 558492 452436 558544
rect 89812 558424 89864 558476
rect 99380 558424 99432 558476
rect 100116 558424 100168 558476
rect 100576 558424 100628 558476
rect 140136 558424 140188 558476
rect 281908 558424 281960 558476
rect 329564 558424 329616 558476
rect 339040 558424 339092 558476
rect 73712 558356 73764 558408
rect 82912 558356 82964 558408
rect 97632 558356 97684 558408
rect 138664 558356 138716 558408
rect 211160 558356 211212 558408
rect 211896 558356 211948 558408
rect 221096 558356 221148 558408
rect 230480 558356 230532 558408
rect 81440 558288 81492 558340
rect 81992 558288 82044 558340
rect 91100 558288 91152 558340
rect 92296 558288 92348 558340
rect 137468 558288 137520 558340
rect 206376 558288 206428 558340
rect 215300 558288 215352 558340
rect 223948 558288 224000 558340
rect 233240 558288 233292 558340
rect 282000 558356 282052 558408
rect 328552 558356 328604 558408
rect 336740 558356 336792 558408
rect 346492 558424 346544 558476
rect 348240 558424 348292 558476
rect 357440 558424 357492 558476
rect 358084 558424 358136 558476
rect 452660 558424 452712 558476
rect 453948 558492 454000 558544
rect 461676 558492 461728 558544
rect 471336 558492 471388 558544
rect 480352 558492 480404 558544
rect 459468 558424 459520 558476
rect 468024 558424 468076 558476
rect 468760 558424 468812 558476
rect 470048 558424 470100 558476
rect 477592 558424 477644 558476
rect 238760 558288 238812 558340
rect 281816 558288 281868 558340
rect 330484 558288 330536 558340
rect 74264 558220 74316 558272
rect 137376 558220 137428 558272
rect 194416 558220 194468 558272
rect 313740 558220 313792 558272
rect 322848 558220 322900 558272
rect 332508 558220 332560 558272
rect 333888 558288 333940 558340
rect 342536 558288 342588 558340
rect 348424 558356 348476 558408
rect 359464 558356 359516 558408
rect 476120 558356 476172 558408
rect 476304 558356 476356 558408
rect 477132 558356 477184 558408
rect 485780 558356 485832 558408
rect 349344 558288 349396 558340
rect 357716 558288 357768 558340
rect 359556 558288 359608 558340
rect 477500 558288 477552 558340
rect 339868 558220 339920 558272
rect 344744 558220 344796 558272
rect 352012 558220 352064 558272
rect 358176 558220 358228 558272
rect 476212 558220 476264 558272
rect 477592 558220 477644 558272
rect 478236 558220 478288 558272
rect 487160 558220 487212 558272
rect 72516 558152 72568 558204
rect 81440 558152 81492 558204
rect 83832 558152 83884 558204
rect 149704 558152 149756 558204
rect 203800 558152 203852 558204
rect 212540 558152 212592 558204
rect 231952 558152 232004 558204
rect 283564 558152 283616 558204
rect 447600 558152 447652 558204
rect 76840 558084 76892 558136
rect 145564 558084 145616 558136
rect 213920 558084 213972 558136
rect 283748 558084 283800 558136
rect 418252 558084 418304 558136
rect 449900 558084 449952 558136
rect 81256 558016 81308 558068
rect 152556 558016 152608 558068
rect 283840 558016 283892 558068
rect 418160 558016 418212 558068
rect 432604 558016 432656 558068
rect 451280 558016 451332 558068
rect 79324 557948 79376 558000
rect 152464 557948 152516 558000
rect 223580 557948 223632 558000
rect 282276 557948 282328 558000
rect 443644 557948 443696 558000
rect 478880 558152 478932 558204
rect 478972 558152 479024 558204
rect 488540 558152 488592 558204
rect 75000 557880 75052 557932
rect 84200 557880 84252 557932
rect 89812 557880 89864 557932
rect 93768 557880 93820 557932
rect 137284 557880 137336 557932
rect 202144 557880 202196 557932
rect 211160 557880 211212 557932
rect 282368 557880 282420 557932
rect 449164 557880 449216 557932
rect 483020 558084 483072 558136
rect 107660 557812 107712 557864
rect 208492 557812 208544 557864
rect 282460 557812 282512 557864
rect 89352 557744 89404 557796
rect 97080 557744 97132 557796
rect 106280 557744 106332 557796
rect 121368 557744 121420 557796
rect 206376 557744 206428 557796
rect 207664 557744 207716 557796
rect 217968 557744 218020 557796
rect 282552 557744 282604 557796
rect 91100 557676 91152 557728
rect 100024 557676 100076 557728
rect 100116 557676 100168 557728
rect 108304 557676 108356 557728
rect 117228 557676 117280 557728
rect 203800 557676 203852 557728
rect 204904 557676 204956 557728
rect 213920 557676 213972 557728
rect 282644 557676 282696 557728
rect 92480 557608 92532 557660
rect 100852 557608 100904 557660
rect 84200 557540 84252 557592
rect 93584 557540 93636 557592
rect 107476 557540 107528 557592
rect 129740 557608 129792 557660
rect 210516 557608 210568 557660
rect 220084 557608 220136 557660
rect 282736 557608 282788 557660
rect 447784 557812 447836 557864
rect 481640 558016 481692 558068
rect 458272 557948 458324 558000
rect 459468 557948 459520 558000
rect 460848 557948 460900 558000
rect 468760 557948 468812 558000
rect 478972 557948 479024 558000
rect 454684 557880 454736 557932
rect 464344 557880 464396 557932
rect 488540 557880 488592 557932
rect 487160 557812 487212 557864
rect 451924 557744 451976 557796
rect 484400 557744 484452 557796
rect 450544 557676 450596 557728
rect 483112 557676 483164 557728
rect 453488 557608 453540 557660
rect 485780 557608 485832 557660
rect 141424 557540 141476 557592
rect 209044 557540 209096 557592
rect 218796 557540 218848 557592
rect 282828 557540 282880 557592
rect 418344 557540 418396 557592
rect 432512 557540 432564 557592
rect 441620 557540 441672 557592
rect 454040 557540 454092 557592
rect 459652 557540 459704 557592
rect 464252 557540 464304 557592
rect 473452 557540 473504 557592
rect 474648 557540 474700 557592
rect 476304 557540 476356 557592
rect 476396 557540 476448 557592
rect 483020 557540 483072 557592
rect 131764 557472 131816 557524
rect 283472 557472 283524 557524
rect 96528 545028 96580 545080
rect 189632 545028 189684 545080
rect 94136 544960 94188 545012
rect 188436 544960 188488 545012
rect 102048 544892 102100 544944
rect 197912 544892 197964 544944
rect 92112 544824 92164 544876
rect 188528 544824 188580 544876
rect 89996 544756 90048 544808
rect 188620 544756 188672 544808
rect 106188 544688 106240 544740
rect 206192 544688 206244 544740
rect 87972 544620 88024 544672
rect 188712 544620 188764 544672
rect 110328 544552 110380 544604
rect 212448 544552 212500 544604
rect 85856 544484 85908 544536
rect 188804 544484 188856 544536
rect 83832 544416 83884 544468
rect 188896 544416 188948 544468
rect 81716 544348 81768 544400
rect 195980 544348 196032 544400
rect 86776 544280 86828 544332
rect 173072 544280 173124 544332
rect 88248 544212 88300 544264
rect 175096 544212 175148 544264
rect 86868 544144 86920 544196
rect 170956 544144 171008 544196
rect 85488 544076 85540 544128
rect 168840 544076 168892 544128
rect 82728 544008 82780 544060
rect 164700 544008 164752 544060
rect 73068 543940 73120 543992
rect 148140 543940 148192 543992
rect 57888 543872 57940 543924
rect 112812 543872 112864 543924
rect 57796 543804 57848 543856
rect 110788 543804 110840 543856
rect 220728 543736 220780 543788
rect 71688 543668 71740 543720
rect 75460 543668 75512 543720
rect 75828 543668 75880 543720
rect 145564 543668 145616 543720
rect 152556 543668 152608 543720
rect 162676 543668 162728 543720
rect 205548 543668 205600 543720
rect 218704 543668 218756 543720
rect 220544 543668 220596 543720
rect 227628 543668 227680 543720
rect 258080 543668 258132 543720
rect 78588 543600 78640 543652
rect 156420 543600 156472 543652
rect 206928 543600 206980 543652
rect 220728 543600 220780 543652
rect 229008 543600 229060 543652
rect 260196 543600 260248 543652
rect 61016 543532 61068 543584
rect 62028 543532 62080 543584
rect 65156 543532 65208 543584
rect 66168 543532 66220 543584
rect 70308 543532 70360 543584
rect 71320 543532 71372 543584
rect 79968 543532 80020 543584
rect 152464 543532 152516 543584
rect 158536 543532 158588 543584
rect 208308 543532 208360 543584
rect 222844 543532 222896 543584
rect 230388 543532 230440 543584
rect 262220 543532 262272 543584
rect 57428 543464 57480 543516
rect 102508 543464 102560 543516
rect 127348 543464 127400 543516
rect 209044 543464 209096 543516
rect 209688 543464 209740 543516
rect 224868 543464 224920 543516
rect 231768 543464 231820 543516
rect 264336 543464 264388 543516
rect 57520 543396 57572 543448
rect 104532 543396 104584 543448
rect 123208 543396 123260 543448
rect 207664 543396 207716 543448
rect 210976 543396 211028 543448
rect 226984 543396 227036 543448
rect 233148 543396 233200 543448
rect 266452 543396 266504 543448
rect 57612 543328 57664 543380
rect 106648 543328 106700 543380
rect 119068 543328 119120 543380
rect 204904 543328 204956 543380
rect 212356 543328 212408 543380
rect 231124 543328 231176 543380
rect 233056 543328 233108 543380
rect 268476 543328 268528 543380
rect 91008 543260 91060 543312
rect 179236 543260 179288 543312
rect 215208 543260 215260 543312
rect 235264 543260 235316 543312
rect 235908 543260 235960 543312
rect 272616 543260 272668 543312
rect 57704 543192 57756 543244
rect 108672 543192 108724 543244
rect 114928 543192 114980 543244
rect 202144 543192 202196 543244
rect 211068 543192 211120 543244
rect 229100 543192 229152 543244
rect 234528 543192 234580 543244
rect 270592 543192 270644 543244
rect 93676 543124 93728 543176
rect 183376 543124 183428 543176
rect 202788 543124 202840 543176
rect 214564 543124 214616 543176
rect 216588 543124 216640 543176
rect 237380 543124 237432 543176
rect 238668 543124 238720 543176
rect 276756 543124 276808 543176
rect 57244 543056 57296 543108
rect 79692 543056 79744 543108
rect 95056 543056 95108 543108
rect 187516 543056 187568 543108
rect 204168 543056 204220 543108
rect 213828 543056 213880 543108
rect 233240 543056 233292 543108
rect 237288 543056 237340 543108
rect 274732 543056 274784 543108
rect 67548 542988 67600 543040
rect 98368 542988 98420 543040
rect 99288 542988 99340 543040
rect 193772 542988 193824 543040
rect 216588 542988 216640 543040
rect 217876 542988 217928 543040
rect 239404 542988 239456 543040
rect 240048 542988 240100 543040
rect 278872 542988 278924 543040
rect 57336 542920 57388 542972
rect 100392 542920 100444 542972
rect 108580 542920 108632 542972
rect 144000 542920 144052 542972
rect 144184 542920 144236 542972
rect 204168 542920 204220 542972
rect 226156 542920 226208 542972
rect 256056 542920 256108 542972
rect 105544 542852 105596 542904
rect 139860 542852 139912 542904
rect 140136 542852 140188 542904
rect 195888 542852 195940 542904
rect 226248 542852 226300 542904
rect 253940 542852 253992 542904
rect 104164 542784 104216 542836
rect 137744 542784 137796 542836
rect 138664 542784 138716 542836
rect 191748 542784 191800 542836
rect 223488 542784 223540 542836
rect 249800 542784 249852 542836
rect 102784 542716 102836 542768
rect 135720 542716 135772 542768
rect 137284 542716 137336 542768
rect 185492 542716 185544 542768
rect 224684 542716 224736 542768
rect 251916 542716 251968 542768
rect 70216 542648 70268 542700
rect 73436 542648 73488 542700
rect 100024 542648 100076 542700
rect 131488 542648 131540 542700
rect 131764 542648 131816 542700
rect 177212 542648 177264 542700
rect 222108 542648 222160 542700
rect 247776 542648 247828 542700
rect 101404 542580 101456 542632
rect 133604 542580 133656 542632
rect 137468 542580 137520 542632
rect 181352 542580 181404 542632
rect 220544 542580 220596 542632
rect 245660 542580 245712 542632
rect 108304 542512 108356 542564
rect 146024 542512 146076 542564
rect 106924 542444 106976 542496
rect 141884 542444 141936 542496
rect 152280 542512 152332 542564
rect 154396 542512 154448 542564
rect 149704 542444 149756 542496
rect 166816 542512 166868 542564
rect 217968 542512 218020 542564
rect 241520 542512 241572 542564
rect 219348 542444 219400 542496
rect 243544 542444 243596 542496
rect 137376 542376 137428 542428
rect 150164 542376 150216 542428
rect 160560 542376 160612 542428
rect 281724 539520 281776 539572
rect 464344 539520 464396 539572
rect 281724 538160 281776 538212
rect 454684 538160 454736 538212
rect 281724 535372 281776 535424
rect 453488 535372 453540 535424
rect 281724 534012 281776 534064
rect 451924 534012 451976 534064
rect 281724 531224 281776 531276
rect 450544 531224 450596 531276
rect 281724 529864 281776 529916
rect 449164 529864 449216 529916
rect 281724 527076 281776 527128
rect 447784 527076 447836 527128
rect 281724 525716 281776 525768
rect 446404 525716 446456 525768
rect 281724 522928 281776 522980
rect 443644 522928 443696 522980
rect 281724 521568 281776 521620
rect 359556 521568 359608 521620
rect 281724 518848 281776 518900
rect 359464 518848 359516 518900
rect 281724 517420 281776 517472
rect 358176 517420 358228 517472
rect 281724 514700 281776 514752
rect 356704 514700 356756 514752
rect 281724 513272 281776 513324
rect 473360 513272 473412 513324
rect 281724 510552 281776 510604
rect 471980 510552 472032 510604
rect 281724 509192 281776 509244
rect 470600 509192 470652 509244
rect 281724 506404 281776 506456
rect 469220 506404 469272 506456
rect 281724 505044 281776 505096
rect 467932 505044 467984 505096
rect 281724 502256 281776 502308
rect 467840 502256 467892 502308
rect 281724 500896 281776 500948
rect 466460 500896 466512 500948
rect 281724 499468 281776 499520
rect 465080 499468 465132 499520
rect 281724 496748 281776 496800
rect 463700 496748 463752 496800
rect 281724 495388 281776 495440
rect 462320 495388 462372 495440
rect 281724 492600 281776 492652
rect 461032 492600 461084 492652
rect 281724 491240 281776 491292
rect 460940 491240 460992 491292
rect 281724 488452 281776 488504
rect 459560 488452 459612 488504
rect 281724 487092 281776 487144
rect 458180 487092 458232 487144
rect 281724 484304 281776 484356
rect 456800 484304 456852 484356
rect 281724 482944 281776 482996
rect 455420 482944 455472 482996
rect 281724 480156 281776 480208
rect 453396 480156 453448 480208
rect 281724 478796 281776 478848
rect 358084 478796 358136 478848
rect 281724 476008 281776 476060
rect 452660 476008 452712 476060
rect 281724 474648 281776 474700
rect 358912 474648 358964 474700
rect 281724 471928 281776 471980
rect 357532 471928 357584 471980
rect 281724 470500 281776 470552
rect 356060 470500 356112 470552
rect 281724 467780 281776 467832
rect 354680 467780 354732 467832
rect 281724 466352 281776 466404
rect 353300 466352 353352 466404
rect 281724 463632 281776 463684
rect 352012 463632 352064 463684
rect 281724 462272 281776 462324
rect 352196 462272 352248 462324
rect 281724 459484 281776 459536
rect 350540 459484 350592 459536
rect 281724 458124 281776 458176
rect 349160 458124 349212 458176
rect 281724 455336 281776 455388
rect 347780 455336 347832 455388
rect 281724 453976 281776 454028
rect 346400 453976 346452 454028
rect 281724 452548 281776 452600
rect 345020 452548 345072 452600
rect 281724 449828 281776 449880
rect 343732 449828 343784 449880
rect 281724 448468 281776 448520
rect 343640 448468 343692 448520
rect 281724 445680 281776 445732
rect 342260 445680 342312 445732
rect 281724 444320 281776 444372
rect 340880 444320 340932 444372
rect 281724 441532 281776 441584
rect 339500 441532 339552 441584
rect 281724 440172 281776 440224
rect 338120 440172 338172 440224
rect 281724 437384 281776 437436
rect 336832 437384 336884 437436
rect 281724 436024 281776 436076
rect 336740 436024 336792 436076
rect 281724 433236 281776 433288
rect 335360 433236 335412 433288
rect 281724 431876 281776 431928
rect 333980 431876 334032 431928
rect 281724 429088 281776 429140
rect 332600 429088 332652 429140
rect 281724 427728 281776 427780
rect 331220 427728 331272 427780
rect 281724 425008 281776 425060
rect 329932 425008 329984 425060
rect 281724 423580 281776 423632
rect 329840 423580 329892 423632
rect 281724 420860 281776 420912
rect 328460 420860 328512 420912
rect 281724 419432 281776 419484
rect 327080 419432 327132 419484
rect 281724 418072 281776 418124
rect 325700 418072 325752 418124
rect 281724 415352 281776 415404
rect 324320 415352 324372 415404
rect 281724 413924 281776 413976
rect 322940 413924 322992 413976
rect 383568 413244 383620 413296
rect 405004 413244 405056 413296
rect 405004 412632 405056 412684
rect 513380 412632 513432 412684
rect 285312 412428 285364 412480
rect 316040 412428 316092 412480
rect 281632 412360 281684 412412
rect 324964 412360 325016 412412
rect 281540 412292 281592 412344
rect 326344 412292 326396 412344
rect 327724 412224 327776 412276
rect 283104 412156 283156 412208
rect 438584 412156 438636 412208
rect 283012 412088 283064 412140
rect 438492 412088 438544 412140
rect 283196 412020 283248 412072
rect 438676 412020 438728 412072
rect 283288 411952 283340 412004
rect 445760 411952 445812 412004
rect 285404 411884 285456 411936
rect 453304 411884 453356 411936
rect 281724 411340 281776 411392
rect 282000 411340 282052 411392
rect 282000 411204 282052 411256
rect 321560 411204 321612 411256
rect 285220 410796 285272 410848
rect 438124 410796 438176 410848
rect 285128 410728 285180 410780
rect 438216 410728 438268 410780
rect 285036 410660 285088 410712
rect 438308 410660 438360 410712
rect 283380 410592 283432 410644
rect 438768 410592 438820 410644
rect 282000 410567 282052 410576
rect 282000 410533 282009 410567
rect 282009 410533 282043 410567
rect 282043 410533 282052 410567
rect 282000 410524 282052 410533
rect 282920 410524 282972 410576
rect 438400 410524 438452 410576
rect 281540 404132 281592 404184
rect 282000 404132 282052 404184
rect 281540 397060 281592 397112
rect 283472 397060 283524 397112
rect 281908 378020 281960 378072
rect 285404 378020 285456 378072
rect 282828 376660 282880 376712
rect 294696 376660 294748 376712
rect 282828 373940 282880 373992
rect 291844 373940 291896 373992
rect 282828 372512 282880 372564
rect 290464 372512 290516 372564
rect 282368 371016 282420 371068
rect 287704 371016 287756 371068
rect 282276 368024 282328 368076
rect 286324 368024 286376 368076
rect 281724 365780 281776 365832
rect 284944 365780 284996 365832
rect 282828 364284 282880 364336
rect 294604 364284 294656 364336
rect 281908 362856 281960 362908
rect 285312 362856 285364 362908
rect 281908 360136 281960 360188
rect 285220 360136 285272 360188
rect 281724 357620 281776 357672
rect 285128 357620 285180 357672
rect 282092 355852 282144 355904
rect 285036 355852 285088 355904
rect 281540 346060 281592 346112
rect 283288 346060 283340 346112
rect 282828 343544 282880 343596
rect 302884 343544 302936 343596
rect 281540 341300 281592 341352
rect 283380 341300 283432 341352
rect 281724 339260 281776 339312
rect 284208 339260 284260 339312
rect 281540 337560 281592 337612
rect 284116 337560 284168 337612
rect 281632 335180 281684 335232
rect 284024 335180 284076 335232
rect 281540 333208 281592 333260
rect 283932 333208 283984 333260
rect 281540 331100 281592 331152
rect 283840 331100 283892 331152
rect 281540 329060 281592 329112
rect 283748 329060 283800 329112
rect 281540 327020 281592 327072
rect 283656 327020 283708 327072
rect 281540 325048 281592 325100
rect 283564 325048 283616 325100
rect 135996 318996 136048 319048
rect 136548 318996 136600 319048
rect 59360 318928 59412 318980
rect 60280 318928 60332 318980
rect 30288 318724 30340 318776
rect 70952 318724 71004 318776
rect 115848 318724 115900 318776
rect 145656 318792 145708 318844
rect 138112 318724 138164 318776
rect 31668 318656 31720 318708
rect 71780 318656 71832 318708
rect 99656 318656 99708 318708
rect 105176 318656 105228 318708
rect 117136 318656 117188 318708
rect 30196 318588 30248 318640
rect 71320 318588 71372 318640
rect 118516 318588 118568 318640
rect 148600 318724 148652 318776
rect 150348 318724 150400 318776
rect 175832 318724 175884 318776
rect 210976 318724 211028 318776
rect 217692 318724 217744 318776
rect 293224 318724 293276 318776
rect 313280 318724 313332 318776
rect 405004 318724 405056 318776
rect 443092 318724 443144 318776
rect 149888 318656 149940 318708
rect 162124 318656 162176 318708
rect 163872 318656 163924 318708
rect 246304 318656 246356 318708
rect 145012 318588 145064 318640
rect 155776 318588 155828 318640
rect 178592 318588 178644 318640
rect 186780 318588 186832 318640
rect 193864 318588 193916 318640
rect 198832 318588 198884 318640
rect 291844 318588 291896 318640
rect 23388 318520 23440 318572
rect 27528 318452 27580 318504
rect 64604 318520 64656 318572
rect 111800 318520 111852 318572
rect 133144 318520 133196 318572
rect 134248 318520 134300 318572
rect 169024 318520 169076 318572
rect 177304 318520 177356 318572
rect 189080 318520 189132 318572
rect 193496 318520 193548 318572
rect 289084 318520 289136 318572
rect 68652 318452 68704 318504
rect 82084 318452 82136 318504
rect 90180 318452 90232 318504
rect 124772 318452 124824 318504
rect 170588 318452 170640 318504
rect 272892 318452 272944 318504
rect 22008 318384 22060 318436
rect 67732 318384 67784 318436
rect 79324 318384 79376 318436
rect 87512 318384 87564 318436
rect 108580 318384 108632 318436
rect 128636 318384 128688 318436
rect 130200 318384 130252 318436
rect 167644 318384 167696 318436
rect 171968 318384 172020 318436
rect 279424 318384 279476 318436
rect 20628 318316 20680 318368
rect 67364 318316 67416 318368
rect 82728 318316 82780 318368
rect 90640 318316 90692 318368
rect 126152 318316 126204 318368
rect 164884 318316 164936 318368
rect 165160 318316 165212 318368
rect 174636 318316 174688 318368
rect 286324 318316 286376 318368
rect 21916 318248 21968 318300
rect 60740 318248 60792 318300
rect 70032 318248 70084 318300
rect 75184 318248 75236 318300
rect 87052 318248 87104 318300
rect 107292 318248 107344 318300
rect 127440 318248 127492 318300
rect 166356 318248 166408 318300
rect 175924 318248 175976 318300
rect 304264 318248 304316 318300
rect 313280 318180 313332 318232
rect 17868 318112 17920 318164
rect 66444 318112 66496 318164
rect 13728 318044 13780 318096
rect 60372 318044 60424 318096
rect 60740 318044 60792 318096
rect 68192 318044 68244 318096
rect 74448 318044 74500 318096
rect 87972 318112 88024 318164
rect 122104 318112 122156 318164
rect 167000 318112 167052 318164
rect 168288 318112 168340 318164
rect 87604 318044 87656 318096
rect 89812 318044 89864 318096
rect 98736 318044 98788 318096
rect 102416 318044 102468 318096
rect 102784 318044 102836 318096
rect 103336 318044 103388 318096
rect 104992 318044 105044 318096
rect 105728 318044 105780 318096
rect 107752 318044 107804 318096
rect 108856 318044 108908 318096
rect 120724 318044 120776 318096
rect 153844 318044 153896 318096
rect 155316 318044 155368 318096
rect 155776 318044 155828 318096
rect 167460 318044 167512 318096
rect 168196 318044 168248 318096
rect 38476 317976 38528 318028
rect 74540 317976 74592 318028
rect 88248 317976 88300 318028
rect 92940 317976 92992 318028
rect 110420 317976 110472 318028
rect 127624 317976 127676 318028
rect 166264 317976 166316 318028
rect 167920 317976 167972 318028
rect 168748 318044 168800 318096
rect 169576 318044 169628 318096
rect 248696 318112 248748 318164
rect 249616 318112 249668 318164
rect 250076 318112 250128 318164
rect 250996 318112 251048 318164
rect 251364 318112 251416 318164
rect 252376 318112 252428 318164
rect 252744 318112 252796 318164
rect 253664 318112 253716 318164
rect 254032 318112 254084 318164
rect 255044 318112 255096 318164
rect 255412 318112 255464 318164
rect 256424 318112 256476 318164
rect 256792 318112 256844 318164
rect 257804 318112 257856 318164
rect 258080 318112 258132 318164
rect 259184 318112 259236 318164
rect 259920 318112 259972 318164
rect 260748 318112 260800 318164
rect 261852 318112 261904 318164
rect 262128 318112 262180 318164
rect 263324 318112 263376 318164
rect 263508 318112 263560 318164
rect 264704 318112 264756 318164
rect 264888 318112 264940 318164
rect 265256 318112 265308 318164
rect 266268 318112 266320 318164
rect 267096 318112 267148 318164
rect 267556 318112 267608 318164
rect 268016 318112 268068 318164
rect 269028 318112 269080 318164
rect 269304 318112 269356 318164
rect 270408 318112 270460 318164
rect 270684 318112 270736 318164
rect 271788 318112 271840 318164
rect 272524 318112 272576 318164
rect 273076 318112 273128 318164
rect 273352 318112 273404 318164
rect 274548 318112 274600 318164
rect 275652 318112 275704 318164
rect 529388 318112 529440 318164
rect 268476 318044 268528 318096
rect 268936 318044 268988 318096
rect 269764 318044 269816 318096
rect 270316 318044 270368 318096
rect 271144 318044 271196 318096
rect 271696 318044 271748 318096
rect 272064 318044 272116 318096
rect 273168 318044 273220 318096
rect 273812 318044 273864 318096
rect 274456 318044 274508 318096
rect 274732 318044 274784 318096
rect 275928 318044 275980 318096
rect 276480 318044 276532 318096
rect 277216 318044 277268 318096
rect 529480 318044 529532 318096
rect 169208 317976 169260 318028
rect 37188 317908 37240 317960
rect 73620 317908 73672 317960
rect 79416 317908 79468 317960
rect 83464 317908 83516 317960
rect 85488 317908 85540 317960
rect 92020 317908 92072 317960
rect 130660 317908 130712 317960
rect 134616 317908 134668 317960
rect 134708 317908 134760 317960
rect 146760 317908 146812 317960
rect 147588 317908 147640 317960
rect 147680 317908 147732 317960
rect 148876 317908 148928 317960
rect 44088 317840 44140 317892
rect 76288 317840 76340 317892
rect 89628 317840 89680 317892
rect 93400 317840 93452 317892
rect 98276 317840 98328 317892
rect 100116 317840 100168 317892
rect 127072 317840 127124 317892
rect 128268 317840 128320 317892
rect 129280 317840 129332 317892
rect 170128 317908 170180 317960
rect 171048 317908 171100 317960
rect 172796 317908 172848 317960
rect 173716 317908 173768 317960
rect 174176 317908 174228 317960
rect 175096 317908 175148 317960
rect 176844 317908 176896 317960
rect 177856 317908 177908 317960
rect 178224 317908 178276 317960
rect 179236 317908 179288 317960
rect 179512 317908 179564 317960
rect 180616 317908 180668 317960
rect 182272 317976 182324 318028
rect 183376 317976 183428 318028
rect 183560 317976 183612 318028
rect 184756 317976 184808 318028
rect 184940 317976 184992 318028
rect 186136 317976 186188 318028
rect 186320 317976 186372 318028
rect 187424 317976 187476 318028
rect 188528 317976 188580 318028
rect 188988 317976 189040 318028
rect 189908 317976 189960 318028
rect 190368 317976 190420 318028
rect 191196 317976 191248 318028
rect 191656 317976 191708 318028
rect 192116 317976 192168 318028
rect 192944 317976 192996 318028
rect 193956 317976 194008 318028
rect 194508 317976 194560 318028
rect 194784 317976 194836 318028
rect 195704 317976 195756 318028
rect 196624 317976 196676 318028
rect 197176 317976 197228 318028
rect 197544 317976 197596 318028
rect 198464 317976 198516 318028
rect 199292 317976 199344 318028
rect 200028 317976 200080 318028
rect 200212 317976 200264 318028
rect 201224 317976 201276 318028
rect 201592 317976 201644 318028
rect 202604 317976 202656 318028
rect 202880 317976 202932 318028
rect 203984 317976 204036 318028
rect 205364 317976 205416 318028
rect 205548 317976 205600 318028
rect 206008 317976 206060 318028
rect 206836 317976 206888 318028
rect 207388 317976 207440 318028
rect 208124 317976 208176 318028
rect 208768 317976 208820 318028
rect 209596 317976 209648 318028
rect 210056 317976 210108 318028
rect 211068 317976 211120 318028
rect 211436 317976 211488 318028
rect 212448 317976 212500 318028
rect 213184 317976 213236 318028
rect 213736 317976 213788 318028
rect 214104 317976 214156 318028
rect 215116 317976 215168 318028
rect 215944 317976 215996 318028
rect 216496 317976 216548 318028
rect 216772 317976 216824 318028
rect 217968 317976 218020 318028
rect 295984 317976 296036 318028
rect 153108 317840 153160 317892
rect 176016 317840 176068 317892
rect 184204 317908 184256 317960
rect 184296 317908 184348 317960
rect 38568 317772 38620 317824
rect 74080 317772 74132 317824
rect 84844 317772 84896 317824
rect 91560 317772 91612 317824
rect 113088 317772 113140 317824
rect 127900 317772 127952 317824
rect 148416 317772 148468 317824
rect 149060 317772 149112 317824
rect 155224 317772 155276 317824
rect 173164 317772 173216 317824
rect 173256 317772 173308 317824
rect 185584 317840 185636 317892
rect 187148 317908 187200 317960
rect 187608 317908 187660 317960
rect 192576 317908 192628 317960
rect 193128 317908 193180 317960
rect 195244 317908 195296 317960
rect 195888 317908 195940 317960
rect 196164 317908 196216 317960
rect 197268 317908 197320 317960
rect 200672 317908 200724 317960
rect 201408 317908 201460 317960
rect 203340 317908 203392 317960
rect 204168 317908 204220 317960
rect 207848 317908 207900 317960
rect 208308 317908 208360 317960
rect 212816 317908 212868 317960
rect 213828 317908 213880 317960
rect 215484 317908 215536 317960
rect 216588 317908 216640 317960
rect 217232 317908 217284 317960
rect 217876 317908 217928 317960
rect 218152 317908 218204 317960
rect 219348 317908 219400 317960
rect 219992 317908 220044 317960
rect 220636 317908 220688 317960
rect 220820 317908 220872 317960
rect 222016 317908 222068 317960
rect 222660 317908 222712 317960
rect 223396 317908 223448 317960
rect 223580 317908 223632 317960
rect 224868 317908 224920 317960
rect 225328 317908 225380 317960
rect 226156 317908 226208 317960
rect 226708 317908 226760 317960
rect 227536 317908 227588 317960
rect 227996 317908 228048 317960
rect 228916 317908 228968 317960
rect 296076 317908 296128 317960
rect 253112 317840 253164 317892
rect 253204 317840 253256 317892
rect 253848 317840 253900 317892
rect 254492 317840 254544 317892
rect 255228 317840 255280 317892
rect 255872 317840 255924 317892
rect 256608 317840 256660 317892
rect 257252 317840 257304 317892
rect 257988 317840 258040 317892
rect 258540 317840 258592 317892
rect 259368 317840 259420 317892
rect 260840 317840 260892 317892
rect 261944 317840 261996 317892
rect 263968 317840 264020 317892
rect 264888 317840 264940 317892
rect 266636 317840 266688 317892
rect 267648 317840 267700 317892
rect 271144 317840 271196 317892
rect 275284 317840 275336 317892
rect 276112 317840 276164 317892
rect 277308 317840 277360 317892
rect 277860 317840 277912 317892
rect 278596 317840 278648 317892
rect 278780 317840 278832 317892
rect 280068 317840 280120 317892
rect 180892 317772 180944 317824
rect 181996 317772 182048 317824
rect 185400 317772 185452 317824
rect 189724 317772 189776 317824
rect 250444 317772 250496 317824
rect 261300 317772 261352 317824
rect 262128 317772 262180 317824
rect 275192 317772 275244 317824
rect 275836 317772 275888 317824
rect 277400 317772 277452 317824
rect 278688 317772 278740 317824
rect 45468 317704 45520 317756
rect 76748 317704 76800 317756
rect 99196 317704 99248 317756
rect 100024 317704 100076 317756
rect 101036 317704 101088 317756
rect 102784 317704 102836 317756
rect 106832 317704 106884 317756
rect 107476 317704 107528 317756
rect 108212 317704 108264 317756
rect 108948 317704 109000 317756
rect 50988 317636 51040 317688
rect 78956 317636 79008 317688
rect 100576 317636 100628 317688
rect 104164 317636 104216 317688
rect 119436 317636 119488 317688
rect 46848 317568 46900 317620
rect 77208 317568 77260 317620
rect 77944 317568 77996 317620
rect 85304 317568 85356 317620
rect 91008 317568 91060 317620
rect 94228 317568 94280 317620
rect 102324 317568 102376 317620
rect 104256 317568 104308 317620
rect 106372 317568 106424 317620
rect 107568 317568 107620 317620
rect 123484 317568 123536 317620
rect 124128 317568 124180 317620
rect 131948 317636 132000 317688
rect 138020 317636 138072 317688
rect 140780 317636 140832 317688
rect 145564 317636 145616 317688
rect 152280 317704 152332 317756
rect 159456 317704 159508 317756
rect 152556 317636 152608 317688
rect 160376 317704 160428 317756
rect 162492 317704 162544 317756
rect 180064 317704 180116 317756
rect 188068 317704 188120 317756
rect 253296 317704 253348 317756
rect 262588 317704 262640 317756
rect 263508 317704 263560 317756
rect 171784 317636 171836 317688
rect 53748 317500 53800 317552
rect 79876 317500 79928 317552
rect 82176 317500 82228 317552
rect 88892 317500 88944 317552
rect 92388 317500 92440 317552
rect 94688 317500 94740 317552
rect 97448 317500 97500 317552
rect 97908 317500 97960 317552
rect 109500 317500 109552 317552
rect 110144 317500 110196 317552
rect 57888 317432 57940 317484
rect 81716 317432 81768 317484
rect 86224 317432 86276 317484
rect 88432 317432 88484 317484
rect 90364 317432 90416 317484
rect 91100 317432 91152 317484
rect 93768 317432 93820 317484
rect 95148 317432 95200 317484
rect 96988 317432 97040 317484
rect 97724 317432 97776 317484
rect 103704 317432 103756 317484
rect 104716 317432 104768 317484
rect 109040 317432 109092 317484
rect 110328 317432 110380 317484
rect 110880 317432 110932 317484
rect 111616 317432 111668 317484
rect 112260 317432 112312 317484
rect 112996 317432 113048 317484
rect 113548 317432 113600 317484
rect 114376 317432 114428 317484
rect 114928 317432 114980 317484
rect 115848 317432 115900 317484
rect 116216 317432 116268 317484
rect 116952 317432 117004 317484
rect 118976 317432 119028 317484
rect 119896 317432 119948 317484
rect 120264 317432 120316 317484
rect 121276 317432 121328 317484
rect 121644 317432 121696 317484
rect 122656 317432 122708 317484
rect 123024 317432 123076 317484
rect 123944 317432 123996 317484
rect 124312 317432 124364 317484
rect 125416 317432 125468 317484
rect 125692 317432 125744 317484
rect 126888 317432 126940 317484
rect 130384 317500 130436 317552
rect 128820 317432 128872 317484
rect 129648 317432 129700 317484
rect 129740 317432 129792 317484
rect 131028 317432 131080 317484
rect 126612 317364 126664 317416
rect 137928 317568 137980 317620
rect 148324 317568 148376 317620
rect 156604 317568 156656 317620
rect 156696 317568 156748 317620
rect 157064 317568 157116 317620
rect 157524 317568 157576 317620
rect 158628 317568 158680 317620
rect 158904 317568 158956 317620
rect 160008 317568 160060 317620
rect 166080 317568 166132 317620
rect 166816 317568 166868 317620
rect 133328 317500 133380 317552
rect 131488 317432 131540 317484
rect 132408 317432 132460 317484
rect 132868 317432 132920 317484
rect 133788 317432 133840 317484
rect 138296 317500 138348 317552
rect 139308 317500 139360 317552
rect 138664 317432 138716 317484
rect 139216 317432 139268 317484
rect 142252 317500 142304 317552
rect 143448 317500 143500 317552
rect 135904 317364 135956 317416
rect 140044 317432 140096 317484
rect 140596 317432 140648 317484
rect 141424 317432 141476 317484
rect 141976 317432 142028 317484
rect 142712 317432 142764 317484
rect 143356 317432 143408 317484
rect 144092 317432 144144 317484
rect 144736 317432 144788 317484
rect 145472 317432 145524 317484
rect 146208 317432 146260 317484
rect 146300 317432 146352 317484
rect 147496 317432 147548 317484
rect 151084 317500 151136 317552
rect 148140 317432 148192 317484
rect 148968 317432 149020 317484
rect 149520 317432 149572 317484
rect 150164 317432 150216 317484
rect 150808 317432 150860 317484
rect 151728 317432 151780 317484
rect 152188 317432 152240 317484
rect 153108 317432 153160 317484
rect 153476 317432 153528 317484
rect 154488 317432 154540 317484
rect 154856 317432 154908 317484
rect 155868 317432 155920 317484
rect 156236 317500 156288 317552
rect 157248 317500 157300 317552
rect 157984 317432 158036 317484
rect 158536 317432 158588 317484
rect 160284 317500 160336 317552
rect 161388 317500 161440 317552
rect 162032 317500 162084 317552
rect 162676 317500 162728 317552
rect 163412 317500 163464 317552
rect 164056 317500 164108 317552
rect 164332 317500 164384 317552
rect 165528 317500 165580 317552
rect 166540 317500 166592 317552
rect 182824 317636 182876 317688
rect 189080 317636 189132 317688
rect 189816 317636 189868 317688
rect 190736 317636 190788 317688
rect 191748 317636 191800 317688
rect 204720 317636 204772 317688
rect 205548 317636 205600 317688
rect 182732 317568 182784 317620
rect 204260 317500 204312 317552
rect 271236 317636 271288 317688
rect 218612 317568 218664 317620
rect 219256 317568 219308 317620
rect 219532 317568 219584 317620
rect 220728 317568 220780 317620
rect 221280 317568 221332 317620
rect 221924 317568 221976 317620
rect 222200 317568 222252 317620
rect 223488 317568 223540 317620
rect 224408 317568 224460 317620
rect 229376 317568 229428 317620
rect 230204 317568 230256 317620
rect 230756 317568 230808 317620
rect 231676 317568 231728 317620
rect 232044 317568 232096 317620
rect 232964 317568 233016 317620
rect 233424 317568 233476 317620
rect 234436 317568 234488 317620
rect 234804 317568 234856 317620
rect 235724 317568 235776 317620
rect 236092 317568 236144 317620
rect 237196 317568 237248 317620
rect 237472 317568 237524 317620
rect 238484 317568 238536 317620
rect 238852 317568 238904 317620
rect 239956 317568 240008 317620
rect 240140 317568 240192 317620
rect 241244 317568 241296 317620
rect 241980 317568 242032 317620
rect 242624 317568 242676 317620
rect 243268 317568 243320 317620
rect 244188 317568 244240 317620
rect 246028 317568 246080 317620
rect 246948 317568 247000 317620
rect 247316 317568 247368 317620
rect 248236 317568 248288 317620
rect 255964 317568 256016 317620
rect 224040 317500 224092 317552
rect 224684 317500 224736 317552
rect 229836 317500 229888 317552
rect 230388 317500 230440 317552
rect 232504 317500 232556 317552
rect 233148 317500 233200 317552
rect 235264 317500 235316 317552
rect 235908 317500 235960 317552
rect 236552 317500 236604 317552
rect 237104 317500 237156 317552
rect 237932 317500 237984 317552
rect 238668 317500 238720 317552
rect 239220 317500 239272 317552
rect 239864 317500 239916 317552
rect 240600 317500 240652 317552
rect 241428 317500 241480 317552
rect 241520 317500 241572 317552
rect 242716 317500 242768 317552
rect 244648 317500 244700 317552
rect 245568 317500 245620 317552
rect 259460 317500 259512 317552
rect 260564 317500 260616 317552
rect 159364 317432 159416 317484
rect 159916 317432 159968 317484
rect 160744 317432 160796 317484
rect 161296 317432 161348 317484
rect 161572 317432 161624 317484
rect 162768 317432 162820 317484
rect 162952 317432 163004 317484
rect 164148 317432 164200 317484
rect 164700 317432 164752 317484
rect 165436 317432 165488 317484
rect 165620 317432 165672 317484
rect 166908 317432 166960 317484
rect 171508 317432 171560 317484
rect 172336 317432 172388 317484
rect 175556 317432 175608 317484
rect 176476 317432 176528 317484
rect 179972 317432 180024 317484
rect 180524 317432 180576 317484
rect 198004 317432 198056 317484
rect 198648 317432 198700 317484
rect 201960 317432 202012 317484
rect 202788 317432 202840 317484
rect 159364 317296 159416 317348
rect 60740 315936 60792 315988
rect 61108 315936 61160 315988
rect 64880 315936 64932 315988
rect 65708 315936 65760 315988
rect 69112 315936 69164 315988
rect 69388 315936 69440 315988
rect 80152 315936 80204 315988
rect 80980 315936 81032 315988
rect 81532 315936 81584 315988
rect 82268 315936 82320 315988
rect 84292 315936 84344 315988
rect 84476 315936 84528 315988
rect 85580 315936 85632 315988
rect 86316 315936 86368 315988
rect 92572 315936 92624 315988
rect 93492 315936 93544 315988
rect 75000 315868 75052 315920
rect 75460 315868 75512 315920
rect 77576 315868 77628 315920
rect 78220 315868 78272 315920
rect 117872 315868 117924 315920
rect 118516 315868 118568 315920
rect 82912 315664 82964 315716
rect 83556 315664 83608 315716
rect 128360 315392 128412 315444
rect 129556 315392 129608 315444
rect 66812 313896 66864 313948
rect 66996 313896 67048 313948
rect 135168 311924 135220 311976
rect 137744 311856 137796 311908
rect 137928 311856 137980 311908
rect 140780 311788 140832 311840
rect 140964 311788 141016 311840
rect 78864 309136 78916 309188
rect 79048 309136 79100 309188
rect 86040 309136 86092 309188
rect 86132 309136 86184 309188
rect 135076 309179 135128 309188
rect 135076 309145 135085 309179
rect 135085 309145 135119 309179
rect 135119 309145 135128 309179
rect 135076 309136 135128 309145
rect 160744 309179 160796 309188
rect 160744 309145 160753 309179
rect 160753 309145 160787 309179
rect 160787 309145 160796 309179
rect 160744 309136 160796 309145
rect 66996 309068 67048 309120
rect 74448 309111 74500 309120
rect 74448 309077 74457 309111
rect 74457 309077 74491 309111
rect 74491 309077 74500 309111
rect 74448 309068 74500 309077
rect 77576 309111 77628 309120
rect 77576 309077 77585 309111
rect 77585 309077 77619 309111
rect 77619 309077 77628 309111
rect 77576 309068 77628 309077
rect 95424 309111 95476 309120
rect 95424 309077 95433 309111
rect 95433 309077 95467 309111
rect 95467 309077 95476 309111
rect 95424 309068 95476 309077
rect 124496 307844 124548 307896
rect 86040 307708 86092 307760
rect 124404 307708 124456 307760
rect 136640 307028 136692 307080
rect 137928 307028 137980 307080
rect 139400 307028 139452 307080
rect 140688 307028 140740 307080
rect 140872 307028 140924 307080
rect 142068 307028 142120 307080
rect 143632 307028 143684 307080
rect 144828 307028 144880 307080
rect 75000 302379 75052 302388
rect 75000 302345 75009 302379
rect 75009 302345 75043 302379
rect 75043 302345 75052 302379
rect 75000 302336 75052 302345
rect 134984 302243 135036 302252
rect 134984 302209 134993 302243
rect 134993 302209 135027 302243
rect 135027 302209 135036 302243
rect 134984 302200 135036 302209
rect 80428 301520 80480 301572
rect 66812 299523 66864 299532
rect 66812 299489 66821 299523
rect 66821 299489 66855 299523
rect 66855 299489 66864 299523
rect 66812 299480 66864 299489
rect 74448 299523 74500 299532
rect 74448 299489 74457 299523
rect 74457 299489 74491 299523
rect 74491 299489 74500 299523
rect 74448 299480 74500 299489
rect 75000 299523 75052 299532
rect 75000 299489 75009 299523
rect 75009 299489 75043 299523
rect 75043 299489 75052 299523
rect 75000 299480 75052 299489
rect 77576 299523 77628 299532
rect 77576 299489 77585 299523
rect 77585 299489 77619 299523
rect 77619 299489 77628 299523
rect 77576 299480 77628 299489
rect 95700 299480 95752 299532
rect 134984 299523 135036 299532
rect 134984 299489 134993 299523
rect 134993 299489 135027 299523
rect 135027 299489 135036 299523
rect 134984 299480 135036 299489
rect 75000 299344 75052 299396
rect 124220 298231 124272 298240
rect 124220 298197 124229 298231
rect 124229 298197 124263 298231
rect 124263 298197 124272 298231
rect 124220 298188 124272 298197
rect 85948 298163 86000 298172
rect 85948 298129 85957 298163
rect 85957 298129 85991 298163
rect 85991 298129 86000 298163
rect 85948 298120 86000 298129
rect 74448 298095 74500 298104
rect 74448 298061 74457 298095
rect 74457 298061 74491 298095
rect 74491 298061 74500 298095
rect 74448 298052 74500 298061
rect 124220 298052 124272 298104
rect 80244 296735 80296 296744
rect 80244 296701 80253 296735
rect 80253 296701 80287 296735
rect 80287 296701 80296 296735
rect 80244 296692 80296 296701
rect 140780 296692 140832 296744
rect 140964 296692 141016 296744
rect 66628 294584 66680 294636
rect 66812 294584 66864 294636
rect 72332 292612 72384 292664
rect 85948 292612 86000 292664
rect 85948 292476 86000 292528
rect 124404 292451 124456 292460
rect 124404 292417 124413 292451
rect 124413 292417 124447 292451
rect 124447 292417 124456 292451
rect 124404 292408 124456 292417
rect 72240 289867 72292 289876
rect 72240 289833 72249 289867
rect 72249 289833 72283 289867
rect 72283 289833 72292 289867
rect 72240 289824 72292 289833
rect 74908 289867 74960 289876
rect 74908 289833 74917 289867
rect 74917 289833 74951 289867
rect 74951 289833 74960 289867
rect 74908 289824 74960 289833
rect 135168 289756 135220 289808
rect 74908 289731 74960 289740
rect 74908 289697 74917 289731
rect 74917 289697 74951 289731
rect 74951 289697 74960 289731
rect 74908 289688 74960 289697
rect 80244 288260 80296 288312
rect 80428 288192 80480 288244
rect 81716 283611 81768 283620
rect 81716 283577 81725 283611
rect 81725 283577 81759 283611
rect 81759 283577 81768 283611
rect 81716 283568 81768 283577
rect 124404 282956 124456 283008
rect 77576 282931 77628 282940
rect 77576 282897 77585 282931
rect 77585 282897 77619 282931
rect 77619 282897 77628 282931
rect 77576 282888 77628 282897
rect 150164 282888 150216 282940
rect 150348 282888 150400 282940
rect 124404 282820 124456 282872
rect 74448 280211 74500 280220
rect 74448 280177 74457 280211
rect 74457 280177 74491 280211
rect 74491 280177 74500 280211
rect 74448 280168 74500 280177
rect 75000 280168 75052 280220
rect 134892 280211 134944 280220
rect 134892 280177 134901 280211
rect 134901 280177 134935 280211
rect 134935 280177 134944 280211
rect 134892 280168 134944 280177
rect 66536 280143 66588 280152
rect 66536 280109 66545 280143
rect 66545 280109 66579 280143
rect 66579 280109 66588 280143
rect 66536 280100 66588 280109
rect 72240 280143 72292 280152
rect 72240 280109 72249 280143
rect 72249 280109 72283 280143
rect 72283 280109 72292 280143
rect 72240 280100 72292 280109
rect 95608 280143 95660 280152
rect 95608 280109 95617 280143
rect 95617 280109 95651 280143
rect 95651 280109 95660 280143
rect 95608 280100 95660 280109
rect 124404 280143 124456 280152
rect 124404 280109 124413 280143
rect 124413 280109 124447 280143
rect 124447 280109 124456 280143
rect 124404 280100 124456 280109
rect 85856 278808 85908 278860
rect 85948 278808 86000 278860
rect 81716 278783 81768 278792
rect 81716 278749 81725 278783
rect 81725 278749 81759 278783
rect 81759 278749 81768 278783
rect 81716 278740 81768 278749
rect 85856 278672 85908 278724
rect 86040 278672 86092 278724
rect 86040 277312 86092 277364
rect 86132 277312 86184 277364
rect 124404 273955 124456 273964
rect 124404 273921 124413 273955
rect 124413 273921 124447 273955
rect 124447 273921 124456 273955
rect 124404 273912 124456 273921
rect 66628 270512 66680 270564
rect 72240 270555 72292 270564
rect 72240 270521 72249 270555
rect 72249 270521 72283 270555
rect 72283 270521 72292 270555
rect 72240 270512 72292 270521
rect 77576 270555 77628 270564
rect 77576 270521 77585 270555
rect 77585 270521 77619 270555
rect 77619 270521 77628 270555
rect 77576 270512 77628 270521
rect 95700 270512 95752 270564
rect 134984 270444 135036 270496
rect 74264 269084 74316 269136
rect 74448 269084 74500 269136
rect 124312 263619 124364 263628
rect 124312 263585 124321 263619
rect 124321 263585 124355 263619
rect 124355 263585 124364 263619
rect 124312 263576 124364 263585
rect 140780 263576 140832 263628
rect 140964 263576 141016 263628
rect 150164 263576 150216 263628
rect 150348 263576 150400 263628
rect 134892 260899 134944 260908
rect 134892 260865 134901 260899
rect 134901 260865 134935 260899
rect 134935 260865 134944 260899
rect 134892 260856 134944 260865
rect 66536 260831 66588 260840
rect 66536 260797 66545 260831
rect 66545 260797 66579 260831
rect 66579 260797 66588 260831
rect 66536 260788 66588 260797
rect 72240 260831 72292 260840
rect 72240 260797 72249 260831
rect 72249 260797 72283 260831
rect 72283 260797 72292 260831
rect 72240 260788 72292 260797
rect 75000 260831 75052 260840
rect 75000 260797 75009 260831
rect 75009 260797 75043 260831
rect 75043 260797 75052 260831
rect 75000 260788 75052 260797
rect 77576 260831 77628 260840
rect 77576 260797 77585 260831
rect 77585 260797 77619 260831
rect 77619 260797 77628 260831
rect 77576 260788 77628 260797
rect 80336 260788 80388 260840
rect 80428 260788 80480 260840
rect 95608 260831 95660 260840
rect 95608 260797 95617 260831
rect 95617 260797 95651 260831
rect 95651 260797 95660 260831
rect 95608 260788 95660 260797
rect 124312 259471 124364 259480
rect 124312 259437 124321 259471
rect 124321 259437 124355 259471
rect 124355 259437 124364 259471
rect 124312 259428 124364 259437
rect 124312 253920 124364 253972
rect 124404 253784 124456 253836
rect 66628 251200 66680 251252
rect 72240 251243 72292 251252
rect 72240 251209 72249 251243
rect 72249 251209 72283 251243
rect 72283 251209 72292 251243
rect 72240 251200 72292 251209
rect 75000 251243 75052 251252
rect 75000 251209 75009 251243
rect 75009 251209 75043 251243
rect 75043 251209 75052 251243
rect 75000 251200 75052 251209
rect 77576 251243 77628 251252
rect 77576 251209 77585 251243
rect 77585 251209 77619 251243
rect 77619 251209 77628 251243
rect 77576 251200 77628 251209
rect 81808 251200 81860 251252
rect 81900 251200 81952 251252
rect 95700 251200 95752 251252
rect 85948 251132 86000 251184
rect 86132 251132 86184 251184
rect 134984 251132 135036 251184
rect 74264 249772 74316 249824
rect 74448 249772 74500 249824
rect 124404 244332 124456 244384
rect 140780 244264 140832 244316
rect 140964 244264 141016 244316
rect 150164 244264 150216 244316
rect 150348 244264 150400 244316
rect 124312 244196 124364 244248
rect 134892 241519 134944 241528
rect 134892 241485 134901 241519
rect 134901 241485 134935 241519
rect 134935 241485 134944 241519
rect 134892 241476 134944 241485
rect 77668 234608 77720 234660
rect 85948 234608 86000 234660
rect 124312 234608 124364 234660
rect 134892 234608 134944 234660
rect 77576 234540 77628 234592
rect 85856 234540 85908 234592
rect 124404 234472 124456 234524
rect 134984 234472 135036 234524
rect 66352 231820 66404 231872
rect 66628 231820 66680 231872
rect 72056 231820 72108 231872
rect 72240 231820 72292 231872
rect 74816 231820 74868 231872
rect 75000 231820 75052 231872
rect 80336 231820 80388 231872
rect 80428 231820 80480 231872
rect 81808 231820 81860 231872
rect 81900 231820 81952 231872
rect 95424 231820 95476 231872
rect 95700 231820 95752 231872
rect 74264 230460 74316 230512
rect 74448 230460 74500 230512
rect 124312 224995 124364 225004
rect 124312 224961 124321 224995
rect 124321 224961 124355 224995
rect 124355 224961 124364 224995
rect 124312 224952 124364 224961
rect 134892 224995 134944 225004
rect 134892 224961 134901 224995
rect 134901 224961 134935 224995
rect 134935 224961 134944 224995
rect 134892 224952 134944 224961
rect 140780 224952 140832 225004
rect 140964 224952 141016 225004
rect 150164 224952 150216 225004
rect 150348 224952 150400 225004
rect 124312 222207 124364 222216
rect 124312 222173 124321 222207
rect 124321 222173 124355 222207
rect 124355 222173 124364 222207
rect 124312 222164 124364 222173
rect 134892 222207 134944 222216
rect 134892 222173 134901 222207
rect 134901 222173 134935 222207
rect 134935 222173 134944 222207
rect 134892 222164 134944 222173
rect 124312 215296 124364 215348
rect 134892 215296 134944 215348
rect 124404 215160 124456 215212
rect 134984 215160 135036 215212
rect 66352 212508 66404 212560
rect 66628 212508 66680 212560
rect 72056 212508 72108 212560
rect 72240 212508 72292 212560
rect 74816 212508 74868 212560
rect 75000 212508 75052 212560
rect 77576 212508 77628 212560
rect 77760 212508 77812 212560
rect 80336 212508 80388 212560
rect 80428 212508 80480 212560
rect 81808 212508 81860 212560
rect 81900 212508 81952 212560
rect 95424 212508 95476 212560
rect 95700 212508 95752 212560
rect 124312 205683 124364 205692
rect 124312 205649 124321 205683
rect 124321 205649 124355 205683
rect 124355 205649 124364 205683
rect 124312 205640 124364 205649
rect 134892 205683 134944 205692
rect 134892 205649 134901 205683
rect 134901 205649 134935 205683
rect 134935 205649 134944 205683
rect 134892 205640 134944 205649
rect 140780 205640 140832 205692
rect 140964 205640 141016 205692
rect 150164 205640 150216 205692
rect 150348 205640 150400 205692
rect 85948 202852 86000 202904
rect 86132 202852 86184 202904
rect 124312 202895 124364 202904
rect 124312 202861 124321 202895
rect 124321 202861 124355 202895
rect 124355 202861 124364 202895
rect 124312 202852 124364 202861
rect 134892 202895 134944 202904
rect 134892 202861 134901 202895
rect 134901 202861 134935 202895
rect 134935 202861 134944 202895
rect 134892 202852 134944 202861
rect 80336 202784 80388 202836
rect 80428 202784 80480 202836
rect 74264 201424 74316 201476
rect 74448 201424 74500 201476
rect 77668 195984 77720 196036
rect 85948 195984 86000 196036
rect 124312 195984 124364 196036
rect 134892 195984 134944 196036
rect 77576 195916 77628 195968
rect 85856 195916 85908 195968
rect 124404 195848 124456 195900
rect 134984 195848 135036 195900
rect 66352 193196 66404 193248
rect 66628 193196 66680 193248
rect 72056 193196 72108 193248
rect 72240 193196 72292 193248
rect 74816 193196 74868 193248
rect 75000 193196 75052 193248
rect 81808 193196 81860 193248
rect 81900 193196 81952 193248
rect 95424 193196 95476 193248
rect 95700 193196 95752 193248
rect 160560 193196 160612 193248
rect 160744 193196 160796 193248
rect 124312 186371 124364 186380
rect 124312 186337 124321 186371
rect 124321 186337 124355 186371
rect 124355 186337 124364 186371
rect 124312 186328 124364 186337
rect 140780 186328 140832 186380
rect 140964 186328 141016 186380
rect 150164 186328 150216 186380
rect 150348 186328 150400 186380
rect 85948 183540 86000 183592
rect 86132 183540 86184 183592
rect 124312 183583 124364 183592
rect 124312 183549 124321 183583
rect 124321 183549 124355 183583
rect 124355 183549 124364 183583
rect 124312 183540 124364 183549
rect 134800 183540 134852 183592
rect 135076 183540 135128 183592
rect 80336 183472 80388 183524
rect 80428 183472 80480 183524
rect 74264 182112 74316 182164
rect 74448 182112 74500 182164
rect 135076 176740 135128 176792
rect 77484 176672 77536 176724
rect 85948 176672 86000 176724
rect 124312 176672 124364 176724
rect 77576 176604 77628 176656
rect 85856 176604 85908 176656
rect 124404 176536 124456 176588
rect 134984 176536 135036 176588
rect 66352 173884 66404 173936
rect 66628 173884 66680 173936
rect 72056 173884 72108 173936
rect 72240 173884 72292 173936
rect 74816 173884 74868 173936
rect 75000 173884 75052 173936
rect 81808 173884 81860 173936
rect 81900 173884 81952 173936
rect 95424 173884 95476 173936
rect 95700 173884 95752 173936
rect 140964 173884 141016 173936
rect 141148 173884 141200 173936
rect 150072 173884 150124 173936
rect 150348 173884 150400 173936
rect 124312 167059 124364 167068
rect 124312 167025 124321 167059
rect 124321 167025 124355 167059
rect 124355 167025 124364 167059
rect 124312 167016 124364 167025
rect 140780 167016 140832 167068
rect 140964 167016 141016 167068
rect 150164 167016 150216 167068
rect 150348 167016 150400 167068
rect 78864 166948 78916 167000
rect 134800 166948 134852 167000
rect 134984 166948 135036 167000
rect 78864 166812 78916 166864
rect 124312 164271 124364 164280
rect 124312 164237 124321 164271
rect 124321 164237 124355 164271
rect 124355 164237 124364 164271
rect 124312 164228 124364 164237
rect 66352 164160 66404 164212
rect 66536 164160 66588 164212
rect 95424 164160 95476 164212
rect 95608 164160 95660 164212
rect 140872 164203 140924 164212
rect 140872 164169 140881 164203
rect 140881 164169 140915 164203
rect 140915 164169 140924 164203
rect 140872 164160 140924 164169
rect 150256 164203 150308 164212
rect 150256 164169 150265 164203
rect 150265 164169 150299 164203
rect 150299 164169 150308 164203
rect 150256 164160 150308 164169
rect 74448 162843 74500 162852
rect 74448 162809 74457 162843
rect 74457 162809 74491 162843
rect 74491 162809 74500 162843
rect 74448 162800 74500 162809
rect 78864 162843 78916 162852
rect 78864 162809 78873 162843
rect 78873 162809 78907 162843
rect 78907 162809 78916 162843
rect 78864 162800 78916 162809
rect 135076 157471 135128 157480
rect 135076 157437 135085 157471
rect 135085 157437 135119 157471
rect 135119 157437 135128 157471
rect 135076 157428 135128 157437
rect 124312 157360 124364 157412
rect 80244 157292 80296 157344
rect 80428 157292 80480 157344
rect 81716 157292 81768 157344
rect 81900 157292 81952 157344
rect 85856 157292 85908 157344
rect 86040 157292 86092 157344
rect 140872 157335 140924 157344
rect 140872 157301 140881 157335
rect 140881 157301 140915 157335
rect 140915 157301 140924 157335
rect 140872 157292 140924 157301
rect 150256 157335 150308 157344
rect 150256 157301 150265 157335
rect 150265 157301 150299 157335
rect 150299 157301 150308 157335
rect 150256 157292 150308 157301
rect 124404 157224 124456 157276
rect 135076 154615 135128 154624
rect 135076 154581 135085 154615
rect 135085 154581 135119 154615
rect 135119 154581 135128 154615
rect 135076 154572 135128 154581
rect 80336 154504 80388 154556
rect 80428 154504 80480 154556
rect 81808 154504 81860 154556
rect 81900 154504 81952 154556
rect 124404 154504 124456 154556
rect 124588 154504 124640 154556
rect 74448 153255 74500 153264
rect 74448 153221 74457 153255
rect 74457 153221 74491 153255
rect 74491 153221 74500 153255
rect 74448 153212 74500 153221
rect 78864 153255 78916 153264
rect 78864 153221 78873 153255
rect 78873 153221 78907 153255
rect 78907 153221 78916 153255
rect 78864 153212 78916 153221
rect 135076 147679 135128 147688
rect 135076 147645 135085 147679
rect 135085 147645 135119 147679
rect 135119 147645 135128 147679
rect 135076 147636 135128 147645
rect 140780 147636 140832 147688
rect 140964 147636 141016 147688
rect 150164 147636 150216 147688
rect 150348 147636 150400 147688
rect 135076 144959 135128 144968
rect 135076 144925 135085 144959
rect 135085 144925 135119 144959
rect 135119 144925 135128 144959
rect 135076 144916 135128 144925
rect 85856 144848 85908 144900
rect 85948 144848 86000 144900
rect 140872 144891 140924 144900
rect 140872 144857 140881 144891
rect 140881 144857 140915 144891
rect 140915 144857 140924 144891
rect 140872 144848 140924 144857
rect 150256 144891 150308 144900
rect 150256 144857 150265 144891
rect 150265 144857 150299 144891
rect 150299 144857 150308 144891
rect 150256 144848 150308 144857
rect 74448 143531 74500 143540
rect 74448 143497 74457 143531
rect 74457 143497 74491 143531
rect 74491 143497 74500 143531
rect 74448 143488 74500 143497
rect 75000 143531 75052 143540
rect 75000 143497 75009 143531
rect 75009 143497 75043 143531
rect 75043 143497 75052 143531
rect 75000 143488 75052 143497
rect 78772 140020 78824 140072
rect 78864 139952 78916 140004
rect 80336 137980 80388 138032
rect 81808 137980 81860 138032
rect 124312 137980 124364 138032
rect 80428 137912 80480 137964
rect 81900 137912 81952 137964
rect 135076 138048 135128 138100
rect 124404 137912 124456 137964
rect 134984 137912 135036 137964
rect 140872 137955 140924 137964
rect 140872 137921 140881 137955
rect 140881 137921 140915 137955
rect 140915 137921 140924 137955
rect 140872 137912 140924 137921
rect 150256 137955 150308 137964
rect 150256 137921 150265 137955
rect 150265 137921 150299 137955
rect 150299 137921 150308 137955
rect 150256 137912 150308 137921
rect 77576 135328 77628 135380
rect 77576 135192 77628 135244
rect 124404 135192 124456 135244
rect 124588 135192 124640 135244
rect 74448 133943 74500 133952
rect 74448 133909 74457 133943
rect 74457 133909 74491 133943
rect 74491 133909 74500 133943
rect 74448 133900 74500 133909
rect 75000 133943 75052 133952
rect 75000 133909 75009 133943
rect 75009 133909 75043 133943
rect 75043 133909 75052 133943
rect 75000 133900 75052 133909
rect 77668 133832 77720 133884
rect 77852 133832 77904 133884
rect 134984 128324 135036 128376
rect 140780 128324 140832 128376
rect 140964 128324 141016 128376
rect 150164 128324 150216 128376
rect 150348 128324 150400 128376
rect 135076 128256 135128 128308
rect 78772 125536 78824 125588
rect 85856 125536 85908 125588
rect 85948 125536 86000 125588
rect 140872 125579 140924 125588
rect 140872 125545 140881 125579
rect 140881 125545 140915 125579
rect 140915 125545 140924 125579
rect 140872 125536 140924 125545
rect 150256 125579 150308 125588
rect 150256 125545 150265 125579
rect 150265 125545 150299 125579
rect 150299 125545 150308 125579
rect 150256 125536 150308 125545
rect 78864 125400 78916 125452
rect 77484 124108 77536 124160
rect 77576 124108 77628 124160
rect 135076 124108 135128 124160
rect 72240 122791 72292 122800
rect 72240 122757 72249 122791
rect 72249 122757 72283 122791
rect 72283 122757 72292 122791
rect 72240 122748 72292 122757
rect 75000 122791 75052 122800
rect 75000 122757 75009 122791
rect 75009 122757 75043 122791
rect 75043 122757 75052 122791
rect 75000 122748 75052 122757
rect 80336 118668 80388 118720
rect 81808 118668 81860 118720
rect 124312 118668 124364 118720
rect 80428 118600 80480 118652
rect 81900 118600 81952 118652
rect 124404 118600 124456 118652
rect 140872 118643 140924 118652
rect 140872 118609 140881 118643
rect 140881 118609 140915 118643
rect 140915 118609 140924 118643
rect 140872 118600 140924 118609
rect 150256 118643 150308 118652
rect 150256 118609 150265 118643
rect 150265 118609 150299 118643
rect 150299 118609 150308 118643
rect 150256 118600 150308 118609
rect 75000 117283 75052 117292
rect 75000 117249 75009 117283
rect 75009 117249 75043 117283
rect 75043 117249 75052 117283
rect 75000 117240 75052 117249
rect 124404 115880 124456 115932
rect 124588 115880 124640 115932
rect 134984 114563 135036 114572
rect 134984 114529 134993 114563
rect 134993 114529 135027 114563
rect 135027 114529 135036 114563
rect 134984 114520 135036 114529
rect 77576 114495 77628 114504
rect 77576 114461 77585 114495
rect 77585 114461 77619 114495
rect 77619 114461 77628 114495
rect 77576 114452 77628 114461
rect 72240 113203 72292 113212
rect 72240 113169 72249 113203
rect 72249 113169 72283 113203
rect 72283 113169 72292 113203
rect 72240 113160 72292 113169
rect 134984 109012 135036 109064
rect 140780 109012 140832 109064
rect 140964 109012 141016 109064
rect 150164 109012 150216 109064
rect 150348 109012 150400 109064
rect 135076 108944 135128 108996
rect 85948 106292 86000 106344
rect 86040 106292 86092 106344
rect 140872 106267 140924 106276
rect 140872 106233 140881 106267
rect 140881 106233 140915 106267
rect 140915 106233 140924 106267
rect 140872 106224 140924 106233
rect 150256 106267 150308 106276
rect 150256 106233 150265 106267
rect 150265 106233 150299 106267
rect 150299 106233 150308 106267
rect 150256 106224 150308 106233
rect 77576 104907 77628 104916
rect 77576 104873 77585 104907
rect 77585 104873 77619 104907
rect 77619 104873 77628 104907
rect 77576 104864 77628 104873
rect 74448 104839 74500 104848
rect 74448 104805 74457 104839
rect 74457 104805 74491 104839
rect 74491 104805 74500 104839
rect 74448 104796 74500 104805
rect 78772 104839 78824 104848
rect 78772 104805 78781 104839
rect 78781 104805 78815 104839
rect 78815 104805 78824 104839
rect 78772 104796 78824 104805
rect 85948 104839 86000 104848
rect 85948 104805 85957 104839
rect 85957 104805 85991 104839
rect 85991 104805 86000 104839
rect 85948 104796 86000 104805
rect 135076 104796 135128 104848
rect 72332 102076 72384 102128
rect 124312 99356 124364 99408
rect 124404 99288 124456 99340
rect 140872 99331 140924 99340
rect 140872 99297 140881 99331
rect 140881 99297 140915 99331
rect 140915 99297 140924 99331
rect 140872 99288 140924 99297
rect 150256 99331 150308 99340
rect 150256 99297 150265 99331
rect 150265 99297 150299 99331
rect 150299 99297 150308 99331
rect 150256 99288 150308 99297
rect 124404 96568 124456 96620
rect 124588 96568 124640 96620
rect 74448 95251 74500 95260
rect 74448 95217 74457 95251
rect 74457 95217 74491 95251
rect 74491 95217 74500 95251
rect 74448 95208 74500 95217
rect 78956 95208 79008 95260
rect 86040 95208 86092 95260
rect 75000 93823 75052 93832
rect 75000 93789 75009 93823
rect 75009 93789 75043 93823
rect 75043 93789 75052 93823
rect 75000 93780 75052 93789
rect 72240 92531 72292 92540
rect 72240 92497 72249 92531
rect 72249 92497 72283 92531
rect 72283 92497 72292 92531
rect 72240 92488 72292 92497
rect 140780 89700 140832 89752
rect 140964 89700 141016 89752
rect 150164 89700 150216 89752
rect 150348 89700 150400 89752
rect 134984 89675 135036 89684
rect 134984 89641 134993 89675
rect 134993 89641 135027 89675
rect 135027 89641 135036 89675
rect 134984 89632 135036 89641
rect 66444 86912 66496 86964
rect 85948 86912 86000 86964
rect 95516 86912 95568 86964
rect 140872 86955 140924 86964
rect 140872 86921 140881 86955
rect 140881 86921 140915 86955
rect 140915 86921 140924 86955
rect 140872 86912 140924 86921
rect 150256 86955 150308 86964
rect 150256 86921 150265 86955
rect 150265 86921 150299 86955
rect 150299 86921 150308 86955
rect 150256 86912 150308 86921
rect 160744 86887 160796 86896
rect 160744 86853 160753 86887
rect 160753 86853 160787 86887
rect 160787 86853 160796 86887
rect 160744 86844 160796 86853
rect 78772 85552 78824 85604
rect 78956 85552 79008 85604
rect 75000 84303 75052 84312
rect 75000 84269 75009 84303
rect 75009 84269 75043 84303
rect 75043 84269 75052 84303
rect 75000 84260 75052 84269
rect 75000 84167 75052 84176
rect 75000 84133 75009 84167
rect 75009 84133 75043 84167
rect 75043 84133 75052 84167
rect 75000 84124 75052 84133
rect 134708 82084 134760 82136
rect 135076 82084 135128 82136
rect 81716 80112 81768 80164
rect 124312 80044 124364 80096
rect 81624 79976 81676 80028
rect 124404 79908 124456 79960
rect 66352 77299 66404 77308
rect 66352 77265 66361 77299
rect 66361 77265 66395 77299
rect 66395 77265 66404 77299
rect 66352 77256 66404 77265
rect 85856 77299 85908 77308
rect 85856 77265 85865 77299
rect 85865 77265 85899 77299
rect 85899 77265 85908 77299
rect 85856 77256 85908 77265
rect 95424 77299 95476 77308
rect 95424 77265 95433 77299
rect 95433 77265 95467 77299
rect 95467 77265 95476 77299
rect 95424 77256 95476 77265
rect 140964 77256 141016 77308
rect 150348 77256 150400 77308
rect 160744 77299 160796 77308
rect 160744 77265 160753 77299
rect 160753 77265 160787 77299
rect 160787 77265 160796 77299
rect 160744 77256 160796 77265
rect 81624 77231 81676 77240
rect 81624 77197 81633 77231
rect 81633 77197 81667 77231
rect 81667 77197 81676 77231
rect 81624 77188 81676 77197
rect 66352 77163 66404 77172
rect 66352 77129 66361 77163
rect 66361 77129 66395 77163
rect 66395 77129 66404 77163
rect 66352 77120 66404 77129
rect 95424 77163 95476 77172
rect 95424 77129 95433 77163
rect 95433 77129 95467 77163
rect 95467 77129 95476 77163
rect 95424 77120 95476 77129
rect 140964 77120 141016 77172
rect 78772 75896 78824 75948
rect 78864 75896 78916 75948
rect 75000 74579 75052 74588
rect 75000 74545 75009 74579
rect 75009 74545 75043 74579
rect 75043 74545 75052 74579
rect 75000 74536 75052 74545
rect 75000 71068 75052 71120
rect 80336 70388 80388 70440
rect 134984 70456 135036 70508
rect 150164 70388 150216 70440
rect 134892 70320 134944 70372
rect 150256 70320 150308 70372
rect 66444 70252 66496 70304
rect 80336 70252 80388 70304
rect 81716 70252 81768 70304
rect 95516 70252 95568 70304
rect 77576 67668 77628 67720
rect 77484 67600 77536 67652
rect 140872 67643 140924 67652
rect 140872 67609 140881 67643
rect 140881 67609 140915 67643
rect 140915 67609 140924 67643
rect 140872 67600 140924 67609
rect 74816 66283 74868 66292
rect 74816 66249 74825 66283
rect 74825 66249 74859 66283
rect 74859 66249 74868 66283
rect 74816 66240 74868 66249
rect 124404 66240 124456 66292
rect 124588 66240 124640 66292
rect 72148 66172 72200 66224
rect 72424 66172 72476 66224
rect 74448 66215 74500 66224
rect 74448 66181 74457 66215
rect 74457 66181 74491 66215
rect 74491 66181 74500 66215
rect 74448 66172 74500 66181
rect 77484 66215 77536 66224
rect 77484 66181 77493 66215
rect 77493 66181 77527 66215
rect 77527 66181 77536 66215
rect 77484 66172 77536 66181
rect 134892 66172 134944 66224
rect 135076 66172 135128 66224
rect 72424 64855 72476 64864
rect 72424 64821 72433 64855
rect 72433 64821 72467 64855
rect 72467 64821 72476 64855
rect 72424 64812 72476 64821
rect 74816 64855 74868 64864
rect 74816 64821 74825 64855
rect 74825 64821 74859 64855
rect 74859 64821 74868 64855
rect 74816 64812 74868 64821
rect 66444 60664 66496 60716
rect 66628 60664 66680 60716
rect 80244 60664 80296 60716
rect 80428 60664 80480 60716
rect 81716 60664 81768 60716
rect 81900 60664 81952 60716
rect 95516 60664 95568 60716
rect 95700 60664 95752 60716
rect 124404 60596 124456 60648
rect 124588 60596 124640 60648
rect 66628 57876 66680 57928
rect 95700 57876 95752 57928
rect 140964 57876 141016 57928
rect 150348 57876 150400 57928
rect 74448 56627 74500 56636
rect 74448 56593 74457 56627
rect 74457 56593 74491 56627
rect 74491 56593 74500 56627
rect 74448 56584 74500 56593
rect 72424 56559 72476 56568
rect 72424 56525 72433 56559
rect 72433 56525 72467 56559
rect 72467 56525 72476 56559
rect 72424 56516 72476 56525
rect 124404 56559 124456 56568
rect 124404 56525 124413 56559
rect 124413 56525 124447 56559
rect 124447 56525 124456 56559
rect 124404 56516 124456 56525
rect 74908 55224 74960 55276
rect 72424 55156 72476 55208
rect 140872 51051 140924 51060
rect 140872 51017 140881 51051
rect 140881 51017 140915 51051
rect 140915 51017 140924 51051
rect 140872 51008 140924 51017
rect 77484 48399 77536 48408
rect 77484 48365 77493 48399
rect 77493 48365 77527 48399
rect 77527 48365 77536 48399
rect 77484 48356 77536 48365
rect 66536 48331 66588 48340
rect 66536 48297 66545 48331
rect 66545 48297 66579 48331
rect 66579 48297 66588 48331
rect 66536 48288 66588 48297
rect 95608 48331 95660 48340
rect 95608 48297 95617 48331
rect 95617 48297 95651 48331
rect 95651 48297 95660 48331
rect 95608 48288 95660 48297
rect 150256 48331 150308 48340
rect 150256 48297 150265 48331
rect 150265 48297 150299 48331
rect 150299 48297 150308 48331
rect 150256 48288 150308 48297
rect 124496 46928 124548 46980
rect 74448 46903 74500 46912
rect 74448 46869 74457 46903
rect 74457 46869 74491 46903
rect 74491 46869 74500 46903
rect 74448 46860 74500 46869
rect 74908 46860 74960 46912
rect 75092 46860 75144 46912
rect 77484 46860 77536 46912
rect 77760 46860 77812 46912
rect 134892 46860 134944 46912
rect 135076 46860 135128 46912
rect 72332 45679 72384 45688
rect 72332 45645 72341 45679
rect 72341 45645 72375 45679
rect 72375 45645 72384 45679
rect 72332 45636 72384 45645
rect 72332 45543 72384 45552
rect 72332 45509 72341 45543
rect 72341 45509 72375 45543
rect 72375 45509 72384 45543
rect 72332 45500 72384 45509
rect 75092 45500 75144 45552
rect 66444 41352 66496 41404
rect 66628 41352 66680 41404
rect 80244 41352 80296 41404
rect 80428 41352 80480 41404
rect 81716 41352 81768 41404
rect 81900 41352 81952 41404
rect 95516 41352 95568 41404
rect 95700 41352 95752 41404
rect 66628 38564 66680 38616
rect 78864 38607 78916 38616
rect 78864 38573 78873 38607
rect 78873 38573 78907 38607
rect 78907 38573 78916 38607
rect 78864 38564 78916 38573
rect 95700 38564 95752 38616
rect 140964 38564 141016 38616
rect 150348 38564 150400 38616
rect 74448 37315 74500 37324
rect 74448 37281 74457 37315
rect 74457 37281 74491 37315
rect 74491 37281 74500 37315
rect 74448 37272 74500 37281
rect 75092 37204 75144 37256
rect 72148 31696 72200 31748
rect 140872 31739 140924 31748
rect 140872 31705 140881 31739
rect 140881 31705 140915 31739
rect 140915 31705 140924 31739
rect 140872 31696 140924 31705
rect 74816 29724 74868 29776
rect 75092 29724 75144 29776
rect 66536 29019 66588 29028
rect 66536 28985 66545 29019
rect 66545 28985 66579 29019
rect 66579 28985 66588 29019
rect 66536 28976 66588 28985
rect 78864 29019 78916 29028
rect 78864 28985 78873 29019
rect 78873 28985 78907 29019
rect 78907 28985 78916 29019
rect 78864 28976 78916 28985
rect 81808 28976 81860 29028
rect 81900 28976 81952 29028
rect 85856 28976 85908 29028
rect 95608 29019 95660 29028
rect 95608 28985 95617 29019
rect 95617 28985 95651 29019
rect 95651 28985 95660 29019
rect 95608 28976 95660 28985
rect 150256 29019 150308 29028
rect 150256 28985 150265 29019
rect 150265 28985 150299 29019
rect 150299 28985 150308 29019
rect 150256 28976 150308 28985
rect 77208 28840 77260 28892
rect 77760 28840 77812 28892
rect 85948 28840 86000 28892
rect 124404 27616 124456 27668
rect 124588 27616 124640 27668
rect 72148 27548 72200 27600
rect 74448 27548 74500 27600
rect 74816 27548 74868 27600
rect 134892 27591 134944 27600
rect 134892 27557 134901 27591
rect 134901 27557 134935 27591
rect 134935 27557 134944 27591
rect 134892 27548 134944 27557
rect 72332 27480 72384 27532
rect 85948 26188 86000 26240
rect 86040 26188 86092 26240
rect 66444 22040 66496 22092
rect 66628 22040 66680 22092
rect 80244 22040 80296 22092
rect 80428 22040 80480 22092
rect 81716 22040 81768 22092
rect 81900 22040 81952 22092
rect 95516 22040 95568 22092
rect 95700 22040 95752 22092
rect 160652 19320 160704 19372
rect 160744 19320 160796 19372
rect 66628 19295 66680 19304
rect 66628 19261 66637 19295
rect 66637 19261 66671 19295
rect 66671 19261 66680 19295
rect 66628 19252 66680 19261
rect 95700 19295 95752 19304
rect 95700 19261 95709 19295
rect 95709 19261 95743 19295
rect 95743 19261 95752 19295
rect 95700 19252 95752 19261
rect 77208 19184 77260 19236
rect 77760 19184 77812 19236
rect 124404 17960 124456 18012
rect 124588 17960 124640 18012
rect 134984 17960 135036 18012
rect 244004 16532 244056 16584
rect 485780 16532 485832 16584
rect 245384 16464 245436 16516
rect 489920 16464 489972 16516
rect 246856 16396 246908 16448
rect 494060 16396 494112 16448
rect 246764 16328 246816 16380
rect 494152 16328 494204 16380
rect 248144 16260 248196 16312
rect 496820 16260 496872 16312
rect 249524 16192 249576 16244
rect 500960 16192 501012 16244
rect 250904 16124 250956 16176
rect 503720 16124 503772 16176
rect 252284 16056 252336 16108
rect 507860 16056 507912 16108
rect 274364 15988 274416 16040
rect 567200 15988 567252 16040
rect 277124 15920 277176 15972
rect 574100 15920 574152 15972
rect 278504 15852 278556 15904
rect 578240 15852 578292 15904
rect 242532 15784 242584 15836
rect 483020 15784 483072 15836
rect 227444 15716 227496 15768
rect 443000 15716 443052 15768
rect 219164 15648 219216 15700
rect 420920 15648 420972 15700
rect 213644 15580 213696 15632
rect 407120 15580 407172 15632
rect 180524 15512 180576 15564
rect 317420 15512 317472 15564
rect 215024 15104 215076 15156
rect 408500 15104 408552 15156
rect 223304 15036 223356 15088
rect 431960 15036 432012 15088
rect 226064 14968 226116 15020
rect 438860 14968 438912 15020
rect 228824 14900 228876 14952
rect 445760 14900 445812 14952
rect 231584 14832 231636 14884
rect 452660 14832 452712 14884
rect 234344 14764 234396 14816
rect 459560 14764 459612 14816
rect 237104 14696 237156 14748
rect 467840 14696 467892 14748
rect 239864 14628 239916 14680
rect 474740 14628 474792 14680
rect 242624 14560 242676 14612
rect 481640 14560 481692 14612
rect 244096 14492 244148 14544
rect 487160 14492 487212 14544
rect 245476 14424 245528 14476
rect 491300 14424 491352 14476
rect 213736 14356 213788 14408
rect 405740 14356 405792 14408
rect 212264 14288 212316 14340
rect 401600 14288 401652 14340
rect 208124 14220 208176 14272
rect 390560 14220 390612 14272
rect 176476 14152 176528 14204
rect 305000 14152 305052 14204
rect 175096 14084 175148 14136
rect 302240 14084 302292 14136
rect 173716 14016 173768 14068
rect 298100 14016 298152 14068
rect 170956 13948 171008 14000
rect 293960 13948 294012 14000
rect 172336 13880 172388 13932
rect 295340 13880 295392 13932
rect 168104 13812 168156 13864
rect 287060 13812 287112 13864
rect 212356 13744 212408 13796
rect 402980 13744 403032 13796
rect 216404 13676 216456 13728
rect 414020 13676 414072 13728
rect 220544 13608 220596 13660
rect 425060 13608 425112 13660
rect 256424 13540 256476 13592
rect 517520 13540 517572 13592
rect 257804 13472 257856 13524
rect 520280 13472 520332 13524
rect 259184 13404 259236 13456
rect 524420 13404 524472 13456
rect 260564 13336 260616 13388
rect 528560 13336 528612 13388
rect 261944 13268 261996 13320
rect 531320 13268 531372 13320
rect 261852 13200 261904 13252
rect 535460 13200 535512 13252
rect 263324 13132 263376 13184
rect 538220 13132 538272 13184
rect 124404 13064 124456 13116
rect 125324 13064 125376 13116
rect 264704 13064 264756 13116
rect 542360 13064 542412 13116
rect 208216 12996 208268 13048
rect 391940 12996 391992 13048
rect 205364 12928 205416 12980
rect 385040 12928 385092 12980
rect 203984 12860 204036 12912
rect 378140 12860 378192 12912
rect 202604 12792 202656 12844
rect 374000 12792 374052 12844
rect 201224 12724 201276 12776
rect 371240 12724 371292 12776
rect 198464 12656 198516 12708
rect 364340 12656 364392 12708
rect 195704 12588 195756 12640
rect 356060 12588 356112 12640
rect 192944 12520 192996 12572
rect 349160 12520 349212 12572
rect 134984 12452 135036 12504
rect 190184 12452 190236 12504
rect 342260 12452 342312 12504
rect 134892 12384 134944 12436
rect 160376 12384 160428 12436
rect 161112 12384 161164 12436
rect 228916 12384 228968 12436
rect 444380 12384 444432 12436
rect 230204 12316 230256 12368
rect 448520 12316 448572 12368
rect 231676 12248 231728 12300
rect 451280 12248 451332 12300
rect 232964 12180 233016 12232
rect 455420 12180 455472 12232
rect 234436 12112 234488 12164
rect 459652 12112 459704 12164
rect 235724 12044 235776 12096
rect 462320 12044 462372 12096
rect 237196 11976 237248 12028
rect 466460 11976 466512 12028
rect 238484 11908 238536 11960
rect 469220 11908 469272 11960
rect 239956 11840 240008 11892
rect 473360 11840 473412 11892
rect 241244 11772 241296 11824
rect 477500 11772 477552 11824
rect 242716 11704 242768 11756
rect 480260 11704 480312 11756
rect 227536 11636 227588 11688
rect 441620 11636 441672 11688
rect 226156 11568 226208 11620
rect 437480 11568 437532 11620
rect 224684 11500 224736 11552
rect 433340 11500 433392 11552
rect 223396 11432 223448 11484
rect 430580 11432 430632 11484
rect 221924 11364 221976 11416
rect 426440 11364 426492 11416
rect 220636 11296 220688 11348
rect 423680 11296 423732 11348
rect 219256 11228 219308 11280
rect 419540 11228 419592 11280
rect 217876 11160 217928 11212
rect 416872 11160 416924 11212
rect 216496 11092 216548 11144
rect 412640 11092 412692 11144
rect 188896 10956 188948 11008
rect 340880 10956 340932 11008
rect 190276 10888 190328 10940
rect 345020 10888 345072 10940
rect 191564 10820 191616 10872
rect 347780 10820 347832 10872
rect 193036 10752 193088 10804
rect 351920 10752 351972 10804
rect 194416 10684 194468 10736
rect 356152 10684 356204 10736
rect 195796 10616 195848 10668
rect 358820 10616 358872 10668
rect 197084 10548 197136 10600
rect 362960 10548 363012 10600
rect 198556 10480 198608 10532
rect 365720 10480 365772 10532
rect 199936 10412 199988 10464
rect 369860 10412 369912 10464
rect 201316 10344 201368 10396
rect 374092 10344 374144 10396
rect 202696 10276 202748 10328
rect 376760 10276 376812 10328
rect 187516 10208 187568 10260
rect 338120 10208 338172 10260
rect 187424 10140 187476 10192
rect 333980 10140 334032 10192
rect 186136 10072 186188 10124
rect 331312 10072 331364 10124
rect 184756 10004 184808 10056
rect 327080 10004 327132 10056
rect 183376 9936 183428 9988
rect 322940 9936 322992 9988
rect 181996 9868 182048 9920
rect 320180 9868 320232 9920
rect 180616 9800 180668 9852
rect 316040 9800 316092 9852
rect 179236 9732 179288 9784
rect 313280 9732 313332 9784
rect 66628 9707 66680 9716
rect 66628 9673 66637 9707
rect 66637 9673 66671 9707
rect 66671 9673 66680 9707
rect 66628 9664 66680 9673
rect 72056 9664 72108 9716
rect 72332 9664 72384 9716
rect 74264 9707 74316 9716
rect 74264 9673 74273 9707
rect 74273 9673 74307 9707
rect 74307 9673 74316 9707
rect 74264 9664 74316 9673
rect 74908 9707 74960 9716
rect 74908 9673 74917 9707
rect 74917 9673 74951 9707
rect 74951 9673 74960 9707
rect 74908 9664 74960 9673
rect 77484 9664 77536 9716
rect 77760 9664 77812 9716
rect 95700 9707 95752 9716
rect 95700 9673 95709 9707
rect 95709 9673 95743 9707
rect 95743 9673 95752 9707
rect 95700 9664 95752 9673
rect 177856 9664 177908 9716
rect 309140 9664 309192 9716
rect 140780 9596 140832 9648
rect 154304 9596 154356 9648
rect 249156 9596 249208 9648
rect 253756 9596 253808 9648
rect 513196 9596 513248 9648
rect 154396 9528 154448 9580
rect 250352 9528 250404 9580
rect 255136 9528 255188 9580
rect 516784 9528 516836 9580
rect 155776 9460 155828 9512
rect 252652 9460 252704 9512
rect 256516 9460 256568 9512
rect 520372 9460 520424 9512
rect 157064 9392 157116 9444
rect 256240 9392 256292 9444
rect 257896 9392 257948 9444
rect 523868 9392 523920 9444
rect 157156 9324 157208 9376
rect 257436 9324 257488 9376
rect 259276 9324 259328 9376
rect 527456 9324 527508 9376
rect 158444 9256 158496 9308
rect 261024 9256 261076 9308
rect 262036 9256 262088 9308
rect 534540 9256 534592 9308
rect 159824 9188 159876 9240
rect 264612 9188 264664 9240
rect 264796 9188 264848 9240
rect 541716 9188 541768 9240
rect 161204 9120 161256 9172
rect 268108 9120 268160 9172
rect 268936 9120 268988 9172
rect 552388 9120 552440 9172
rect 162676 9052 162728 9104
rect 270500 9052 270552 9104
rect 271696 9052 271748 9104
rect 559564 9052 559616 9104
rect 164056 8984 164108 9036
rect 274088 8984 274140 9036
rect 274456 8984 274508 9036
rect 566740 8984 566792 9036
rect 165436 8916 165488 8968
rect 277676 8916 277728 8968
rect 278596 8916 278648 8968
rect 577412 8916 577464 8968
rect 151636 8848 151688 8900
rect 243176 8848 243228 8900
rect 252468 8848 252520 8900
rect 509608 8848 509660 8900
rect 153016 8780 153068 8832
rect 245568 8780 245620 8832
rect 251088 8780 251140 8832
rect 506020 8780 506072 8832
rect 151544 8712 151596 8764
rect 241980 8712 242032 8764
rect 249708 8712 249760 8764
rect 502432 8712 502484 8764
rect 248328 8644 248380 8696
rect 498936 8644 498988 8696
rect 206744 8576 206796 8628
rect 388260 8576 388312 8628
rect 171048 8508 171100 8560
rect 291936 8508 291988 8560
rect 169576 8440 169628 8492
rect 288348 8440 288400 8492
rect 168196 8372 168248 8424
rect 284760 8372 284812 8424
rect 166816 8304 166868 8356
rect 281264 8304 281316 8356
rect 222016 8236 222068 8288
rect 426348 8236 426400 8288
rect 137744 8168 137796 8220
rect 206284 8168 206336 8220
rect 223488 8168 223540 8220
rect 429936 8168 429988 8220
rect 139124 8100 139176 8152
rect 209872 8100 209924 8152
rect 224868 8100 224920 8152
rect 433524 8100 433576 8152
rect 140504 8032 140556 8084
rect 213460 8032 213512 8084
rect 224776 8032 224828 8084
rect 437020 8032 437072 8084
rect 141884 7964 141936 8016
rect 217048 7964 217100 8016
rect 226248 7964 226300 8016
rect 440608 7964 440660 8016
rect 143264 7896 143316 7948
rect 220544 7896 220596 7948
rect 227628 7896 227680 7948
rect 444196 7896 444248 7948
rect 144644 7828 144696 7880
rect 224132 7828 224184 7880
rect 229008 7828 229060 7880
rect 447784 7828 447836 7880
rect 147496 7760 147548 7812
rect 228916 7760 228968 7812
rect 230296 7760 230348 7812
rect 451372 7760 451424 7812
rect 146116 7692 146168 7744
rect 227720 7692 227772 7744
rect 231768 7692 231820 7744
rect 454868 7692 454920 7744
rect 148876 7624 148928 7676
rect 232504 7624 232556 7676
rect 233056 7624 233108 7676
rect 458456 7624 458508 7676
rect 147404 7556 147456 7608
rect 231308 7556 231360 7608
rect 234528 7556 234580 7608
rect 462044 7556 462096 7608
rect 220728 7488 220780 7540
rect 422760 7488 422812 7540
rect 219348 7420 219400 7472
rect 419172 7420 419224 7472
rect 217968 7352 218020 7404
rect 415676 7352 415728 7404
rect 216588 7284 216640 7336
rect 412088 7284 412140 7336
rect 215116 7216 215168 7268
rect 408592 7216 408644 7268
rect 213828 7148 213880 7200
rect 404912 7148 404964 7200
rect 212448 7080 212500 7132
rect 401324 7080 401376 7132
rect 211068 7012 211120 7064
rect 397828 7012 397880 7064
rect 161296 6944 161348 6996
rect 267004 6944 267056 6996
rect 202788 6919 202840 6928
rect 202788 6885 202797 6919
rect 202797 6885 202831 6919
rect 202831 6885 202840 6919
rect 202788 6876 202840 6885
rect 125416 6808 125468 6860
rect 170588 6808 170640 6860
rect 184848 6808 184900 6860
rect 330024 6808 330076 6860
rect 126888 6740 126940 6792
rect 174176 6740 174228 6792
rect 186228 6740 186280 6792
rect 333612 6740 333664 6792
rect 128268 6672 128320 6724
rect 177764 6672 177816 6724
rect 187608 6672 187660 6724
rect 337108 6672 337160 6724
rect 129556 6604 129608 6656
rect 181352 6604 181404 6656
rect 188988 6604 189040 6656
rect 340696 6604 340748 6656
rect 131028 6536 131080 6588
rect 184848 6536 184900 6588
rect 190368 6536 190420 6588
rect 344284 6536 344336 6588
rect 130936 6468 130988 6520
rect 188436 6468 188488 6520
rect 193128 6468 193180 6520
rect 351368 6468 351420 6520
rect 132316 6400 132368 6452
rect 192024 6400 192076 6452
rect 194508 6400 194560 6452
rect 354956 6400 355008 6452
rect 133696 6332 133748 6384
rect 195612 6332 195664 6384
rect 195888 6332 195940 6384
rect 358544 6332 358596 6384
rect 134892 6264 134944 6316
rect 199200 6264 199252 6316
rect 200028 6264 200080 6316
rect 369216 6264 369268 6316
rect 158536 6196 158588 6248
rect 259828 6196 259880 6248
rect 273076 6196 273128 6248
rect 563152 6196 563204 6248
rect 159916 6128 159968 6180
rect 263416 6128 263468 6180
rect 277216 6128 277268 6180
rect 573824 6128 573876 6180
rect 123944 6060 123996 6112
rect 167092 6060 167144 6112
rect 175924 6060 175976 6112
rect 183468 6060 183520 6112
rect 326436 6060 326488 6112
rect 122656 5992 122708 6044
rect 163504 5992 163556 6044
rect 182088 5992 182140 6044
rect 322848 5992 322900 6044
rect 180708 5924 180760 5976
rect 319260 5924 319312 5976
rect 179328 5856 179380 5908
rect 315764 5856 315816 5908
rect 177948 5788 178000 5840
rect 312176 5788 312228 5840
rect 176568 5720 176620 5772
rect 308588 5720 308640 5772
rect 175188 5652 175240 5704
rect 305092 5652 305144 5704
rect 173808 5584 173860 5636
rect 301412 5584 301464 5636
rect 172428 5516 172480 5568
rect 297916 5516 297968 5568
rect 148968 5448 149020 5500
rect 233700 5448 233752 5500
rect 262128 5448 262180 5500
rect 533436 5448 533488 5500
rect 150164 5380 150216 5432
rect 237196 5380 237248 5432
rect 263508 5380 263560 5432
rect 536932 5380 536984 5432
rect 151728 5312 151780 5364
rect 240784 5312 240836 5364
rect 264888 5312 264940 5364
rect 540520 5312 540572 5364
rect 153108 5244 153160 5296
rect 244372 5244 244424 5296
rect 266268 5244 266320 5296
rect 544108 5244 544160 5296
rect 71872 5176 71924 5228
rect 154488 5176 154540 5228
rect 247960 5176 248012 5228
rect 267648 5176 267700 5228
rect 547696 5176 547748 5228
rect 155868 5108 155920 5160
rect 251456 5108 251508 5160
rect 269028 5108 269080 5160
rect 551192 5108 551244 5160
rect 157248 5040 157300 5092
rect 255044 5040 255096 5092
rect 270408 5040 270460 5092
rect 554780 5040 554832 5092
rect 158628 4972 158680 5024
rect 258632 4972 258684 5024
rect 271788 4972 271840 5024
rect 558368 4972 558420 5024
rect 160008 4904 160060 4956
rect 262220 4904 262272 4956
rect 273168 4904 273220 4956
rect 561956 4904 562008 4956
rect 161388 4836 161440 4888
rect 265808 4836 265860 4888
rect 274548 4836 274600 4888
rect 565544 4836 565596 4888
rect 55220 4768 55272 4820
rect 80428 4768 80480 4820
rect 90364 4768 90416 4820
rect 162768 4768 162820 4820
rect 269304 4768 269356 4820
rect 275928 4768 275980 4820
rect 569040 4768 569092 4820
rect 147588 4700 147640 4752
rect 230112 4700 230164 4752
rect 260748 4700 260800 4752
rect 529848 4700 529900 4752
rect 146208 4632 146260 4684
rect 226524 4632 226576 4684
rect 259368 4632 259420 4684
rect 526260 4632 526312 4684
rect 144736 4564 144788 4616
rect 222936 4564 222988 4616
rect 257988 4564 258040 4616
rect 522672 4564 522724 4616
rect 143356 4496 143408 4548
rect 219348 4496 219400 4548
rect 256608 4496 256660 4548
rect 519084 4496 519136 4548
rect 141976 4428 142028 4480
rect 215852 4428 215904 4480
rect 255228 4428 255280 4480
rect 515588 4428 515640 4480
rect 140596 4360 140648 4412
rect 212264 4360 212316 4412
rect 253848 4360 253900 4412
rect 512000 4360 512052 4412
rect 139216 4292 139268 4344
rect 208676 4292 208728 4344
rect 209596 4292 209648 4344
rect 394240 4292 394292 4344
rect 70584 4224 70636 4276
rect 137836 4224 137888 4276
rect 205088 4224 205140 4276
rect 205548 4224 205600 4276
rect 383568 4224 383620 4276
rect 37372 4088 37424 4140
rect 38568 4088 38620 4140
rect 119896 4156 119948 4208
rect 136548 4156 136600 4208
rect 201500 4156 201552 4208
rect 376392 4156 376444 4208
rect 72148 4088 72200 4140
rect 75184 4088 75236 4140
rect 29092 4020 29144 4072
rect 30288 4020 30340 4072
rect 78772 4020 78824 4072
rect 79048 4020 79100 4072
rect 80244 4088 80296 4140
rect 82084 4088 82136 4140
rect 83832 4088 83884 4140
rect 84844 4088 84896 4140
rect 84936 4088 84988 4140
rect 85488 4088 85540 4140
rect 88524 4088 88576 4140
rect 89628 4088 89680 4140
rect 93308 4088 93360 4140
rect 93768 4088 93820 4140
rect 96528 4088 96580 4140
rect 96896 4088 96948 4140
rect 97908 4088 97960 4140
rect 99288 4088 99340 4140
rect 100024 4088 100076 4140
rect 103980 4088 104032 4140
rect 104624 4088 104676 4140
rect 117136 4088 117188 4140
rect 117228 4088 117280 4140
rect 148324 4088 148376 4140
rect 151544 4088 151596 4140
rect 152464 4088 152516 4140
rect 155132 4088 155184 4140
rect 155224 4088 155276 4140
rect 82912 4020 82964 4072
rect 104808 4020 104860 4072
rect 118240 4020 118292 4072
rect 118516 4020 118568 4072
rect 153844 4020 153896 4072
rect 25504 3952 25556 4004
rect 69112 3952 69164 4004
rect 72056 3952 72108 4004
rect 73068 3952 73120 4004
rect 79324 3952 79376 4004
rect 85580 3952 85632 4004
rect 106096 3952 106148 4004
rect 120632 3952 120684 4004
rect 121276 3952 121328 4004
rect 159916 3952 159968 4004
rect 167644 3952 167696 4004
rect 18328 3884 18380 3936
rect 66628 3884 66680 3936
rect 67180 3884 67232 3936
rect 16028 3816 16080 3868
rect 64880 3816 64932 3868
rect 75460 3884 75512 3936
rect 85764 3884 85816 3936
rect 107568 3884 107620 3936
rect 14832 3748 14884 3800
rect 64972 3748 65024 3800
rect 10048 3680 10100 3732
rect 63592 3680 63644 3732
rect 7656 3612 7708 3664
rect 62212 3612 62264 3664
rect 62396 3612 62448 3664
rect 77944 3816 77996 3868
rect 87604 3816 87656 3868
rect 89720 3816 89772 3868
rect 92572 3816 92624 3868
rect 94504 3816 94556 3868
rect 95332 3816 95384 3868
rect 106188 3816 106240 3868
rect 121828 3816 121880 3868
rect 68284 3748 68336 3800
rect 79416 3748 79468 3800
rect 81900 3748 81952 3800
rect 107476 3748 107528 3800
rect 124220 3884 124272 3936
rect 125508 3884 125560 3936
rect 168196 3884 168248 3936
rect 169024 3952 169076 4004
rect 176476 3952 176528 4004
rect 169944 3884 169996 3936
rect 172980 3884 173032 3936
rect 182548 3952 182600 4004
rect 300308 4088 300360 4140
rect 304264 4088 304316 4140
rect 307392 4088 307444 4140
rect 193220 4020 193272 4072
rect 190828 3952 190880 4004
rect 122748 3816 122800 3868
rect 159456 3816 159508 3868
rect 164700 3816 164752 3868
rect 166264 3816 166316 3868
rect 176568 3816 176620 3868
rect 81440 3680 81492 3732
rect 82728 3680 82780 3732
rect 104716 3680 104768 3732
rect 65984 3612 66036 3664
rect 84292 3612 84344 3664
rect 102784 3612 102836 3664
rect 108764 3612 108816 3664
rect 108948 3680 109000 3732
rect 123024 3680 123076 3732
rect 6460 3544 6512 3596
rect 62120 3544 62172 3596
rect 63592 3544 63644 3596
rect 64788 3544 64840 3596
rect 84384 3544 84436 3596
rect 87328 3544 87380 3596
rect 88248 3544 88300 3596
rect 100668 3544 100720 3596
rect 106372 3544 106424 3596
rect 1676 3476 1728 3528
rect 59360 3476 59412 3528
rect 60004 3476 60056 3528
rect 572 3408 624 3460
rect 59912 3408 59964 3460
rect 61200 3408 61252 3460
rect 76656 3476 76708 3528
rect 82176 3476 82228 3528
rect 100116 3476 100168 3528
rect 101588 3476 101640 3528
rect 101956 3476 102008 3528
rect 109960 3476 110012 3528
rect 110144 3612 110196 3664
rect 131396 3748 131448 3800
rect 124128 3680 124180 3732
rect 127624 3680 127676 3732
rect 130384 3612 130436 3664
rect 169944 3748 169996 3800
rect 176844 3884 176896 3936
rect 189816 3884 189868 3936
rect 310980 4020 311032 4072
rect 289544 3952 289596 4004
rect 295984 3952 296036 4004
rect 417976 3952 418028 4004
rect 176752 3816 176804 3868
rect 332416 3884 332468 3936
rect 133788 3680 133840 3732
rect 150440 3680 150492 3732
rect 151084 3680 151136 3732
rect 157984 3680 158036 3732
rect 176016 3680 176068 3732
rect 181536 3748 181588 3800
rect 185584 3748 185636 3800
rect 190460 3748 190512 3800
rect 193864 3816 193916 3868
rect 335912 3816 335964 3868
rect 191748 3748 191800 3800
rect 346676 3748 346728 3800
rect 176936 3680 176988 3732
rect 183744 3680 183796 3732
rect 184204 3680 184256 3732
rect 200396 3680 200448 3732
rect 360936 3748 360988 3800
rect 132408 3612 132460 3664
rect 110236 3544 110288 3596
rect 132592 3544 132644 3596
rect 133144 3612 133196 3664
rect 137284 3612 137336 3664
rect 189632 3612 189684 3664
rect 189724 3612 189776 3664
rect 190276 3612 190328 3664
rect 194416 3612 194468 3664
rect 197268 3612 197320 3664
rect 356060 3680 356112 3732
rect 357348 3680 357400 3732
rect 374000 3680 374052 3732
rect 375196 3680 375248 3732
rect 206928 3612 206980 3664
rect 389456 3612 389508 3664
rect 186412 3544 186464 3596
rect 187240 3544 187292 3596
rect 196808 3544 196860 3596
rect 209688 3544 209740 3596
rect 396632 3544 396684 3596
rect 408500 3544 408552 3596
rect 409696 3544 409748 3596
rect 485780 3544 485832 3596
rect 486976 3544 487028 3596
rect 81532 3408 81584 3460
rect 82636 3408 82688 3460
rect 97816 3408 97868 3460
rect 100484 3408 100536 3460
rect 102048 3408 102100 3460
rect 111156 3408 111208 3460
rect 111708 3476 111760 3528
rect 136088 3476 136140 3528
rect 137928 3476 137980 3528
rect 203892 3476 203944 3528
rect 215208 3476 215260 3528
rect 410892 3476 410944 3528
rect 433340 3476 433392 3528
rect 434628 3476 434680 3528
rect 451280 3476 451332 3528
rect 452476 3476 452528 3528
rect 459560 3476 459612 3528
rect 460848 3476 460900 3528
rect 502340 3476 502392 3528
rect 503628 3476 503680 3528
rect 520280 3476 520332 3528
rect 521476 3476 521528 3528
rect 529480 3476 529532 3528
rect 564348 3476 564400 3528
rect 11244 3340 11296 3392
rect 12348 3340 12400 3392
rect 17224 3340 17276 3392
rect 17868 3340 17920 3392
rect 19524 3340 19576 3392
rect 20628 3340 20680 3392
rect 26700 3340 26752 3392
rect 27528 3340 27580 3392
rect 27896 3340 27948 3392
rect 33876 3340 33928 3392
rect 32680 3272 32732 3324
rect 12440 3136 12492 3188
rect 13728 3136 13780 3188
rect 36176 3272 36228 3324
rect 37188 3272 37240 3324
rect 43352 3272 43404 3324
rect 44088 3272 44140 3324
rect 44548 3272 44600 3324
rect 45468 3272 45520 3324
rect 45744 3272 45796 3324
rect 46848 3272 46900 3324
rect 50528 3272 50580 3324
rect 50988 3272 51040 3324
rect 52828 3272 52880 3324
rect 53748 3272 53800 3324
rect 42156 3204 42208 3256
rect 70676 3340 70728 3392
rect 86224 3340 86276 3392
rect 104256 3340 104308 3392
rect 112352 3340 112404 3392
rect 69480 3272 69532 3324
rect 86040 3272 86092 3324
rect 106004 3272 106056 3324
rect 112996 3408 113048 3460
rect 133696 3408 133748 3460
rect 207480 3408 207532 3460
rect 222108 3408 222160 3460
rect 428740 3408 428792 3460
rect 494060 3408 494112 3460
rect 495348 3408 495400 3460
rect 529388 3408 529440 3460
rect 571432 3408 571484 3460
rect 119436 3340 119488 3392
rect 127808 3340 127860 3392
rect 115940 3272 115992 3324
rect 116952 3272 117004 3324
rect 145840 3272 145892 3324
rect 148048 3272 148100 3324
rect 166356 3340 166408 3392
rect 178960 3340 179012 3392
rect 180064 3340 180116 3392
rect 182824 3340 182876 3392
rect 186136 3340 186188 3392
rect 271696 3340 271748 3392
rect 275284 3340 275336 3392
rect 382372 3340 382424 3392
rect 390652 3340 390704 3392
rect 391848 3340 391900 3392
rect 156328 3272 156380 3324
rect 48136 3136 48188 3188
rect 74908 3204 74960 3256
rect 77484 3204 77536 3256
rect 77852 3204 77904 3256
rect 88432 3204 88484 3256
rect 103428 3204 103480 3256
rect 114744 3204 114796 3256
rect 115848 3204 115900 3256
rect 145656 3204 145708 3256
rect 152556 3204 152608 3256
rect 186320 3272 186372 3324
rect 186412 3272 186464 3324
rect 282460 3272 282512 3324
rect 293132 3272 293184 3324
rect 293224 3272 293276 3324
rect 400220 3272 400272 3324
rect 176660 3204 176712 3256
rect 186044 3204 186096 3256
rect 253848 3204 253900 3256
rect 255964 3204 256016 3256
rect 339500 3204 339552 3256
rect 347780 3204 347832 3256
rect 349068 3204 349120 3256
rect 77300 3136 77352 3188
rect 103336 3136 103388 3188
rect 113548 3136 113600 3188
rect 114284 3136 114336 3188
rect 143264 3136 143316 3188
rect 152740 3136 152792 3188
rect 157524 3136 157576 3188
rect 246764 3136 246816 3188
rect 253204 3136 253256 3188
rect 328828 3136 328880 3188
rect 8852 3068 8904 3120
rect 9588 3068 9640 3120
rect 49332 3068 49384 3120
rect 104164 3068 104216 3120
rect 107568 3068 107620 3120
rect 110328 3068 110380 3120
rect 130200 3068 130252 3120
rect 138480 3068 138532 3120
rect 160744 3068 160796 3120
rect 164884 3068 164936 3120
rect 175372 3068 175424 3120
rect 51632 3000 51684 3052
rect 77392 3000 77444 3052
rect 86132 3000 86184 3052
rect 92664 3000 92716 3052
rect 114376 3000 114428 3052
rect 142068 3000 142120 3052
rect 149244 3000 149296 3052
rect 20720 2932 20772 2984
rect 22008 2932 22060 2984
rect 54024 2932 54076 2984
rect 80060 2932 80112 2984
rect 113088 2932 113140 2984
rect 139676 2932 139728 2984
rect 46940 2864 46992 2916
rect 56416 2864 56468 2916
rect 80152 2864 80204 2916
rect 111616 2864 111668 2916
rect 134892 2864 134944 2916
rect 139308 2864 139360 2916
rect 145564 2864 145616 2916
rect 176568 3000 176620 3052
rect 236000 3068 236052 3120
rect 271236 3068 271288 3120
rect 291844 3068 291896 3120
rect 368020 3068 368072 3120
rect 58808 2796 58860 2848
rect 83096 2796 83148 2848
rect 95424 2796 95476 2848
rect 95700 2796 95752 2848
rect 108856 2796 108908 2848
rect 126612 2796 126664 2848
rect 129556 2796 129608 2848
rect 129648 2796 129700 2848
rect 133972 2796 134024 2848
rect 148416 2796 148468 2848
rect 171784 2932 171836 2984
rect 173164 2932 173216 2984
rect 239588 3000 239640 3052
rect 250444 3000 250496 3052
rect 325240 3000 325292 3052
rect 176752 2932 176804 2984
rect 225328 2932 225380 2984
rect 253296 2932 253348 2984
rect 278872 2932 278924 2984
rect 289084 2932 289136 2984
rect 353760 2932 353812 2984
rect 165896 2864 165948 2916
rect 202696 2864 202748 2916
rect 246304 2864 246356 2916
rect 275284 2864 275336 2916
rect 156604 2796 156656 2848
rect 198004 2796 198056 2848
rect 271144 2796 271196 2848
rect 285956 2864 286008 2916
rect 286324 2864 286376 2916
rect 303804 2864 303856 2916
rect 305000 2864 305052 2916
rect 306196 2864 306248 2916
rect 279424 2796 279476 2848
rect 296720 2796 296772 2848
rect 180156 2728 180208 2780
rect 273444 2320 273496 2372
rect 280068 2320 280120 2372
rect 365720 1368 365772 1420
rect 366916 1368 366968 1420
rect 5264 552 5316 604
rect 5448 552 5500 604
rect 23112 552 23164 604
rect 23388 552 23440 604
rect 92112 552 92164 604
rect 92388 552 92440 604
rect 95424 552 95476 604
rect 95700 552 95752 604
rect 128636 552 128688 604
rect 129004 552 129056 604
rect 140872 595 140924 604
rect 140872 561 140881 595
rect 140881 561 140915 595
rect 140915 561 140924 595
rect 140872 552 140924 561
rect 295340 552 295392 604
rect 295524 552 295576 604
rect 298100 552 298152 604
rect 299112 552 299164 604
rect 309140 552 309192 604
rect 309784 552 309836 604
rect 316040 552 316092 604
rect 316960 552 317012 604
rect 317420 552 317472 604
rect 318064 552 318116 604
rect 322940 552 322992 604
rect 324044 552 324096 604
rect 327080 552 327132 604
rect 327632 552 327684 604
rect 333980 552 334032 604
rect 334716 552 334768 604
rect 340880 552 340932 604
rect 341892 552 341944 604
rect 342260 552 342312 604
rect 343088 552 343140 604
rect 364340 552 364392 604
rect 364524 552 364576 604
rect 369860 552 369912 604
rect 370412 552 370464 604
rect 376760 552 376812 604
rect 377588 552 377640 604
rect 378140 552 378192 604
rect 378784 552 378836 604
rect 412640 552 412692 604
rect 413284 552 413336 604
rect 419540 552 419592 604
rect 420368 552 420420 604
rect 420920 552 420972 604
rect 421564 552 421616 604
rect 423680 552 423732 604
rect 423956 552 424008 604
rect 426440 552 426492 604
rect 427544 552 427596 604
rect 430580 552 430632 604
rect 431132 552 431184 604
rect 438860 552 438912 604
rect 439412 552 439464 604
rect 441620 552 441672 604
rect 441804 552 441856 604
rect 444380 552 444432 604
rect 445392 552 445444 604
rect 445760 552 445812 604
rect 446588 552 446640 604
rect 448520 552 448572 604
rect 448980 552 449032 604
rect 452660 552 452712 604
rect 453672 552 453724 604
rect 455420 552 455472 604
rect 456064 552 456116 604
rect 462320 552 462372 604
rect 463240 552 463292 604
rect 466460 552 466512 604
rect 466828 552 466880 604
rect 469220 552 469272 604
rect 470324 552 470376 604
rect 489920 552 489972 604
rect 490564 552 490616 604
rect 495440 552 495492 604
rect 496544 552 496596 604
rect 496820 552 496872 604
rect 497740 552 497792 604
rect 499580 552 499632 604
rect 500132 552 500184 604
rect 500960 552 501012 604
rect 501236 552 501288 604
rect 503720 552 503772 604
rect 504824 552 504876 604
rect 506480 552 506532 604
rect 507216 552 507268 604
rect 507860 552 507912 604
rect 508412 552 508464 604
rect 510620 552 510672 604
rect 510804 552 510856 604
rect 513380 552 513432 604
rect 514392 552 514444 604
rect 524420 552 524472 604
rect 525064 552 525116 604
rect 538220 552 538272 604
rect 539324 552 539376 604
rect 542360 552 542412 604
rect 542912 552 542964 604
rect 549260 552 549312 604
rect 550088 552 550140 604
rect 556160 552 556212 604
rect 557172 552 557224 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 264888 653404 264940 653410
rect 264888 653346 264940 653352
rect 378140 653404 378192 653410
rect 378140 653346 378192 653352
rect 383568 653404 383620 653410
rect 383568 653346 383620 653352
rect 508412 653404 508464 653410
rect 508412 653346 508464 653352
rect 264900 652934 264928 653346
rect 378152 652934 378180 653346
rect 383580 652934 383608 653346
rect 259184 652928 259236 652934
rect 129278 652896 129334 652905
rect 129278 652831 129334 652840
rect 133694 652896 133750 652905
rect 133694 652831 133750 652840
rect 259182 652896 259184 652905
rect 263600 652928 263652 652934
rect 259236 652896 259238 652905
rect 259182 652831 259238 652840
rect 263598 652896 263600 652905
rect 264888 652928 264940 652934
rect 263652 652896 263654 652905
rect 378140 652928 378192 652934
rect 264888 652870 264940 652876
rect 378138 652896 378140 652905
rect 383568 652928 383620 652934
rect 378192 652896 378194 652905
rect 263598 652831 263654 652840
rect 378138 652831 378194 652840
rect 383566 652896 383568 652905
rect 508424 652905 508452 653346
rect 383620 652896 383622 652905
rect 383566 652831 383622 652840
rect 508410 652896 508466 652905
rect 508410 652831 508412 652840
rect 129292 652798 129320 652831
rect 133708 652798 133736 652831
rect 383580 652805 383608 652831
rect 508464 652831 508466 652840
rect 513378 652896 513434 652905
rect 513378 652831 513380 652840
rect 508412 652802 508464 652808
rect 513432 652831 513434 652840
rect 513380 652802 513432 652808
rect 129280 652792 129332 652798
rect 129280 652734 129332 652740
rect 133696 652792 133748 652798
rect 133696 652734 133748 652740
rect 139400 652792 139452 652798
rect 508424 652771 508452 652802
rect 518900 652792 518952 652798
rect 139400 652734 139452 652740
rect 518900 652734 518952 652740
rect 139412 650570 139440 652734
rect 139320 650542 139440 650570
rect 266452 650548 266504 650554
rect 137652 650480 137704 650486
rect 137652 650422 137704 650428
rect 137664 649720 137692 650422
rect 139320 649754 139348 650542
rect 266452 650490 266504 650496
rect 266464 650282 266492 650490
rect 282828 650480 282880 650486
rect 282828 650422 282880 650428
rect 516416 650480 516468 650486
rect 516416 650422 516468 650428
rect 266452 650276 266504 650282
rect 266452 650218 266504 650224
rect 266464 649913 266492 650218
rect 282840 650214 282868 650422
rect 387156 650276 387208 650282
rect 387156 650218 387208 650224
rect 282276 650208 282328 650214
rect 282276 650150 282328 650156
rect 282828 650208 282880 650214
rect 282828 650150 282880 650156
rect 266450 649904 266506 649913
rect 266450 649839 266506 649848
rect 139320 649726 139440 649754
rect 137650 649711 137706 649720
rect 137650 649646 137706 649655
rect 57886 646096 57942 646105
rect 57886 646031 57942 646040
rect 57794 645008 57850 645017
rect 57794 644943 57850 644952
rect 57702 643240 57758 643249
rect 57702 643175 57758 643184
rect 57610 642016 57666 642025
rect 57610 641951 57666 641960
rect 57518 640384 57574 640393
rect 57518 640319 57574 640328
rect 57426 639296 57482 639305
rect 57426 639231 57482 639240
rect 57334 637664 57390 637673
rect 57334 637599 57390 637608
rect 57242 579728 57298 579737
rect 57242 579663 57298 579672
rect 57256 543114 57284 579663
rect 57244 543108 57296 543114
rect 57244 543050 57296 543056
rect 57348 542978 57376 637599
rect 57440 543522 57468 639231
rect 57428 543516 57480 543522
rect 57428 543458 57480 543464
rect 57532 543454 57560 640319
rect 57520 543448 57572 543454
rect 57520 543390 57572 543396
rect 57624 543386 57652 641951
rect 57612 543380 57664 543386
rect 57612 543322 57664 543328
rect 57716 543250 57744 643175
rect 57808 543862 57836 644943
rect 57900 543930 57928 646031
rect 139412 589665 139440 649726
rect 282288 648689 282316 650150
rect 387168 649913 387196 650218
rect 516428 649913 516456 650422
rect 387154 649904 387210 649913
rect 387154 649839 387210 649848
rect 516414 649904 516470 649913
rect 516414 649839 516470 649848
rect 282274 648680 282330 648689
rect 282274 648615 282330 648624
rect 188342 646096 188398 646105
rect 188342 646031 188398 646040
rect 307390 646096 307446 646105
rect 307390 646031 307446 646040
rect 438122 646096 438178 646105
rect 438122 646031 438178 646040
rect 139398 589656 139454 589665
rect 139398 589591 139454 589600
rect 139398 580408 139454 580417
rect 139398 580343 139454 580352
rect 139412 579630 139440 580343
rect 139400 579624 139452 579630
rect 139400 579566 139452 579572
rect 187700 579624 187752 579630
rect 187700 579566 187752 579572
rect 187712 579057 187740 579566
rect 187698 579048 187754 579057
rect 187698 578983 187754 578992
rect 67546 558920 67602 558929
rect 66168 558884 66220 558890
rect 67546 558855 67602 558864
rect 68926 558920 68982 558929
rect 68926 558855 68982 558864
rect 70214 558920 70270 558929
rect 70214 558855 70270 558864
rect 71686 558920 71742 558929
rect 71686 558855 71742 558864
rect 72514 558920 72570 558929
rect 72514 558855 72570 558864
rect 73066 558920 73122 558929
rect 73066 558855 73122 558864
rect 73710 558920 73766 558929
rect 73710 558855 73766 558864
rect 74262 558920 74318 558929
rect 74262 558855 74318 558864
rect 74998 558920 75054 558929
rect 74998 558855 75054 558864
rect 75826 558920 75882 558929
rect 75826 558855 75882 558864
rect 76838 558920 76894 558929
rect 76838 558855 76894 558864
rect 77390 558920 77446 558929
rect 77390 558855 77446 558864
rect 78586 558920 78642 558929
rect 78586 558855 78642 558864
rect 79322 558920 79378 558929
rect 79322 558855 79378 558864
rect 79966 558920 80022 558929
rect 79966 558855 80022 558864
rect 80794 558920 80850 558929
rect 80794 558855 80850 558864
rect 81254 558920 81310 558929
rect 81254 558855 81310 558864
rect 81990 558920 82046 558929
rect 81990 558855 82046 558864
rect 82726 558920 82782 558929
rect 82726 558855 82782 558864
rect 83830 558920 83886 558929
rect 83830 558855 83886 558864
rect 84198 558920 84254 558929
rect 84198 558855 84254 558864
rect 85486 558920 85542 558929
rect 85486 558855 85542 558864
rect 86774 558920 86830 558929
rect 86774 558855 86830 558864
rect 87878 558920 87934 558929
rect 87878 558855 87934 558864
rect 88246 558920 88302 558929
rect 88246 558855 88302 558864
rect 88890 558920 88946 558929
rect 88890 558855 88946 558864
rect 89350 558920 89406 558929
rect 89350 558855 89406 558864
rect 89810 558920 89866 558929
rect 89810 558855 89866 558864
rect 91006 558920 91062 558929
rect 91006 558855 91062 558864
rect 92294 558920 92350 558929
rect 92294 558855 92350 558864
rect 92478 558920 92534 558929
rect 92478 558855 92534 558864
rect 93674 558920 93730 558929
rect 93674 558855 93730 558864
rect 94870 558920 94926 558929
rect 94870 558855 94926 558864
rect 95054 558920 95110 558929
rect 95054 558855 95110 558864
rect 95698 558920 95754 558929
rect 95698 558855 95754 558864
rect 96526 558920 96582 558929
rect 96526 558855 96582 558864
rect 97078 558920 97134 558929
rect 97078 558855 97134 558864
rect 97630 558920 97686 558929
rect 97630 558855 97686 558864
rect 98550 558920 98606 558929
rect 98550 558855 98606 558864
rect 99286 558920 99342 558929
rect 99286 558855 99342 558864
rect 100574 558920 100630 558929
rect 100574 558855 100630 558864
rect 102046 558920 102102 558929
rect 102046 558855 102102 558864
rect 104806 558920 104862 558929
rect 104806 558855 104862 558864
rect 107474 558920 107530 558929
rect 107474 558855 107530 558864
rect 108486 558920 108542 558929
rect 108486 558855 108542 558864
rect 66168 558826 66220 558832
rect 62026 558376 62082 558385
rect 62026 558311 62082 558320
rect 57888 543924 57940 543930
rect 57888 543866 57940 543872
rect 57796 543856 57848 543862
rect 57796 543798 57848 543804
rect 62040 543590 62068 558311
rect 63406 558240 63462 558249
rect 63406 558175 63462 558184
rect 61016 543584 61068 543590
rect 61016 543526 61068 543532
rect 62028 543584 62080 543590
rect 62028 543526 62080 543532
rect 57704 543244 57756 543250
rect 57704 543186 57756 543192
rect 57336 542972 57388 542978
rect 57336 542914 57388 542920
rect 61028 539988 61056 543526
rect 63420 540002 63448 558175
rect 66180 543590 66208 558826
rect 67456 558816 67508 558822
rect 67456 558758 67508 558764
rect 65156 543584 65208 543590
rect 65156 543526 65208 543532
rect 66168 543584 66220 543590
rect 66168 543526 66220 543532
rect 63066 539974 63448 540002
rect 65168 539988 65196 543526
rect 67468 540002 67496 558758
rect 67560 543046 67588 558855
rect 67548 543040 67600 543046
rect 67548 542982 67600 542988
rect 68940 542450 68968 558855
rect 70228 542706 70256 558855
rect 70306 558784 70362 558793
rect 70306 558719 70362 558728
rect 70320 543590 70348 558719
rect 71700 543726 71728 558855
rect 72528 558210 72556 558855
rect 72516 558204 72568 558210
rect 72516 558146 72568 558152
rect 73080 543998 73108 558855
rect 73724 558414 73752 558855
rect 73712 558408 73764 558414
rect 73712 558350 73764 558356
rect 74276 558278 74304 558855
rect 74264 558272 74316 558278
rect 74264 558214 74316 558220
rect 75012 557938 75040 558855
rect 75000 557932 75052 557938
rect 75000 557874 75052 557880
rect 73068 543992 73120 543998
rect 73068 543934 73120 543940
rect 75840 543726 75868 558855
rect 75918 558784 75974 558793
rect 75918 558719 75974 558728
rect 75932 558550 75960 558719
rect 75920 558544 75972 558550
rect 75920 558486 75972 558492
rect 76852 558142 76880 558855
rect 77404 558618 77432 558855
rect 78494 558784 78550 558793
rect 78494 558719 78550 558728
rect 78508 558686 78536 558719
rect 78496 558680 78548 558686
rect 78496 558622 78548 558628
rect 77392 558612 77444 558618
rect 77392 558554 77444 558560
rect 76840 558136 76892 558142
rect 76840 558078 76892 558084
rect 71688 543720 71740 543726
rect 71688 543662 71740 543668
rect 75460 543720 75512 543726
rect 75460 543662 75512 543668
rect 75828 543720 75880 543726
rect 75828 543662 75880 543668
rect 70308 543584 70360 543590
rect 70308 543526 70360 543532
rect 71320 543584 71372 543590
rect 71320 543526 71372 543532
rect 70216 542700 70268 542706
rect 70216 542642 70268 542648
rect 68940 542422 69060 542450
rect 67206 539974 67496 540002
rect 69032 540002 69060 542422
rect 69032 539974 69322 540002
rect 71332 539988 71360 543526
rect 73436 542700 73488 542706
rect 73436 542642 73488 542648
rect 73448 539988 73476 542642
rect 75472 539988 75500 543662
rect 78600 543658 78628 558855
rect 79336 558006 79364 558855
rect 79506 558784 79562 558793
rect 79506 558719 79508 558728
rect 79560 558719 79562 558728
rect 79508 558690 79560 558696
rect 79324 558000 79376 558006
rect 79324 557942 79376 557948
rect 78588 543652 78640 543658
rect 78588 543594 78640 543600
rect 79980 543590 80008 558855
rect 80808 558482 80836 558855
rect 80796 558476 80848 558482
rect 80796 558418 80848 558424
rect 81268 558074 81296 558855
rect 82004 558346 82032 558855
rect 81440 558340 81492 558346
rect 81440 558282 81492 558288
rect 81992 558340 82044 558346
rect 81992 558282 82044 558288
rect 81452 558210 81480 558282
rect 81440 558204 81492 558210
rect 81440 558146 81492 558152
rect 81256 558068 81308 558074
rect 81256 558010 81308 558016
rect 81716 544400 81768 544406
rect 81716 544342 81768 544348
rect 79968 543584 80020 543590
rect 79968 543526 80020 543532
rect 79692 543108 79744 543114
rect 79692 543050 79744 543056
rect 77574 543008 77630 543017
rect 77574 542943 77630 542952
rect 77588 539988 77616 542943
rect 79704 539988 79732 543050
rect 81728 539988 81756 544342
rect 82740 544066 82768 558855
rect 82910 558784 82966 558793
rect 82910 558719 82966 558728
rect 82924 558414 82952 558719
rect 82912 558408 82964 558414
rect 82912 558350 82964 558356
rect 83844 558210 83872 558855
rect 83832 558204 83884 558210
rect 83832 558146 83884 558152
rect 84212 557938 84240 558855
rect 85394 558784 85450 558793
rect 85394 558719 85450 558728
rect 85408 558550 85436 558719
rect 85396 558544 85448 558550
rect 85396 558486 85448 558492
rect 84200 557932 84252 557938
rect 84200 557874 84252 557880
rect 84212 557598 84240 557874
rect 84200 557592 84252 557598
rect 84200 557534 84252 557540
rect 83832 544468 83884 544474
rect 83832 544410 83884 544416
rect 82728 544060 82780 544066
rect 82728 544002 82780 544008
rect 83844 539988 83872 544410
rect 85500 544134 85528 558855
rect 86682 558648 86738 558657
rect 86682 558583 86684 558592
rect 86736 558583 86738 558592
rect 86684 558554 86736 558560
rect 86696 558482 86724 558554
rect 86684 558476 86736 558482
rect 86684 558418 86736 558424
rect 85856 544536 85908 544542
rect 85856 544478 85908 544484
rect 85488 544128 85540 544134
rect 85488 544070 85540 544076
rect 85868 539988 85896 544478
rect 86788 544338 86816 558855
rect 86866 558784 86922 558793
rect 86866 558719 86922 558728
rect 86776 544332 86828 544338
rect 86776 544274 86828 544280
rect 86880 544202 86908 558719
rect 87892 558686 87920 558855
rect 87880 558680 87932 558686
rect 87880 558622 87932 558628
rect 87972 544672 88024 544678
rect 87972 544614 88024 544620
rect 86868 544196 86920 544202
rect 86868 544138 86920 544144
rect 87984 539988 88012 544614
rect 88260 544270 88288 558855
rect 88904 558754 88932 558855
rect 88892 558748 88944 558754
rect 88892 558690 88944 558696
rect 89364 557802 89392 558855
rect 89824 558482 89852 558855
rect 89812 558476 89864 558482
rect 89812 558418 89864 558424
rect 89824 557938 89852 558418
rect 89812 557932 89864 557938
rect 89812 557874 89864 557880
rect 89352 557796 89404 557802
rect 89352 557738 89404 557744
rect 89996 544808 90048 544814
rect 89996 544750 90048 544756
rect 88248 544264 88300 544270
rect 88248 544206 88300 544212
rect 90008 539988 90036 544750
rect 91020 543318 91048 558855
rect 91098 558784 91154 558793
rect 91098 558719 91154 558728
rect 91112 558346 91140 558719
rect 92308 558346 92336 558855
rect 91100 558340 91152 558346
rect 91100 558282 91152 558288
rect 92296 558340 92348 558346
rect 92296 558282 92348 558288
rect 91112 557734 91140 558282
rect 91100 557728 91152 557734
rect 91100 557670 91152 557676
rect 92492 557666 92520 558855
rect 93582 558648 93638 558657
rect 93582 558583 93638 558592
rect 92480 557660 92532 557666
rect 92480 557602 92532 557608
rect 93596 557598 93624 558583
rect 93584 557592 93636 557598
rect 93584 557534 93636 557540
rect 92112 544876 92164 544882
rect 92112 544818 92164 544824
rect 91008 543312 91060 543318
rect 91008 543254 91060 543260
rect 92124 539988 92152 544818
rect 93688 543182 93716 558855
rect 93766 558784 93822 558793
rect 93766 558719 93822 558728
rect 93780 557938 93808 558719
rect 94884 558618 94912 558855
rect 94872 558612 94924 558618
rect 94872 558554 94924 558560
rect 93768 557932 93820 557938
rect 93768 557874 93820 557880
rect 94136 545012 94188 545018
rect 94136 544954 94188 544960
rect 93676 543176 93728 543182
rect 93676 543118 93728 543124
rect 94148 539988 94176 544954
rect 95068 543114 95096 558855
rect 95712 558550 95740 558855
rect 95700 558544 95752 558550
rect 95700 558486 95752 558492
rect 96540 545086 96568 558855
rect 97092 558686 97120 558855
rect 97080 558680 97132 558686
rect 97080 558622 97132 558628
rect 97092 557802 97120 558622
rect 97644 558414 97672 558855
rect 98564 558754 98592 558855
rect 98552 558748 98604 558754
rect 98552 558690 98604 558696
rect 97632 558408 97684 558414
rect 97632 558350 97684 558356
rect 97080 557796 97132 557802
rect 97080 557738 97132 557744
rect 96528 545080 96580 545086
rect 96528 545022 96580 545028
rect 96250 543280 96306 543289
rect 96250 543215 96306 543224
rect 95056 543108 95108 543114
rect 95056 543050 95108 543056
rect 96264 539988 96292 543215
rect 99300 543046 99328 558855
rect 99378 558512 99434 558521
rect 100588 558482 100616 558855
rect 102060 558686 102088 558855
rect 102048 558680 102100 558686
rect 102048 558622 102100 558628
rect 104820 558618 104848 558855
rect 104898 558784 104954 558793
rect 104898 558719 104900 558728
rect 104952 558719 104954 558728
rect 104900 558690 104952 558696
rect 102784 558612 102836 558618
rect 102784 558554 102836 558560
rect 104808 558612 104860 558618
rect 104808 558554 104860 558560
rect 99378 558447 99380 558456
rect 99432 558447 99434 558456
rect 100116 558476 100168 558482
rect 99380 558418 99432 558424
rect 100116 558418 100168 558424
rect 100576 558476 100628 558482
rect 100576 558418 100628 558424
rect 100022 557832 100078 557841
rect 100022 557767 100078 557776
rect 100036 557734 100064 557767
rect 100128 557734 100156 558418
rect 100024 557728 100076 557734
rect 100024 557670 100076 557676
rect 100116 557728 100168 557734
rect 100116 557670 100168 557676
rect 100850 557696 100906 557705
rect 98368 543040 98420 543046
rect 98368 542982 98420 542988
rect 99288 543040 99340 543046
rect 99288 542982 99340 542988
rect 98380 539988 98408 542982
rect 100036 542706 100064 557670
rect 100850 557631 100852 557640
rect 100904 557631 100906 557640
rect 101402 557696 101458 557705
rect 101402 557631 101458 557640
rect 100852 557602 100904 557608
rect 100392 542972 100444 542978
rect 100392 542914 100444 542920
rect 100024 542700 100076 542706
rect 100024 542642 100076 542648
rect 100404 539988 100432 542914
rect 101416 542638 101444 557631
rect 102796 557569 102824 558554
rect 104164 558544 104216 558550
rect 104164 558486 104216 558492
rect 104176 557569 104204 558486
rect 106280 557796 106332 557802
rect 106280 557738 106332 557744
rect 106292 557705 106320 557738
rect 106278 557696 106334 557705
rect 106278 557631 106334 557640
rect 106922 557696 106978 557705
rect 106922 557631 106978 557640
rect 102046 557560 102102 557569
rect 102046 557495 102102 557504
rect 102782 557560 102838 557569
rect 102782 557495 102838 557504
rect 103426 557560 103482 557569
rect 103426 557495 103482 557504
rect 104162 557560 104218 557569
rect 104162 557495 104218 557504
rect 105542 557560 105598 557569
rect 105542 557495 105598 557504
rect 106186 557560 106242 557569
rect 106186 557495 106242 557504
rect 102060 544950 102088 557495
rect 102048 544944 102100 544950
rect 102048 544886 102100 544892
rect 102508 543516 102560 543522
rect 102508 543458 102560 543464
rect 101404 542632 101456 542638
rect 101404 542574 101456 542580
rect 102520 539988 102548 543458
rect 102796 542774 102824 557495
rect 103440 543153 103468 557495
rect 103426 543144 103482 543153
rect 103426 543079 103482 543088
rect 104176 542842 104204 557495
rect 104532 543448 104584 543454
rect 104532 543390 104584 543396
rect 104164 542836 104216 542842
rect 104164 542778 104216 542784
rect 102784 542768 102836 542774
rect 102784 542710 102836 542716
rect 104544 539988 104572 543390
rect 105556 542910 105584 557495
rect 106200 544746 106228 557495
rect 106188 544740 106240 544746
rect 106188 544682 106240 544688
rect 106648 543380 106700 543386
rect 106648 543322 106700 543328
rect 105544 542904 105596 542910
rect 105544 542846 105596 542852
rect 106660 539988 106688 543322
rect 106936 542502 106964 557631
rect 107488 557598 107516 558855
rect 108500 558550 108528 558855
rect 125508 558748 125560 558754
rect 125508 558690 125560 558696
rect 108488 558544 108540 558550
rect 108302 558512 108358 558521
rect 108488 558486 108540 558492
rect 108302 558447 108358 558456
rect 107660 557864 107712 557870
rect 107660 557806 107712 557812
rect 107476 557592 107528 557598
rect 107672 557569 107700 557806
rect 108316 557734 108344 558447
rect 121368 557796 121420 557802
rect 121368 557738 121420 557744
rect 108304 557728 108356 557734
rect 108304 557670 108356 557676
rect 117228 557728 117280 557734
rect 117228 557670 117280 557676
rect 107476 557534 107528 557540
rect 107658 557560 107714 557569
rect 107658 557495 107714 557504
rect 108316 542570 108344 557670
rect 108486 557560 108542 557569
rect 108486 557495 108542 557504
rect 110326 557560 110382 557569
rect 110326 557495 110382 557504
rect 108500 547890 108528 557495
rect 108500 547862 108620 547890
rect 108592 542978 108620 547862
rect 110340 544610 110368 557495
rect 110328 544604 110380 544610
rect 110328 544546 110380 544552
rect 112812 543924 112864 543930
rect 112812 543866 112864 543872
rect 110788 543856 110840 543862
rect 110788 543798 110840 543804
rect 108672 543244 108724 543250
rect 108672 543186 108724 543192
rect 108580 542972 108632 542978
rect 108580 542914 108632 542920
rect 108304 542564 108356 542570
rect 108304 542506 108356 542512
rect 106924 542496 106976 542502
rect 106924 542438 106976 542444
rect 108684 539988 108712 543186
rect 110800 539988 110828 543798
rect 112824 539988 112852 543866
rect 114928 543244 114980 543250
rect 114928 543186 114980 543192
rect 114940 539988 114968 543186
rect 117240 540002 117268 557670
rect 119068 543380 119120 543386
rect 119068 543322 119120 543328
rect 117070 539974 117268 540002
rect 119080 539988 119108 543322
rect 121380 540002 121408 557738
rect 123208 543448 123260 543454
rect 123208 543390 123260 543396
rect 121210 539974 121408 540002
rect 123220 539988 123248 543390
rect 125520 540002 125548 558690
rect 140044 558680 140096 558686
rect 140044 558622 140096 558628
rect 138664 558408 138716 558414
rect 138664 558350 138716 558356
rect 137468 558340 137520 558346
rect 137468 558282 137520 558288
rect 137376 558272 137428 558278
rect 137376 558214 137428 558220
rect 137284 557932 137336 557938
rect 137284 557874 137336 557880
rect 129740 557660 129792 557666
rect 129740 557602 129792 557608
rect 129752 557546 129780 557602
rect 129660 557518 129780 557546
rect 131764 557524 131816 557530
rect 127348 543516 127400 543522
rect 127348 543458 127400 543464
rect 125350 539974 125548 540002
rect 127360 539988 127388 543458
rect 129660 540002 129688 557518
rect 131764 557466 131816 557472
rect 131776 542706 131804 557466
rect 137296 542774 137324 557874
rect 135720 542768 135772 542774
rect 135720 542710 135772 542716
rect 137284 542768 137336 542774
rect 137284 542710 137336 542716
rect 131488 542700 131540 542706
rect 131488 542642 131540 542648
rect 131764 542700 131816 542706
rect 131764 542642 131816 542648
rect 129490 539974 129688 540002
rect 131500 539988 131528 542642
rect 133604 542632 133656 542638
rect 133604 542574 133656 542580
rect 133616 539988 133644 542574
rect 135732 539988 135760 542710
rect 137388 542434 137416 558214
rect 137480 542638 137508 558282
rect 138676 542842 138704 558350
rect 140056 543697 140084 558622
rect 144184 558612 144236 558618
rect 144184 558554 144236 558560
rect 140136 558476 140188 558482
rect 140136 558418 140188 558424
rect 140042 543688 140098 543697
rect 140042 543623 140098 543632
rect 140148 542910 140176 558418
rect 141424 557592 141476 557598
rect 141424 557534 141476 557540
rect 141436 543425 141464 557534
rect 141422 543416 141478 543425
rect 141422 543351 141478 543360
rect 144196 542978 144224 558554
rect 148324 558544 148376 558550
rect 148324 558486 148376 558492
rect 145564 558136 145616 558142
rect 145564 558078 145616 558084
rect 145576 543726 145604 558078
rect 148140 543992 148192 543998
rect 148140 543934 148192 543940
rect 145564 543720 145616 543726
rect 145564 543662 145616 543668
rect 144000 542972 144052 542978
rect 144000 542914 144052 542920
rect 144184 542972 144236 542978
rect 144184 542914 144236 542920
rect 139860 542904 139912 542910
rect 139860 542846 139912 542852
rect 140136 542904 140188 542910
rect 140136 542846 140188 542852
rect 137744 542836 137796 542842
rect 137744 542778 137796 542784
rect 138664 542836 138716 542842
rect 138664 542778 138716 542784
rect 137468 542632 137520 542638
rect 137468 542574 137520 542580
rect 137376 542428 137428 542434
rect 137376 542370 137428 542376
rect 137756 539988 137784 542778
rect 139872 539988 139900 542846
rect 141884 542496 141936 542502
rect 141884 542438 141936 542444
rect 141896 539988 141924 542438
rect 144012 539988 144040 542914
rect 146024 542564 146076 542570
rect 146024 542506 146076 542512
rect 146036 539988 146064 542506
rect 148152 539988 148180 543934
rect 148336 543561 148364 558486
rect 149704 558204 149756 558210
rect 149704 558146 149756 558152
rect 148322 543552 148378 543561
rect 148322 543487 148378 543496
rect 149716 542502 149744 558146
rect 152556 558068 152608 558074
rect 152556 558010 152608 558016
rect 152464 558000 152516 558006
rect 152464 557942 152516 557948
rect 152476 543590 152504 557942
rect 152568 543726 152596 558010
rect 173072 544332 173124 544338
rect 173072 544274 173124 544280
rect 170956 544196 171008 544202
rect 170956 544138 171008 544144
rect 168840 544128 168892 544134
rect 168840 544070 168892 544076
rect 164700 544060 164752 544066
rect 164700 544002 164752 544008
rect 152556 543720 152608 543726
rect 152556 543662 152608 543668
rect 162676 543720 162728 543726
rect 162676 543662 162728 543668
rect 156420 543652 156472 543658
rect 156420 543594 156472 543600
rect 152464 543584 152516 543590
rect 152464 543526 152516 543532
rect 152280 542564 152332 542570
rect 152280 542506 152332 542512
rect 154396 542564 154448 542570
rect 154396 542506 154448 542512
rect 149704 542496 149756 542502
rect 149704 542438 149756 542444
rect 150164 542428 150216 542434
rect 150164 542370 150216 542376
rect 150176 539988 150204 542370
rect 152292 539988 152320 542506
rect 154408 539988 154436 542506
rect 156432 539988 156460 543594
rect 158536 543584 158588 543590
rect 158536 543526 158588 543532
rect 158548 539988 158576 543526
rect 160560 542428 160612 542434
rect 160560 542370 160612 542376
rect 160572 539988 160600 542370
rect 162688 539988 162716 543662
rect 164712 539988 164740 544002
rect 166816 542564 166868 542570
rect 166816 542506 166868 542512
rect 166828 539988 166856 542506
rect 168852 539988 168880 544070
rect 170968 539988 170996 544138
rect 173084 539988 173112 544274
rect 175096 544264 175148 544270
rect 175096 544206 175148 544212
rect 175108 539988 175136 544206
rect 179236 543312 179288 543318
rect 188356 543289 188384 646031
rect 307404 645930 307432 646031
rect 294696 645924 294748 645930
rect 294696 645866 294748 645872
rect 307392 645924 307444 645930
rect 307392 645866 307444 645872
rect 188434 645008 188490 645017
rect 188434 644943 188490 644952
rect 188448 545018 188476 644943
rect 291844 644496 291896 644502
rect 291844 644438 291896 644444
rect 188526 643240 188582 643249
rect 188526 643175 188582 643184
rect 188436 545012 188488 545018
rect 188436 544954 188488 544960
rect 188540 544882 188568 643175
rect 290464 643136 290516 643142
rect 290464 643078 290516 643084
rect 188618 642016 188674 642025
rect 188618 641951 188674 641960
rect 188528 544876 188580 544882
rect 188528 544818 188580 544824
rect 188632 544814 188660 641951
rect 287704 641776 287756 641782
rect 287704 641718 287756 641724
rect 188710 640384 188766 640393
rect 188710 640319 188766 640328
rect 286324 640348 286376 640354
rect 188620 544808 188672 544814
rect 188620 544750 188672 544756
rect 188724 544678 188752 640319
rect 286324 640290 286376 640296
rect 188802 639296 188858 639305
rect 188802 639231 188858 639240
rect 188712 544672 188764 544678
rect 188712 544614 188764 544620
rect 188816 544542 188844 639231
rect 284944 638988 284996 638994
rect 284944 638930 284996 638936
rect 188894 637664 188950 637673
rect 188894 637599 188950 637608
rect 188804 544536 188856 544542
rect 188804 544478 188856 544484
rect 188908 544474 188936 637599
rect 282182 587208 282238 587217
rect 282182 587143 282238 587152
rect 282196 586537 282224 587143
rect 282182 586528 282238 586537
rect 282182 586463 282238 586472
rect 188986 579728 189042 579737
rect 188986 579663 189042 579672
rect 188896 544468 188948 544474
rect 188896 544410 188948 544416
rect 179236 543254 179288 543260
rect 188342 543280 188398 543289
rect 177212 542700 177264 542706
rect 177212 542642 177264 542648
rect 177224 539988 177252 542642
rect 179248 539988 179276 543254
rect 188342 543215 188398 543224
rect 183376 543176 183428 543182
rect 183376 543118 183428 543124
rect 181352 542632 181404 542638
rect 181352 542574 181404 542580
rect 181364 539988 181392 542574
rect 183388 539988 183416 543118
rect 187516 543108 187568 543114
rect 187516 543050 187568 543056
rect 185492 542768 185544 542774
rect 185492 542710 185544 542716
rect 185504 539988 185532 542710
rect 187528 539988 187556 543050
rect 189000 543017 189028 579663
rect 282196 578950 282224 586463
rect 282184 578944 282236 578950
rect 282184 578886 282236 578892
rect 229374 560008 229430 560017
rect 229374 559943 229430 559952
rect 225970 559872 226026 559881
rect 225970 559807 226026 559816
rect 194414 558920 194470 558929
rect 194414 558855 194470 558864
rect 195978 558920 196034 558929
rect 195978 558855 196034 558864
rect 200210 558920 200266 558929
rect 200210 558855 200212 558864
rect 194428 558278 194456 558855
rect 194416 558272 194468 558278
rect 194416 558214 194468 558220
rect 194428 558113 194456 558214
rect 194414 558104 194470 558113
rect 194414 558039 194470 558048
rect 189632 545080 189684 545086
rect 189632 545022 189684 545028
rect 188986 543008 189042 543017
rect 188986 542943 189042 542952
rect 189644 539988 189672 545022
rect 195992 544406 196020 558855
rect 200264 558855 200266 558864
rect 201498 558920 201554 558929
rect 201498 558855 201554 558864
rect 202786 558920 202842 558929
rect 202786 558855 202842 558864
rect 203798 558920 203854 558929
rect 203798 558855 203854 558864
rect 204166 558920 204222 558929
rect 204166 558855 204222 558864
rect 205546 558920 205602 558929
rect 205546 558855 205602 558864
rect 206374 558920 206430 558929
rect 206374 558855 206430 558864
rect 208490 558920 208546 558929
rect 208490 558855 208546 558864
rect 211894 558920 211950 558929
rect 211894 558855 211950 558864
rect 213090 558920 213146 558929
rect 213090 558855 213146 558864
rect 213918 558920 213974 558929
rect 213918 558855 213974 558864
rect 215298 558920 215354 558929
rect 215298 558855 215354 558864
rect 218794 558920 218850 558929
rect 218794 558855 218850 558864
rect 220082 558920 220138 558929
rect 220082 558855 220138 558864
rect 221094 558920 221150 558929
rect 221094 558855 221150 558864
rect 222290 558920 222346 558929
rect 222290 558855 222346 558864
rect 223578 558920 223634 558929
rect 223578 558855 223634 558864
rect 223946 558920 224002 558929
rect 223946 558855 224002 558864
rect 200212 558826 200264 558832
rect 201512 558822 201540 558855
rect 201500 558816 201552 558822
rect 201500 558758 201552 558764
rect 202142 558784 202198 558793
rect 202142 558719 202198 558728
rect 202156 557938 202184 558719
rect 202144 557932 202196 557938
rect 202144 557874 202196 557880
rect 197912 544944 197964 544950
rect 197912 544886 197964 544892
rect 195980 544400 196032 544406
rect 195980 544342 196032 544348
rect 193772 543040 193824 543046
rect 193772 542982 193824 542988
rect 191748 542836 191800 542842
rect 191748 542778 191800 542784
rect 191760 539988 191788 542778
rect 193784 539988 193812 542982
rect 195888 542904 195940 542910
rect 195888 542846 195940 542852
rect 195900 539988 195928 542846
rect 197924 539988 197952 544886
rect 200026 543688 200082 543697
rect 200026 543623 200082 543632
rect 200040 539988 200068 543623
rect 202156 543250 202184 557874
rect 202144 543244 202196 543250
rect 202144 543186 202196 543192
rect 202800 543182 202828 558855
rect 203812 558210 203840 558855
rect 203800 558204 203852 558210
rect 203800 558146 203852 558152
rect 203812 557734 203840 558146
rect 203800 557728 203852 557734
rect 203800 557670 203852 557676
rect 202788 543176 202840 543182
rect 202050 543144 202106 543153
rect 202788 543118 202840 543124
rect 204180 543114 204208 558855
rect 204902 558648 204958 558657
rect 204902 558583 204958 558592
rect 204916 557734 204944 558583
rect 204904 557728 204956 557734
rect 204904 557670 204956 557676
rect 204916 543386 204944 557670
rect 205560 543726 205588 558855
rect 206388 558346 206416 558855
rect 208504 558754 208532 558855
rect 208492 558748 208544 558754
rect 208492 558690 208544 558696
rect 211160 558748 211212 558754
rect 211160 558690 211212 558696
rect 206376 558340 206428 558346
rect 206376 558282 206428 558288
rect 206388 557802 206416 558282
rect 208504 557870 208532 558690
rect 211172 558657 211200 558690
rect 210514 558648 210570 558657
rect 210514 558583 210570 558592
rect 211158 558648 211214 558657
rect 211158 558583 211214 558592
rect 208492 557864 208544 557870
rect 208492 557806 208544 557812
rect 206376 557796 206428 557802
rect 206376 557738 206428 557744
rect 207664 557796 207716 557802
rect 207664 557738 207716 557744
rect 207676 557705 207704 557738
rect 207662 557696 207718 557705
rect 207662 557631 207718 557640
rect 209042 557696 209098 557705
rect 210528 557666 210556 558583
rect 211908 558414 211936 558855
rect 213104 558618 213132 558855
rect 212540 558612 212592 558618
rect 212540 558554 212592 558560
rect 213092 558612 213144 558618
rect 213092 558554 213144 558560
rect 211160 558408 211212 558414
rect 211160 558350 211212 558356
rect 211896 558408 211948 558414
rect 211896 558350 211948 558356
rect 211172 557938 211200 558350
rect 212552 558210 212580 558554
rect 212540 558204 212592 558210
rect 212540 558146 212592 558152
rect 213932 558142 213960 558855
rect 215312 558346 215340 558855
rect 217966 558784 218022 558793
rect 217966 558719 217968 558728
rect 218020 558719 218022 558728
rect 217968 558690 218020 558696
rect 215300 558340 215352 558346
rect 215300 558282 215352 558288
rect 213920 558136 213972 558142
rect 213920 558078 213972 558084
rect 211160 557932 211212 557938
rect 211160 557874 211212 557880
rect 213932 557734 213960 558078
rect 217980 557802 218008 558690
rect 218808 558550 218836 558855
rect 220096 558822 220124 558855
rect 220084 558816 220136 558822
rect 220084 558758 220136 558764
rect 218796 558544 218848 558550
rect 218796 558486 218848 558492
rect 217968 557796 218020 557802
rect 217968 557738 218020 557744
rect 213920 557728 213972 557734
rect 210974 557696 211030 557705
rect 209042 557631 209098 557640
rect 210516 557660 210568 557666
rect 206926 557560 206982 557569
rect 206926 557495 206982 557504
rect 206192 544740 206244 544746
rect 206192 544682 206244 544688
rect 205548 543720 205600 543726
rect 205548 543662 205600 543668
rect 204904 543380 204956 543386
rect 204904 543322 204956 543328
rect 202050 543079 202106 543088
rect 204168 543108 204220 543114
rect 202064 539988 202092 543079
rect 204168 543050 204220 543056
rect 204168 542972 204220 542978
rect 204168 542914 204220 542920
rect 204180 539988 204208 542914
rect 206204 539988 206232 544682
rect 206940 543658 206968 557495
rect 206928 543652 206980 543658
rect 206928 543594 206980 543600
rect 207676 543454 207704 557631
rect 209056 557598 209084 557631
rect 213920 557670 213972 557676
rect 217874 557696 217930 557705
rect 210974 557631 211030 557640
rect 217874 557631 217930 557640
rect 210516 557602 210568 557608
rect 209044 557592 209096 557598
rect 208306 557560 208362 557569
rect 209044 557534 209096 557540
rect 209686 557560 209742 557569
rect 208306 557495 208362 557504
rect 208320 543590 208348 557495
rect 208308 543584 208360 543590
rect 208308 543526 208360 543532
rect 209056 543522 209084 557534
rect 209686 557495 209742 557504
rect 209700 543522 209728 557495
rect 210422 543552 210478 543561
rect 209044 543516 209096 543522
rect 209044 543458 209096 543464
rect 209688 543516 209740 543522
rect 210422 543487 210478 543496
rect 209688 543458 209740 543464
rect 207664 543448 207716 543454
rect 207664 543390 207716 543396
rect 208306 543416 208362 543425
rect 208306 543351 208362 543360
rect 208320 539988 208348 543351
rect 210436 539988 210464 543487
rect 210988 543454 211016 557631
rect 211066 557560 211122 557569
rect 211066 557495 211122 557504
rect 212446 557560 212502 557569
rect 212446 557495 212502 557504
rect 213826 557560 213882 557569
rect 213826 557495 213882 557504
rect 215206 557560 215262 557569
rect 215206 557495 215262 557504
rect 216586 557560 216642 557569
rect 216586 557495 216642 557504
rect 210976 543448 211028 543454
rect 210976 543390 211028 543396
rect 211080 543250 211108 557495
rect 212460 545578 212488 557495
rect 212368 545550 212488 545578
rect 212368 543386 212396 545550
rect 212448 544604 212500 544610
rect 212448 544546 212500 544552
rect 212356 543380 212408 543386
rect 212356 543322 212408 543328
rect 211068 543244 211120 543250
rect 211068 543186 211120 543192
rect 212460 539988 212488 544546
rect 213840 543114 213868 557495
rect 215220 543318 215248 557495
rect 215208 543312 215260 543318
rect 215208 543254 215260 543260
rect 216600 543182 216628 557495
rect 214564 543176 214616 543182
rect 214564 543118 214616 543124
rect 216588 543176 216640 543182
rect 216588 543118 216640 543124
rect 213828 543108 213880 543114
rect 213828 543050 213880 543056
rect 214576 539988 214604 543118
rect 217888 543046 217916 557631
rect 218808 557598 218836 558486
rect 220096 557666 220124 558758
rect 220728 558680 220780 558686
rect 220726 558648 220728 558657
rect 220780 558648 220782 558657
rect 220726 558583 220782 558592
rect 221108 558414 221136 558855
rect 222304 558618 222332 558855
rect 222292 558612 222344 558618
rect 222292 558554 222344 558560
rect 221096 558408 221148 558414
rect 221096 558350 221148 558356
rect 223592 558006 223620 558855
rect 223960 558346 223988 558855
rect 225984 558754 226012 559807
rect 227258 559328 227314 559337
rect 227258 559263 227314 559272
rect 225972 558748 226024 558754
rect 225972 558690 226024 558696
rect 227272 558686 227300 559263
rect 228086 558920 228142 558929
rect 228086 558855 228142 558864
rect 227260 558680 227312 558686
rect 227260 558622 227312 558628
rect 228100 558550 228128 558855
rect 229388 558822 229416 559943
rect 235906 558920 235962 558929
rect 235906 558855 235962 558864
rect 237286 558920 237342 558929
rect 237286 558855 237342 558864
rect 240046 558920 240102 558929
rect 240046 558855 240102 558864
rect 282092 558884 282144 558890
rect 229376 558816 229428 558822
rect 229376 558758 229428 558764
rect 231950 558784 232006 558793
rect 231950 558719 232006 558728
rect 233238 558784 233294 558793
rect 233238 558719 233294 558728
rect 234618 558784 234674 558793
rect 234618 558719 234620 558728
rect 231858 558648 231914 558657
rect 231858 558583 231860 558592
rect 231912 558583 231914 558592
rect 231860 558554 231912 558560
rect 228088 558544 228140 558550
rect 228088 558486 228140 558492
rect 230478 558512 230534 558521
rect 230478 558447 230534 558456
rect 230492 558414 230520 558447
rect 230480 558408 230532 558414
rect 230480 558350 230532 558356
rect 223948 558340 224000 558346
rect 223948 558282 224000 558288
rect 231964 558210 231992 558719
rect 233252 558346 233280 558719
rect 234672 558719 234674 558728
rect 234620 558690 234672 558696
rect 233240 558340 233292 558346
rect 233240 558282 233292 558288
rect 231952 558204 232004 558210
rect 231952 558146 232004 558152
rect 223580 558000 223632 558006
rect 223580 557942 223632 557948
rect 226246 557696 226302 557705
rect 220084 557660 220136 557666
rect 226246 557631 226302 557640
rect 233146 557696 233202 557705
rect 233146 557631 233202 557640
rect 220084 557602 220136 557608
rect 218796 557592 218848 557598
rect 217966 557560 218022 557569
rect 218796 557534 218848 557540
rect 219346 557560 219402 557569
rect 217966 557495 218022 557504
rect 219346 557495 219402 557504
rect 220726 557560 220782 557569
rect 220726 557495 220782 557504
rect 222106 557560 222162 557569
rect 222106 557495 222162 557504
rect 223486 557560 223542 557569
rect 223486 557495 223542 557504
rect 224866 557560 224922 557569
rect 224866 557495 224922 557504
rect 226154 557560 226210 557569
rect 226154 557495 226210 557504
rect 216588 543040 216640 543046
rect 216588 542982 216640 542988
rect 217876 543040 217928 543046
rect 217876 542982 217928 542988
rect 216600 539988 216628 542982
rect 217980 542570 218008 557495
rect 218704 543720 218756 543726
rect 218704 543662 218756 543668
rect 217968 542564 218020 542570
rect 217968 542506 218020 542512
rect 218716 539988 218744 543662
rect 219360 542502 219388 557495
rect 220740 543794 220768 557495
rect 220728 543788 220780 543794
rect 220728 543730 220780 543736
rect 220544 543720 220596 543726
rect 220544 543662 220596 543668
rect 220556 542638 220584 543662
rect 220728 543652 220780 543658
rect 220728 543594 220780 543600
rect 220544 542632 220596 542638
rect 220544 542574 220596 542580
rect 219348 542496 219400 542502
rect 219348 542438 219400 542444
rect 220740 539988 220768 543594
rect 222120 542706 222148 557495
rect 222844 543584 222896 543590
rect 222844 543526 222896 543532
rect 222108 542700 222160 542706
rect 222108 542642 222160 542648
rect 222856 539988 222884 543526
rect 223500 542842 223528 557495
rect 224880 545306 224908 557495
rect 224696 545278 224908 545306
rect 223488 542836 223540 542842
rect 223488 542778 223540 542784
rect 224696 542774 224724 545278
rect 224868 543516 224920 543522
rect 224868 543458 224920 543464
rect 224684 542768 224736 542774
rect 224684 542710 224736 542716
rect 224880 539988 224908 543458
rect 226168 542978 226196 557495
rect 226156 542972 226208 542978
rect 226156 542914 226208 542920
rect 226260 542910 226288 557631
rect 227626 557560 227682 557569
rect 227626 557495 227682 557504
rect 229006 557560 229062 557569
rect 229006 557495 229062 557504
rect 230386 557560 230442 557569
rect 230386 557495 230442 557504
rect 231766 557560 231822 557569
rect 231766 557495 231822 557504
rect 233054 557560 233110 557569
rect 233054 557495 233110 557504
rect 227640 543726 227668 557495
rect 227628 543720 227680 543726
rect 227628 543662 227680 543668
rect 229020 543658 229048 557495
rect 229008 543652 229060 543658
rect 229008 543594 229060 543600
rect 230400 543590 230428 557495
rect 230388 543584 230440 543590
rect 230388 543526 230440 543532
rect 231780 543522 231808 557495
rect 231768 543516 231820 543522
rect 231768 543458 231820 543464
rect 226984 543448 227036 543454
rect 226984 543390 227036 543396
rect 226248 542904 226300 542910
rect 226248 542846 226300 542852
rect 226996 539988 227024 543390
rect 233068 543386 233096 557495
rect 233160 543454 233188 557631
rect 234526 557560 234582 557569
rect 234526 557495 234582 557504
rect 233148 543448 233200 543454
rect 233148 543390 233200 543396
rect 231124 543380 231176 543386
rect 231124 543322 231176 543328
rect 233056 543380 233108 543386
rect 233056 543322 233108 543328
rect 229100 543244 229152 543250
rect 229100 543186 229152 543192
rect 229112 539988 229140 543186
rect 231136 539988 231164 543322
rect 234540 543250 234568 557495
rect 235920 543318 235948 558855
rect 235998 558784 236054 558793
rect 235998 558719 236054 558728
rect 236012 558686 236040 558719
rect 236000 558680 236052 558686
rect 236000 558622 236052 558628
rect 235264 543312 235316 543318
rect 235264 543254 235316 543260
rect 235908 543312 235960 543318
rect 235908 543254 235960 543260
rect 234528 543244 234580 543250
rect 234528 543186 234580 543192
rect 233240 543108 233292 543114
rect 233240 543050 233292 543056
rect 233252 539988 233280 543050
rect 235276 539988 235304 543254
rect 237300 543114 237328 558855
rect 237378 558648 237434 558657
rect 237378 558583 237434 558592
rect 237392 558550 237420 558583
rect 237380 558544 237432 558550
rect 237380 558486 237432 558492
rect 238758 558376 238814 558385
rect 238758 558311 238760 558320
rect 238812 558311 238814 558320
rect 238760 558282 238812 558288
rect 238666 558104 238722 558113
rect 238666 558039 238722 558048
rect 238680 543182 238708 558039
rect 237380 543176 237432 543182
rect 237380 543118 237432 543124
rect 238668 543176 238720 543182
rect 238668 543118 238720 543124
rect 237288 543108 237340 543114
rect 237288 543050 237340 543056
rect 237392 539988 237420 543118
rect 240060 543046 240088 558855
rect 282092 558826 282144 558832
rect 281908 558476 281960 558482
rect 281908 558418 281960 558424
rect 281816 558340 281868 558346
rect 281816 558282 281868 558288
rect 258080 543720 258132 543726
rect 258080 543662 258132 543668
rect 239404 543040 239456 543046
rect 239404 542982 239456 542988
rect 240048 543040 240100 543046
rect 240048 542982 240100 542988
rect 239416 539988 239444 542982
rect 256056 542972 256108 542978
rect 256056 542914 256108 542920
rect 253940 542904 253992 542910
rect 253940 542846 253992 542852
rect 249800 542836 249852 542842
rect 249800 542778 249852 542784
rect 247776 542700 247828 542706
rect 247776 542642 247828 542648
rect 245660 542632 245712 542638
rect 245660 542574 245712 542580
rect 241520 542564 241572 542570
rect 241520 542506 241572 542512
rect 241532 539988 241560 542506
rect 243544 542496 243596 542502
rect 243544 542438 243596 542444
rect 243556 539988 243584 542438
rect 245672 539988 245700 542574
rect 247788 539988 247816 542642
rect 249812 539988 249840 542778
rect 251916 542768 251968 542774
rect 251916 542710 251968 542716
rect 251928 539988 251956 542710
rect 253952 539988 253980 542846
rect 256068 539988 256096 542914
rect 258092 539988 258120 543662
rect 260196 543652 260248 543658
rect 260196 543594 260248 543600
rect 260208 539988 260236 543594
rect 262220 543584 262272 543590
rect 262220 543526 262272 543532
rect 262232 539988 262260 543526
rect 264336 543516 264388 543522
rect 264336 543458 264388 543464
rect 264348 539988 264376 543458
rect 266452 543448 266504 543454
rect 266452 543390 266504 543396
rect 266464 539988 266492 543390
rect 268476 543380 268528 543386
rect 268476 543322 268528 543328
rect 268488 539988 268516 543322
rect 272616 543312 272668 543318
rect 272616 543254 272668 543260
rect 270592 543244 270644 543250
rect 270592 543186 270644 543192
rect 270604 539988 270632 543186
rect 272628 539988 272656 543254
rect 276756 543176 276808 543182
rect 276756 543118 276808 543124
rect 274732 543108 274784 543114
rect 274732 543050 274784 543056
rect 274744 539988 274772 543050
rect 276768 539988 276796 543118
rect 278872 543040 278924 543046
rect 278872 542982 278924 542988
rect 278884 539988 278912 542982
rect 281724 539572 281776 539578
rect 281724 539514 281776 539520
rect 281736 539073 281764 539514
rect 281722 539064 281778 539073
rect 281722 538999 281778 539008
rect 281724 538212 281776 538218
rect 281724 538154 281776 538160
rect 281736 537033 281764 538154
rect 281722 537024 281778 537033
rect 281722 536959 281778 536968
rect 281724 535424 281776 535430
rect 281724 535366 281776 535372
rect 281736 534993 281764 535366
rect 281722 534984 281778 534993
rect 281722 534919 281778 534928
rect 281724 534064 281776 534070
rect 281724 534006 281776 534012
rect 281736 532953 281764 534006
rect 281722 532944 281778 532953
rect 281722 532879 281778 532888
rect 281724 531276 281776 531282
rect 281724 531218 281776 531224
rect 281736 530913 281764 531218
rect 281722 530904 281778 530913
rect 281722 530839 281778 530848
rect 281724 529916 281776 529922
rect 281724 529858 281776 529864
rect 281736 528873 281764 529858
rect 281722 528864 281778 528873
rect 281722 528799 281778 528808
rect 281724 527128 281776 527134
rect 281724 527070 281776 527076
rect 281736 526833 281764 527070
rect 281722 526824 281778 526833
rect 281722 526759 281778 526768
rect 281724 525768 281776 525774
rect 281724 525710 281776 525716
rect 281736 524793 281764 525710
rect 281722 524784 281778 524793
rect 281722 524719 281778 524728
rect 281724 522980 281776 522986
rect 281724 522922 281776 522928
rect 281736 522753 281764 522922
rect 281722 522744 281778 522753
rect 281722 522679 281778 522688
rect 281724 521620 281776 521626
rect 281724 521562 281776 521568
rect 281736 520713 281764 521562
rect 281722 520704 281778 520713
rect 281722 520639 281778 520648
rect 281724 518900 281776 518906
rect 281724 518842 281776 518848
rect 281736 518673 281764 518842
rect 281722 518664 281778 518673
rect 281722 518599 281778 518608
rect 281724 517472 281776 517478
rect 281724 517414 281776 517420
rect 281736 516633 281764 517414
rect 281722 516624 281778 516633
rect 281722 516559 281778 516568
rect 281724 514752 281776 514758
rect 281724 514694 281776 514700
rect 281736 514593 281764 514694
rect 281722 514584 281778 514593
rect 281722 514519 281778 514528
rect 281724 513324 281776 513330
rect 281724 513266 281776 513272
rect 281736 512553 281764 513266
rect 281722 512544 281778 512553
rect 281722 512479 281778 512488
rect 281724 510604 281776 510610
rect 281724 510546 281776 510552
rect 281736 510513 281764 510546
rect 281722 510504 281778 510513
rect 281722 510439 281778 510448
rect 281724 509244 281776 509250
rect 281724 509186 281776 509192
rect 281736 508473 281764 509186
rect 281722 508464 281778 508473
rect 281722 508399 281778 508408
rect 281724 506456 281776 506462
rect 281722 506424 281724 506433
rect 281776 506424 281778 506433
rect 281722 506359 281778 506368
rect 281724 505096 281776 505102
rect 281724 505038 281776 505044
rect 281736 504393 281764 505038
rect 281722 504384 281778 504393
rect 281722 504319 281778 504328
rect 281722 502344 281778 502353
rect 281722 502279 281724 502288
rect 281776 502279 281778 502288
rect 281724 502250 281776 502256
rect 281724 500948 281776 500954
rect 281724 500890 281776 500896
rect 281736 500313 281764 500890
rect 281722 500304 281778 500313
rect 281722 500239 281778 500248
rect 281724 499520 281776 499526
rect 281724 499462 281776 499468
rect 281736 498273 281764 499462
rect 281722 498264 281778 498273
rect 281722 498199 281778 498208
rect 281724 496800 281776 496806
rect 281724 496742 281776 496748
rect 281736 496233 281764 496742
rect 281722 496224 281778 496233
rect 281722 496159 281778 496168
rect 281724 495440 281776 495446
rect 281724 495382 281776 495388
rect 281736 494193 281764 495382
rect 281722 494184 281778 494193
rect 281722 494119 281778 494128
rect 281724 492652 281776 492658
rect 281724 492594 281776 492600
rect 281736 492153 281764 492594
rect 281722 492144 281778 492153
rect 281722 492079 281778 492088
rect 281724 491292 281776 491298
rect 281724 491234 281776 491240
rect 281736 490113 281764 491234
rect 281722 490104 281778 490113
rect 281722 490039 281778 490048
rect 281724 488504 281776 488510
rect 281724 488446 281776 488452
rect 281736 488073 281764 488446
rect 281722 488064 281778 488073
rect 281722 487999 281778 488008
rect 281724 487144 281776 487150
rect 281724 487086 281776 487092
rect 281736 486033 281764 487086
rect 281722 486024 281778 486033
rect 281722 485959 281778 485968
rect 281724 484356 281776 484362
rect 281724 484298 281776 484304
rect 281736 483993 281764 484298
rect 281722 483984 281778 483993
rect 281722 483919 281778 483928
rect 281724 482996 281776 483002
rect 281724 482938 281776 482944
rect 281736 481953 281764 482938
rect 281722 481944 281778 481953
rect 281722 481879 281778 481888
rect 281724 480208 281776 480214
rect 281724 480150 281776 480156
rect 281736 479913 281764 480150
rect 281722 479904 281778 479913
rect 281722 479839 281778 479848
rect 281724 478848 281776 478854
rect 281724 478790 281776 478796
rect 281736 477873 281764 478790
rect 281722 477864 281778 477873
rect 281722 477799 281778 477808
rect 281724 476060 281776 476066
rect 281724 476002 281776 476008
rect 281736 475833 281764 476002
rect 281722 475824 281778 475833
rect 281722 475759 281778 475768
rect 281724 474700 281776 474706
rect 281724 474642 281776 474648
rect 281736 473793 281764 474642
rect 281722 473784 281778 473793
rect 281722 473719 281778 473728
rect 281724 471980 281776 471986
rect 281724 471922 281776 471928
rect 281736 471753 281764 471922
rect 281722 471744 281778 471753
rect 281722 471679 281778 471688
rect 281724 470552 281776 470558
rect 281724 470494 281776 470500
rect 281736 469713 281764 470494
rect 281722 469704 281778 469713
rect 281722 469639 281778 469648
rect 281724 467832 281776 467838
rect 281724 467774 281776 467780
rect 281736 467673 281764 467774
rect 281722 467664 281778 467673
rect 281722 467599 281778 467608
rect 281724 466404 281776 466410
rect 281724 466346 281776 466352
rect 281736 465633 281764 466346
rect 281722 465624 281778 465633
rect 281722 465559 281778 465568
rect 281724 463684 281776 463690
rect 281724 463626 281776 463632
rect 281736 463593 281764 463626
rect 281722 463584 281778 463593
rect 281722 463519 281778 463528
rect 281724 462324 281776 462330
rect 281724 462266 281776 462272
rect 281736 461553 281764 462266
rect 281722 461544 281778 461553
rect 281722 461479 281778 461488
rect 281724 459536 281776 459542
rect 281722 459504 281724 459513
rect 281776 459504 281778 459513
rect 281722 459439 281778 459448
rect 281724 458176 281776 458182
rect 281724 458118 281776 458124
rect 281736 457473 281764 458118
rect 281722 457464 281778 457473
rect 281722 457399 281778 457408
rect 281722 455424 281778 455433
rect 281722 455359 281724 455368
rect 281776 455359 281778 455368
rect 281724 455330 281776 455336
rect 281724 454028 281776 454034
rect 281724 453970 281776 453976
rect 281736 453393 281764 453970
rect 281722 453384 281778 453393
rect 281722 453319 281778 453328
rect 281724 452600 281776 452606
rect 281724 452542 281776 452548
rect 281736 451353 281764 452542
rect 281722 451344 281778 451353
rect 281722 451279 281778 451288
rect 281724 449880 281776 449886
rect 281724 449822 281776 449828
rect 281736 449313 281764 449822
rect 281722 449304 281778 449313
rect 281722 449239 281778 449248
rect 281724 448520 281776 448526
rect 281724 448462 281776 448468
rect 281736 447273 281764 448462
rect 281722 447264 281778 447273
rect 281722 447199 281778 447208
rect 281724 445732 281776 445738
rect 281724 445674 281776 445680
rect 281736 445233 281764 445674
rect 281722 445224 281778 445233
rect 281722 445159 281778 445168
rect 281724 444372 281776 444378
rect 281724 444314 281776 444320
rect 281736 443193 281764 444314
rect 281722 443184 281778 443193
rect 281722 443119 281778 443128
rect 281724 441584 281776 441590
rect 281724 441526 281776 441532
rect 281736 441153 281764 441526
rect 281722 441144 281778 441153
rect 281722 441079 281778 441088
rect 281724 440224 281776 440230
rect 281724 440166 281776 440172
rect 281736 439113 281764 440166
rect 281722 439104 281778 439113
rect 281722 439039 281778 439048
rect 281724 437436 281776 437442
rect 281724 437378 281776 437384
rect 281736 437073 281764 437378
rect 281722 437064 281778 437073
rect 281722 436999 281778 437008
rect 281724 436076 281776 436082
rect 281724 436018 281776 436024
rect 281736 435033 281764 436018
rect 281722 435024 281778 435033
rect 281722 434959 281778 434968
rect 281724 433288 281776 433294
rect 281724 433230 281776 433236
rect 281736 432993 281764 433230
rect 281722 432984 281778 432993
rect 281722 432919 281778 432928
rect 281724 431928 281776 431934
rect 281724 431870 281776 431876
rect 281736 431089 281764 431870
rect 281722 431080 281778 431089
rect 281722 431015 281778 431024
rect 281724 429140 281776 429146
rect 281724 429082 281776 429088
rect 281736 429049 281764 429082
rect 281722 429040 281778 429049
rect 281722 428975 281778 428984
rect 281724 427780 281776 427786
rect 281724 427722 281776 427728
rect 281736 427009 281764 427722
rect 281722 427000 281778 427009
rect 281722 426935 281778 426944
rect 281724 425060 281776 425066
rect 281724 425002 281776 425008
rect 281736 424969 281764 425002
rect 281722 424960 281778 424969
rect 281722 424895 281778 424904
rect 281724 423632 281776 423638
rect 281724 423574 281776 423580
rect 281736 422929 281764 423574
rect 281722 422920 281778 422929
rect 281722 422855 281778 422864
rect 281724 420912 281776 420918
rect 281722 420880 281724 420889
rect 281776 420880 281778 420889
rect 281722 420815 281778 420824
rect 281724 419484 281776 419490
rect 281724 419426 281776 419432
rect 281736 418849 281764 419426
rect 281722 418840 281778 418849
rect 281722 418775 281778 418784
rect 281724 418124 281776 418130
rect 281724 418066 281776 418072
rect 281736 416809 281764 418066
rect 281722 416800 281778 416809
rect 281722 416735 281778 416744
rect 281724 415404 281776 415410
rect 281724 415346 281776 415352
rect 281736 414769 281764 415346
rect 281722 414760 281778 414769
rect 281722 414695 281778 414704
rect 281724 413976 281776 413982
rect 281724 413918 281776 413924
rect 281736 412729 281764 413918
rect 281722 412720 281778 412729
rect 281722 412655 281778 412664
rect 281632 412412 281684 412418
rect 281632 412354 281684 412360
rect 281540 412344 281592 412350
rect 281540 412286 281592 412292
rect 281552 404274 281580 412286
rect 281644 404410 281672 412354
rect 281724 411392 281776 411398
rect 281724 411334 281776 411340
rect 281736 404569 281764 411334
rect 281828 408649 281856 558282
rect 281814 408640 281870 408649
rect 281814 408575 281870 408584
rect 281920 406609 281948 558418
rect 282000 558408 282052 558414
rect 282000 558350 282052 558356
rect 282012 411398 282040 558350
rect 282000 411392 282052 411398
rect 282000 411334 282052 411340
rect 282000 411256 282052 411262
rect 282000 411198 282052 411204
rect 282012 410689 282040 411198
rect 281998 410680 282054 410689
rect 281998 410615 282054 410624
rect 282000 410576 282052 410582
rect 282000 410518 282052 410524
rect 281906 406600 281962 406609
rect 281906 406535 281962 406544
rect 281722 404560 281778 404569
rect 281722 404495 281778 404504
rect 281644 404382 281764 404410
rect 281552 404246 281672 404274
rect 281540 404184 281592 404190
rect 281540 404126 281592 404132
rect 281552 402529 281580 404126
rect 281538 402520 281594 402529
rect 281538 402455 281594 402464
rect 281644 400489 281672 404246
rect 281630 400480 281686 400489
rect 281630 400415 281686 400424
rect 281736 398449 281764 404382
rect 282012 404190 282040 410518
rect 282000 404184 282052 404190
rect 282000 404126 282052 404132
rect 281722 398440 281778 398449
rect 281722 398375 281778 398384
rect 281540 397112 281592 397118
rect 281540 397054 281592 397060
rect 281552 396409 281580 397054
rect 281538 396400 281594 396409
rect 281538 396335 281594 396344
rect 282104 394369 282132 558826
rect 282090 394360 282146 394369
rect 282090 394295 282146 394304
rect 281908 378072 281960 378078
rect 281906 378040 281908 378049
rect 281960 378040 281962 378049
rect 281906 377975 281962 377984
rect 281724 365832 281776 365838
rect 281722 365800 281724 365809
rect 281776 365800 281778 365809
rect 281722 365735 281778 365744
rect 281908 362908 281960 362914
rect 281908 362850 281960 362856
rect 281920 361729 281948 362850
rect 281906 361720 281962 361729
rect 281906 361655 281962 361664
rect 281908 360188 281960 360194
rect 281908 360130 281960 360136
rect 281920 359689 281948 360130
rect 281906 359680 281962 359689
rect 281906 359615 281962 359624
rect 281724 357672 281776 357678
rect 281722 357640 281724 357649
rect 281776 357640 281778 357649
rect 281722 357575 281778 357584
rect 282092 355904 282144 355910
rect 282092 355846 282144 355852
rect 282104 355609 282132 355846
rect 282090 355600 282146 355609
rect 282090 355535 282146 355544
rect 281540 346112 281592 346118
rect 281540 346054 281592 346060
rect 281552 345409 281580 346054
rect 281538 345400 281594 345409
rect 281538 345335 281594 345344
rect 281540 341352 281592 341358
rect 281538 341320 281540 341329
rect 281592 341320 281594 341329
rect 281538 341255 281594 341264
rect 281724 339312 281776 339318
rect 281722 339280 281724 339289
rect 281776 339280 281778 339289
rect 281722 339215 281778 339224
rect 281540 337612 281592 337618
rect 281540 337554 281592 337560
rect 281552 337249 281580 337554
rect 281538 337240 281594 337249
rect 281538 337175 281594 337184
rect 281632 335232 281684 335238
rect 281630 335200 281632 335209
rect 281684 335200 281686 335209
rect 281630 335135 281686 335144
rect 281540 333260 281592 333266
rect 281540 333202 281592 333208
rect 281552 333169 281580 333202
rect 281538 333160 281594 333169
rect 281538 333095 281594 333104
rect 281540 331152 281592 331158
rect 281538 331120 281540 331129
rect 281592 331120 281594 331129
rect 281538 331055 281594 331064
rect 281540 329112 281592 329118
rect 281538 329080 281540 329089
rect 281592 329080 281594 329089
rect 281538 329015 281594 329024
rect 281540 327072 281592 327078
rect 281538 327040 281540 327049
rect 281592 327040 281594 327049
rect 281538 326975 281594 326984
rect 281540 325100 281592 325106
rect 281540 325042 281592 325048
rect 281552 325009 281580 325042
rect 281538 325000 281594 325009
rect 281538 324935 281594 324944
rect 282196 321065 282224 578886
rect 283932 558884 283984 558890
rect 283932 558826 283984 558832
rect 283654 558240 283710 558249
rect 283564 558204 283616 558210
rect 283654 558175 283710 558184
rect 283564 558146 283616 558152
rect 282276 558000 282328 558006
rect 282276 557942 282328 557948
rect 282288 380089 282316 557942
rect 282368 557932 282420 557938
rect 282368 557874 282420 557880
rect 282380 382129 282408 557874
rect 282460 557864 282512 557870
rect 282460 557806 282512 557812
rect 282472 384169 282500 557806
rect 282552 557796 282604 557802
rect 282552 557738 282604 557744
rect 282564 386209 282592 557738
rect 282644 557728 282696 557734
rect 282644 557670 282696 557676
rect 282656 388249 282684 557670
rect 282736 557660 282788 557666
rect 282736 557602 282788 557608
rect 282748 390289 282776 557602
rect 282828 557592 282880 557598
rect 282828 557534 282880 557540
rect 282840 392329 282868 557534
rect 283472 557524 283524 557530
rect 283472 557466 283524 557472
rect 283104 412208 283156 412214
rect 283104 412150 283156 412156
rect 283012 412140 283064 412146
rect 283012 412082 283064 412088
rect 282920 410576 282972 410582
rect 282920 410518 282972 410524
rect 282826 392320 282882 392329
rect 282826 392255 282882 392264
rect 282734 390280 282790 390289
rect 282734 390215 282790 390224
rect 282642 388240 282698 388249
rect 282642 388175 282698 388184
rect 282550 386200 282606 386209
rect 282550 386135 282606 386144
rect 282458 384160 282514 384169
rect 282458 384095 282514 384104
rect 282366 382120 282422 382129
rect 282366 382055 282422 382064
rect 282274 380080 282330 380089
rect 282274 380015 282330 380024
rect 282828 376712 282880 376718
rect 282828 376654 282880 376660
rect 282840 376009 282868 376654
rect 282826 376000 282882 376009
rect 282826 375935 282882 375944
rect 282828 373992 282880 373998
rect 282826 373960 282828 373969
rect 282880 373960 282882 373969
rect 282826 373895 282882 373904
rect 282828 372564 282880 372570
rect 282828 372506 282880 372512
rect 282840 371929 282868 372506
rect 282826 371920 282882 371929
rect 282826 371855 282882 371864
rect 282368 371068 282420 371074
rect 282368 371010 282420 371016
rect 282380 369889 282408 371010
rect 282366 369880 282422 369889
rect 282366 369815 282422 369824
rect 282276 368076 282328 368082
rect 282276 368018 282328 368024
rect 282288 367849 282316 368018
rect 282274 367840 282330 367849
rect 282274 367775 282330 367784
rect 282828 364336 282880 364342
rect 282828 364278 282880 364284
rect 282840 363769 282868 364278
rect 282826 363760 282882 363769
rect 282826 363695 282882 363704
rect 282826 353560 282882 353569
rect 282932 353546 282960 410518
rect 282882 353518 282960 353546
rect 282826 353495 282882 353504
rect 282826 351520 282882 351529
rect 283024 351506 283052 412082
rect 282882 351478 283052 351506
rect 282826 351455 282882 351464
rect 282826 349480 282882 349489
rect 283116 349466 283144 412150
rect 283196 412072 283248 412078
rect 283196 412014 283248 412020
rect 282882 349438 283144 349466
rect 282826 349415 282882 349424
rect 282826 347712 282882 347721
rect 283208 347698 283236 412014
rect 283288 412004 283340 412010
rect 283288 411946 283340 411952
rect 282882 347670 283236 347698
rect 282826 347647 282882 347656
rect 283300 346118 283328 411946
rect 283380 410644 283432 410650
rect 283380 410586 283432 410592
rect 283288 346112 283340 346118
rect 283288 346054 283340 346060
rect 282828 343596 282880 343602
rect 282828 343538 282880 343544
rect 282840 343369 282868 343538
rect 282826 343360 282882 343369
rect 282826 343295 282882 343304
rect 283392 341358 283420 410586
rect 283484 397118 283512 557466
rect 283472 397112 283524 397118
rect 283472 397054 283524 397060
rect 283380 341352 283432 341358
rect 283380 341294 283432 341300
rect 283576 325106 283604 558146
rect 283668 327078 283696 558175
rect 283748 558136 283800 558142
rect 283748 558078 283800 558084
rect 283760 329118 283788 558078
rect 283840 558068 283892 558074
rect 283840 558010 283892 558016
rect 283852 331158 283880 558010
rect 283944 333266 283972 558826
rect 284208 558816 284260 558822
rect 284208 558758 284260 558764
rect 284116 558748 284168 558754
rect 284116 558690 284168 558696
rect 284024 558544 284076 558550
rect 284024 558486 284076 558492
rect 284036 335238 284064 558486
rect 284128 337618 284156 558690
rect 284220 339318 284248 558758
rect 284956 365838 284984 638930
rect 285312 412480 285364 412486
rect 285312 412422 285364 412428
rect 285220 410848 285272 410854
rect 285220 410790 285272 410796
rect 285128 410780 285180 410786
rect 285128 410722 285180 410728
rect 285036 410712 285088 410718
rect 285036 410654 285088 410660
rect 284944 365832 284996 365838
rect 284944 365774 284996 365780
rect 285048 355910 285076 410654
rect 285140 357678 285168 410722
rect 285232 360194 285260 410790
rect 285324 362914 285352 412422
rect 285404 411936 285456 411942
rect 285404 411878 285456 411884
rect 285416 378078 285444 411878
rect 285404 378072 285456 378078
rect 285404 378014 285456 378020
rect 286336 368082 286364 640290
rect 287716 371074 287744 641718
rect 290476 372570 290504 643078
rect 291856 373998 291884 644438
rect 294604 637628 294656 637634
rect 294604 637570 294656 637576
rect 292578 558648 292634 558657
rect 292578 558583 292580 558592
rect 292632 558583 292634 558592
rect 292580 558554 292632 558560
rect 291844 373992 291896 373998
rect 291844 373934 291896 373940
rect 290464 372564 290516 372570
rect 290464 372506 290516 372512
rect 287704 371068 287756 371074
rect 287704 371010 287756 371016
rect 286324 368076 286376 368082
rect 286324 368018 286376 368024
rect 294616 364342 294644 637570
rect 294708 376718 294736 645866
rect 307114 645008 307170 645017
rect 307114 644943 307170 644952
rect 307128 644502 307156 644943
rect 307116 644496 307168 644502
rect 307116 644438 307168 644444
rect 307114 643512 307170 643521
rect 307114 643447 307170 643456
rect 307128 643142 307156 643447
rect 307116 643136 307168 643142
rect 307116 643078 307168 643084
rect 307666 642152 307722 642161
rect 307666 642087 307722 642096
rect 307680 641782 307708 642087
rect 307668 641776 307720 641782
rect 307668 641718 307720 641724
rect 307666 640520 307722 640529
rect 307666 640455 307722 640464
rect 307680 640354 307708 640455
rect 307668 640348 307720 640354
rect 307668 640290 307720 640296
rect 306654 639432 306710 639441
rect 306654 639367 306710 639376
rect 306668 638994 306696 639367
rect 306656 638988 306708 638994
rect 306656 638930 306708 638936
rect 306838 637936 306894 637945
rect 306838 637871 306894 637880
rect 306852 637634 306880 637871
rect 306840 637628 306892 637634
rect 306840 637570 306892 637576
rect 389178 580952 389234 580961
rect 389178 580887 389234 580896
rect 389192 580310 389220 580887
rect 389180 580304 389232 580310
rect 389180 580246 389232 580252
rect 437848 580304 437900 580310
rect 437848 580246 437900 580252
rect 306930 580000 306986 580009
rect 306930 579935 306986 579944
rect 306944 579698 306972 579935
rect 302884 579692 302936 579698
rect 302884 579634 302936 579640
rect 306932 579692 306984 579698
rect 306932 579634 306984 579640
rect 302146 558648 302202 558657
rect 302146 558583 302202 558592
rect 302160 558550 302188 558583
rect 302148 558544 302200 558550
rect 302148 558486 302200 558492
rect 294696 376712 294748 376718
rect 294696 376654 294748 376660
rect 294604 364336 294656 364342
rect 294604 364278 294656 364284
rect 285312 362908 285364 362914
rect 285312 362850 285364 362856
rect 285220 360188 285272 360194
rect 285220 360130 285272 360136
rect 285128 357672 285180 357678
rect 285128 357614 285180 357620
rect 285036 355904 285088 355910
rect 285036 355846 285088 355852
rect 302896 343602 302924 579634
rect 437860 579193 437888 580246
rect 437846 579184 437902 579193
rect 437846 579119 437902 579128
rect 307668 578944 307720 578950
rect 307666 578912 307668 578921
rect 307720 578912 307722 578921
rect 307666 578847 307722 578856
rect 348422 559328 348478 559337
rect 348422 559263 348478 559272
rect 357714 559328 357770 559337
rect 357714 559263 357770 559272
rect 313738 558920 313794 558929
rect 313738 558855 313794 558864
rect 316038 558920 316094 558929
rect 316038 558855 316094 558864
rect 317418 558920 317474 558929
rect 317418 558855 317420 558864
rect 313752 558278 313780 558855
rect 313740 558272 313792 558278
rect 313740 558214 313792 558220
rect 316052 412486 316080 558855
rect 317472 558855 317474 558864
rect 320270 558920 320326 558929
rect 320270 558855 320326 558864
rect 322846 558920 322902 558929
rect 322846 558855 322902 558864
rect 323490 558920 323546 558929
rect 328550 558920 328606 558929
rect 323490 558855 323546 558864
rect 326344 558884 326396 558890
rect 317420 558826 317472 558832
rect 320284 558822 320312 558855
rect 320272 558816 320324 558822
rect 320178 558784 320234 558793
rect 320272 558758 320324 558764
rect 320178 558719 320180 558728
rect 320232 558719 320234 558728
rect 320180 558690 320232 558696
rect 322860 558686 322888 558855
rect 322848 558680 322900 558686
rect 318798 558648 318854 558657
rect 322848 558622 322900 558628
rect 318798 558583 318854 558592
rect 318812 558550 318840 558583
rect 318800 558544 318852 558550
rect 318800 558486 318852 558492
rect 322860 558278 322888 558622
rect 323504 558618 323532 558855
rect 328550 558855 328606 558864
rect 329562 558920 329618 558929
rect 329562 558855 329618 558864
rect 330482 558920 330538 558929
rect 330482 558855 330538 558864
rect 332506 558920 332562 558929
rect 332506 558855 332562 558864
rect 333150 558920 333206 558929
rect 333150 558855 333206 558864
rect 334254 558920 334310 558929
rect 334254 558855 334256 558864
rect 326344 558826 326396 558832
rect 324964 558748 325016 558754
rect 324964 558690 325016 558696
rect 323492 558612 323544 558618
rect 323492 558554 323544 558560
rect 322848 558272 322900 558278
rect 322848 558214 322900 558220
rect 324976 557705 325004 558690
rect 326356 557705 326384 558826
rect 327724 558680 327776 558686
rect 327724 558622 327776 558628
rect 327736 557705 327764 558622
rect 328564 558414 328592 558855
rect 329576 558482 329604 558855
rect 329564 558476 329616 558482
rect 329564 558418 329616 558424
rect 328552 558408 328604 558414
rect 328552 558350 328604 558356
rect 330496 558346 330524 558855
rect 332520 558822 332548 558855
rect 332508 558816 332560 558822
rect 332508 558758 332560 558764
rect 330484 558340 330536 558346
rect 330484 558282 330536 558288
rect 332520 558278 332548 558758
rect 333164 558618 333192 558855
rect 334308 558855 334310 558864
rect 335910 558920 335966 558929
rect 335910 558855 335966 558864
rect 336278 558920 336334 558929
rect 336278 558855 336334 558864
rect 337750 558920 337806 558929
rect 337750 558855 337806 558864
rect 339038 558920 339094 558929
rect 339038 558855 339094 558864
rect 339866 558920 339922 558929
rect 339866 558855 339922 558864
rect 341246 558920 341302 558929
rect 341246 558855 341302 558864
rect 342534 558920 342590 558929
rect 342534 558855 342590 558864
rect 343638 558920 343694 558929
rect 344834 558920 344890 558929
rect 343638 558855 343640 558864
rect 334256 558826 334308 558832
rect 334268 558754 334296 558826
rect 334256 558748 334308 558754
rect 334256 558690 334308 558696
rect 335924 558686 335952 558855
rect 336292 558754 336320 558855
rect 336280 558748 336332 558754
rect 336280 558690 336332 558696
rect 335912 558680 335964 558686
rect 335912 558622 335964 558628
rect 336292 558618 336320 558690
rect 337764 558618 337792 558855
rect 333152 558612 333204 558618
rect 333152 558554 333204 558560
rect 333888 558612 333940 558618
rect 333888 558554 333940 558560
rect 336280 558612 336332 558618
rect 336280 558554 336332 558560
rect 336740 558612 336792 558618
rect 336740 558554 336792 558560
rect 337752 558612 337804 558618
rect 337752 558554 337804 558560
rect 333900 558346 333928 558554
rect 336752 558414 336780 558554
rect 339052 558482 339080 558855
rect 339040 558476 339092 558482
rect 339040 558418 339092 558424
rect 336740 558408 336792 558414
rect 336740 558350 336792 558356
rect 333888 558340 333940 558346
rect 333888 558282 333940 558288
rect 339880 558278 339908 558855
rect 341260 558822 341288 558855
rect 341248 558816 341300 558822
rect 341248 558758 341300 558764
rect 342548 558346 342576 558855
rect 343692 558855 343694 558864
rect 344744 558884 344796 558890
rect 343640 558826 343692 558832
rect 344834 558855 344836 558864
rect 344744 558826 344796 558832
rect 344888 558855 344890 558864
rect 345754 558920 345810 558929
rect 345754 558855 345810 558864
rect 346490 558920 346546 558929
rect 346490 558855 346546 558864
rect 348238 558920 348294 558929
rect 348238 558855 348294 558864
rect 344836 558826 344888 558832
rect 342536 558340 342588 558346
rect 342536 558282 342588 558288
rect 344756 558278 344784 558826
rect 344848 558686 344876 558826
rect 345768 558754 345796 558855
rect 345756 558748 345808 558754
rect 345756 558690 345808 558696
rect 346504 558686 346532 558855
rect 344836 558680 344888 558686
rect 344836 558622 344888 558628
rect 346492 558680 346544 558686
rect 346492 558622 346544 558628
rect 346504 558482 346532 558622
rect 348252 558482 348280 558855
rect 346492 558476 346544 558482
rect 346492 558418 346544 558424
rect 348240 558476 348292 558482
rect 348240 558418 348292 558424
rect 348436 558414 348464 559263
rect 349342 558920 349398 558929
rect 349342 558855 349398 558864
rect 350538 558920 350594 558929
rect 350538 558855 350594 558864
rect 352010 558920 352066 558929
rect 352010 558855 352066 558864
rect 353298 558920 353354 558929
rect 353298 558855 353300 558864
rect 349356 558754 349384 558855
rect 350552 558822 350580 558855
rect 350540 558816 350592 558822
rect 350540 558758 350592 558764
rect 349344 558748 349396 558754
rect 349344 558690 349396 558696
rect 348424 558408 348476 558414
rect 348424 558350 348476 558356
rect 349356 558346 349384 558690
rect 349344 558340 349396 558346
rect 349344 558282 349396 558288
rect 352024 558278 352052 558855
rect 353352 558855 353354 558864
rect 353300 558826 353352 558832
rect 354678 558784 354734 558793
rect 354678 558719 354734 558728
rect 356058 558784 356114 558793
rect 356058 558719 356114 558728
rect 354692 558618 354720 558719
rect 356072 558686 356100 558719
rect 356060 558680 356112 558686
rect 356060 558622 356112 558628
rect 354680 558612 354732 558618
rect 354680 558554 354732 558560
rect 357438 558512 357494 558521
rect 357438 558447 357440 558456
rect 357492 558447 357494 558456
rect 357440 558418 357492 558424
rect 356702 558376 356758 558385
rect 357728 558346 357756 559263
rect 418252 558680 418304 558686
rect 418252 558622 418304 558628
rect 383568 558544 383620 558550
rect 383568 558486 383620 558492
rect 358084 558476 358136 558482
rect 358084 558418 358136 558424
rect 356702 558311 356758 558320
rect 357716 558340 357768 558346
rect 332508 558272 332560 558278
rect 332508 558214 332560 558220
rect 339868 558272 339920 558278
rect 339868 558214 339920 558220
rect 344744 558272 344796 558278
rect 344744 558214 344796 558220
rect 352012 558272 352064 558278
rect 352012 558214 352064 558220
rect 324962 557696 325018 557705
rect 324962 557631 325018 557640
rect 326342 557696 326398 557705
rect 326342 557631 326398 557640
rect 327722 557696 327778 557705
rect 327722 557631 327778 557640
rect 329930 557696 329986 557705
rect 329930 557631 329986 557640
rect 336830 557696 336886 557705
rect 336830 557631 336886 557640
rect 343730 557696 343786 557705
rect 343730 557631 343786 557640
rect 352010 557696 352066 557705
rect 352010 557631 352066 557640
rect 321558 557560 321614 557569
rect 321558 557495 321614 557504
rect 322938 557560 322994 557569
rect 322938 557495 322994 557504
rect 324318 557560 324374 557569
rect 324318 557495 324374 557504
rect 316040 412480 316092 412486
rect 316040 412422 316092 412428
rect 321572 411262 321600 557495
rect 322952 413982 322980 557495
rect 324332 415410 324360 557495
rect 324320 415404 324372 415410
rect 324320 415346 324372 415352
rect 322940 413976 322992 413982
rect 322940 413918 322992 413924
rect 324976 412418 325004 557631
rect 325698 557560 325754 557569
rect 325698 557495 325754 557504
rect 325712 418130 325740 557495
rect 325700 418124 325752 418130
rect 325700 418066 325752 418072
rect 324964 412412 325016 412418
rect 324964 412354 325016 412360
rect 326356 412350 326384 557631
rect 327078 557560 327134 557569
rect 327078 557495 327134 557504
rect 327092 419490 327120 557495
rect 327080 419484 327132 419490
rect 327080 419426 327132 419432
rect 326344 412344 326396 412350
rect 326344 412286 326396 412292
rect 327736 412282 327764 557631
rect 328458 557560 328514 557569
rect 328458 557495 328514 557504
rect 329838 557560 329894 557569
rect 329838 557495 329894 557504
rect 328472 420918 328500 557495
rect 329852 423638 329880 557495
rect 329944 425066 329972 557631
rect 331218 557560 331274 557569
rect 331218 557495 331274 557504
rect 332598 557560 332654 557569
rect 332598 557495 332654 557504
rect 333978 557560 334034 557569
rect 333978 557495 334034 557504
rect 335358 557560 335414 557569
rect 335358 557495 335414 557504
rect 336738 557560 336794 557569
rect 336738 557495 336794 557504
rect 331232 427786 331260 557495
rect 332612 429146 332640 557495
rect 333992 431934 334020 557495
rect 335372 433294 335400 557495
rect 336752 436082 336780 557495
rect 336844 437442 336872 557631
rect 338118 557560 338174 557569
rect 338118 557495 338174 557504
rect 339498 557560 339554 557569
rect 339498 557495 339554 557504
rect 340878 557560 340934 557569
rect 340878 557495 340934 557504
rect 342258 557560 342314 557569
rect 342258 557495 342314 557504
rect 343638 557560 343694 557569
rect 343638 557495 343694 557504
rect 338132 440230 338160 557495
rect 339512 441590 339540 557495
rect 340892 444378 340920 557495
rect 342272 445738 342300 557495
rect 343652 448526 343680 557495
rect 343744 449886 343772 557631
rect 345018 557560 345074 557569
rect 345018 557495 345074 557504
rect 346398 557560 346454 557569
rect 346398 557495 346454 557504
rect 347778 557560 347834 557569
rect 347778 557495 347834 557504
rect 349158 557560 349214 557569
rect 349158 557495 349214 557504
rect 350538 557560 350594 557569
rect 350538 557495 350594 557504
rect 345032 452606 345060 557495
rect 346412 454034 346440 557495
rect 347792 455394 347820 557495
rect 349172 458182 349200 557495
rect 350552 459542 350580 557495
rect 352024 463690 352052 557631
rect 353298 557560 353354 557569
rect 353298 557495 353354 557504
rect 354678 557560 354734 557569
rect 354678 557495 354734 557504
rect 356058 557560 356114 557569
rect 356058 557495 356114 557504
rect 352194 555520 352250 555529
rect 352194 555455 352250 555464
rect 352012 463684 352064 463690
rect 352012 463626 352064 463632
rect 352208 462330 352236 555455
rect 353312 466410 353340 557495
rect 354692 467838 354720 557495
rect 356072 470558 356100 557495
rect 356716 514758 356744 558311
rect 357716 558282 357768 558288
rect 357530 557560 357586 557569
rect 357530 557495 357586 557504
rect 356704 514752 356756 514758
rect 356704 514694 356756 514700
rect 357544 471986 357572 557495
rect 358096 478854 358124 558418
rect 359464 558408 359516 558414
rect 359464 558350 359516 558356
rect 358176 558272 358228 558278
rect 358176 558214 358228 558220
rect 358188 517478 358216 558214
rect 358910 555520 358966 555529
rect 358910 555455 358966 555464
rect 358176 517472 358228 517478
rect 358176 517414 358228 517420
rect 358084 478848 358136 478854
rect 358084 478790 358136 478796
rect 358924 474706 358952 555455
rect 359476 518906 359504 558350
rect 359556 558340 359608 558346
rect 359556 558282 359608 558288
rect 359568 521626 359596 558282
rect 359556 521620 359608 521626
rect 359556 521562 359608 521568
rect 359464 518900 359516 518906
rect 359464 518842 359516 518848
rect 358912 474700 358964 474706
rect 358912 474642 358964 474648
rect 357532 471980 357584 471986
rect 357532 471922 357584 471928
rect 356060 470552 356112 470558
rect 356060 470494 356112 470500
rect 354680 467832 354732 467838
rect 354680 467774 354732 467780
rect 353300 466404 353352 466410
rect 353300 466346 353352 466352
rect 352196 462324 352248 462330
rect 352196 462266 352248 462272
rect 350540 459536 350592 459542
rect 350540 459478 350592 459484
rect 349160 458176 349212 458182
rect 349160 458118 349212 458124
rect 347780 455388 347832 455394
rect 347780 455330 347832 455336
rect 346400 454028 346452 454034
rect 346400 453970 346452 453976
rect 345020 452600 345072 452606
rect 345020 452542 345072 452548
rect 343732 449880 343784 449886
rect 343732 449822 343784 449828
rect 343640 448520 343692 448526
rect 343640 448462 343692 448468
rect 342260 445732 342312 445738
rect 342260 445674 342312 445680
rect 340880 444372 340932 444378
rect 340880 444314 340932 444320
rect 339500 441584 339552 441590
rect 339500 441526 339552 441532
rect 338120 440224 338172 440230
rect 338120 440166 338172 440172
rect 336832 437436 336884 437442
rect 336832 437378 336884 437384
rect 336740 436076 336792 436082
rect 336740 436018 336792 436024
rect 335360 433288 335412 433294
rect 335360 433230 335412 433236
rect 333980 431928 334032 431934
rect 333980 431870 334032 431876
rect 332600 429140 332652 429146
rect 332600 429082 332652 429088
rect 331220 427780 331272 427786
rect 331220 427722 331272 427728
rect 329932 425060 329984 425066
rect 329932 425002 329984 425008
rect 329840 423632 329892 423638
rect 329840 423574 329892 423580
rect 328460 420912 328512 420918
rect 328460 420854 328512 420860
rect 383580 413302 383608 558486
rect 418264 558142 418292 558622
rect 418252 558136 418304 558142
rect 418252 558078 418304 558084
rect 418160 558068 418212 558074
rect 418160 558010 418212 558016
rect 432604 558068 432656 558074
rect 432604 558010 432656 558016
rect 418172 557954 418200 558010
rect 418172 557926 418384 557954
rect 418356 557598 418384 557926
rect 432616 557682 432644 558010
rect 432524 557654 432644 557682
rect 432524 557598 432552 557654
rect 418344 557592 418396 557598
rect 418344 557534 418396 557540
rect 432512 557592 432564 557598
rect 432512 557534 432564 557540
rect 383568 413296 383620 413302
rect 383566 413264 383568 413273
rect 405004 413296 405056 413302
rect 383620 413264 383622 413273
rect 405004 413238 405056 413244
rect 383566 413199 383622 413208
rect 405016 412690 405044 413238
rect 405004 412684 405056 412690
rect 405004 412626 405056 412632
rect 327724 412276 327776 412282
rect 327724 412218 327776 412224
rect 321560 411256 321612 411262
rect 321560 411198 321612 411204
rect 302884 343596 302936 343602
rect 302884 343538 302936 343544
rect 284208 339312 284260 339318
rect 284208 339254 284260 339260
rect 284116 337612 284168 337618
rect 284116 337554 284168 337560
rect 284024 335232 284076 335238
rect 284024 335174 284076 335180
rect 283932 333260 283984 333266
rect 283932 333202 283984 333208
rect 283840 331152 283892 331158
rect 283840 331094 283892 331100
rect 283748 329112 283800 329118
rect 283748 329054 283800 329060
rect 283656 327072 283708 327078
rect 283656 327014 283708 327020
rect 283564 325100 283616 325106
rect 283564 325042 283616 325048
rect 282182 321056 282238 321065
rect 282182 320991 282238 321000
rect 62500 320198 62882 320226
rect 79060 320198 79442 320226
rect 88996 320198 89378 320226
rect 100142 320198 100524 320226
rect 101430 320198 101812 320226
rect 104190 320198 104572 320226
rect 210542 320198 210924 320226
rect 214590 320198 214972 320226
rect 233910 320198 234292 320226
rect 250470 320198 250852 320226
rect 60016 320062 60214 320090
rect 60292 320062 60582 320090
rect 60844 320062 61042 320090
rect 61120 320062 61502 320090
rect 59360 318980 59412 318986
rect 59360 318922 59412 318928
rect 30288 318776 30340 318782
rect 30288 318718 30340 318724
rect 30196 318640 30248 318646
rect 30196 318582 30248 318588
rect 23388 318572 23440 318578
rect 23388 318514 23440 318520
rect 12346 318472 12402 318481
rect 12346 318407 12402 318416
rect 22008 318436 22060 318442
rect 9586 318200 9642 318209
rect 9586 318135 9642 318144
rect 5446 318064 5502 318073
rect 5446 317999 5502 318008
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 4066 3496 4122 3505
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 4066 3431 4122 3440
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 2884 480 2912 3295
rect 4080 480 4108 3431
rect 5460 610 5488 317999
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5448 604 5500 610
rect 5448 546 5500 552
rect 5276 480 5304 546
rect 6472 480 6500 3538
rect 7668 480 7696 3606
rect 9600 3126 9628 318135
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 8864 480 8892 3062
rect 10060 480 10088 3674
rect 12360 3398 12388 318407
rect 22008 318378 22060 318384
rect 20628 318368 20680 318374
rect 13634 318336 13690 318345
rect 20628 318310 20680 318316
rect 13634 318271 13690 318280
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 11256 480 11284 3334
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12452 480 12480 3130
rect 13648 480 13676 318271
rect 17868 318164 17920 318170
rect 17868 318106 17920 318112
rect 13728 318096 13780 318102
rect 13728 318038 13780 318044
rect 13740 3194 13768 318038
rect 16028 3868 16080 3874
rect 16028 3810 16080 3816
rect 14832 3800 14884 3806
rect 14832 3742 14884 3748
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 14844 480 14872 3742
rect 16040 480 16068 3810
rect 17880 3398 17908 318106
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17236 480 17264 3334
rect 18340 480 18368 3878
rect 20640 3398 20668 318310
rect 21916 318300 21968 318306
rect 21916 318242 21968 318248
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 19536 480 19564 3334
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20732 480 20760 2926
rect 21928 480 21956 318242
rect 22020 2990 22048 318378
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 23400 610 23428 318514
rect 27528 318504 27580 318510
rect 27528 318446 27580 318452
rect 25504 4004 25556 4010
rect 25504 3946 25556 3952
rect 24306 3632 24362 3641
rect 24306 3567 24362 3576
rect 23112 604 23164 610
rect 23112 546 23164 552
rect 23388 604 23440 610
rect 23388 546 23440 552
rect 23124 480 23152 546
rect 24320 480 24348 3567
rect 25516 480 25544 3946
rect 27540 3398 27568 318446
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 26712 480 26740 3334
rect 27908 480 27936 3334
rect 29104 480 29132 4014
rect 30208 3482 30236 318582
rect 30300 4078 30328 318718
rect 31668 318708 31720 318714
rect 31668 318650 31720 318656
rect 30288 4072 30340 4078
rect 30288 4014 30340 4020
rect 31680 3482 31708 318650
rect 38476 318028 38528 318034
rect 38476 317970 38528 317976
rect 37188 317960 37240 317966
rect 37188 317902 37240 317908
rect 34978 3768 35034 3777
rect 34978 3703 35034 3712
rect 30208 3454 30328 3482
rect 30300 480 30328 3454
rect 31496 3454 31708 3482
rect 31496 480 31524 3454
rect 33876 3392 33928 3398
rect 33876 3334 33928 3340
rect 32680 3324 32732 3330
rect 32680 3266 32732 3272
rect 32692 480 32720 3266
rect 33888 480 33916 3334
rect 34992 480 35020 3703
rect 37200 3330 37228 317902
rect 37372 4140 37424 4146
rect 37372 4082 37424 4088
rect 36176 3324 36228 3330
rect 36176 3266 36228 3272
rect 37188 3324 37240 3330
rect 37188 3266 37240 3272
rect 36188 480 36216 3266
rect 37384 480 37412 4082
rect 38488 3482 38516 317970
rect 44088 317892 44140 317898
rect 44088 317834 44140 317840
rect 38568 317824 38620 317830
rect 38568 317766 38620 317772
rect 38580 4146 38608 317766
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 40958 4040 41014 4049
rect 40958 3975 41014 3984
rect 39762 3904 39818 3913
rect 39762 3839 39818 3848
rect 38488 3454 38608 3482
rect 38580 480 38608 3454
rect 39776 480 39804 3839
rect 40972 480 41000 3975
rect 44100 3330 44128 317834
rect 45468 317756 45520 317762
rect 45468 317698 45520 317704
rect 45480 3330 45508 317698
rect 50988 317688 51040 317694
rect 50988 317630 51040 317636
rect 46848 317620 46900 317626
rect 46848 317562 46900 317568
rect 46860 3330 46888 317562
rect 51000 3330 51028 317630
rect 53748 317552 53800 317558
rect 53748 317494 53800 317500
rect 53760 3330 53788 317494
rect 57888 317484 57940 317490
rect 57888 317426 57940 317432
rect 55220 4820 55272 4826
rect 55220 4762 55272 4768
rect 43352 3324 43404 3330
rect 43352 3266 43404 3272
rect 44088 3324 44140 3330
rect 44088 3266 44140 3272
rect 44548 3324 44600 3330
rect 44548 3266 44600 3272
rect 45468 3324 45520 3330
rect 45468 3266 45520 3272
rect 45744 3324 45796 3330
rect 45744 3266 45796 3272
rect 46848 3324 46900 3330
rect 46848 3266 46900 3272
rect 50528 3324 50580 3330
rect 50528 3266 50580 3272
rect 50988 3324 51040 3330
rect 50988 3266 51040 3272
rect 52828 3324 52880 3330
rect 52828 3266 52880 3272
rect 53748 3324 53800 3330
rect 53748 3266 53800 3272
rect 42156 3256 42208 3262
rect 42156 3198 42208 3204
rect 42168 480 42196 3198
rect 43364 480 43392 3266
rect 44560 480 44588 3266
rect 45756 480 45784 3266
rect 48136 3188 48188 3194
rect 48136 3130 48188 3136
rect 46940 2916 46992 2922
rect 46940 2858 46992 2864
rect 46952 480 46980 2858
rect 48148 480 48176 3130
rect 49332 3120 49384 3126
rect 49332 3062 49384 3068
rect 49344 480 49372 3062
rect 50540 480 50568 3266
rect 51632 3052 51684 3058
rect 51632 2994 51684 3000
rect 51644 480 51672 2994
rect 52840 480 52868 3266
rect 54024 2984 54076 2990
rect 54024 2926 54076 2932
rect 54036 480 54064 2926
rect 55232 480 55260 4762
rect 56416 2916 56468 2922
rect 56416 2858 56468 2864
rect 56428 480 56456 2858
rect 57900 626 57928 317426
rect 59372 3534 59400 318922
rect 60016 317914 60044 320062
rect 60292 318986 60320 320062
rect 60280 318980 60332 318986
rect 60280 318922 60332 318928
rect 60740 318300 60792 318306
rect 60740 318242 60792 318248
rect 60752 318102 60780 318242
rect 60372 318096 60424 318102
rect 60372 318038 60424 318044
rect 60740 318096 60792 318102
rect 60740 318038 60792 318044
rect 60384 317914 60412 318038
rect 60016 317886 60412 317914
rect 60016 3618 60044 317886
rect 60740 315988 60792 315994
rect 60740 315930 60792 315936
rect 59924 3590 60044 3618
rect 59360 3528 59412 3534
rect 59360 3470 59412 3476
rect 59924 3466 59952 3590
rect 60004 3528 60056 3534
rect 60752 3505 60780 315930
rect 60004 3470 60056 3476
rect 60738 3496 60794 3505
rect 59912 3460 59964 3466
rect 59912 3402 59964 3408
rect 58808 2848 58860 2854
rect 58808 2790 58860 2796
rect 57624 598 57928 626
rect 57624 480 57652 598
rect 58820 480 58848 2790
rect 60016 480 60044 3470
rect 60738 3431 60794 3440
rect 60844 3369 60872 320062
rect 61120 315994 61148 320062
rect 61948 318073 61976 320076
rect 62132 320062 62422 320090
rect 61934 318064 61990 318073
rect 61934 317999 61990 318008
rect 61108 315988 61160 315994
rect 61108 315930 61160 315936
rect 62132 3602 62160 320062
rect 62500 316010 62528 320198
rect 63328 318209 63356 320076
rect 63604 320062 63802 320090
rect 63314 318200 63370 318209
rect 63314 318135 63370 318144
rect 62224 315982 62528 316010
rect 62224 3670 62252 315982
rect 63604 3738 63632 320062
rect 64156 318481 64184 320076
rect 64616 318578 64644 320076
rect 64604 318572 64656 318578
rect 64604 318514 64656 318520
rect 64142 318472 64198 318481
rect 64142 318407 64198 318416
rect 65076 318345 65104 320076
rect 65260 320062 65550 320090
rect 65720 320062 66010 320090
rect 65062 318336 65118 318345
rect 65062 318271 65118 318280
rect 65260 316010 65288 320062
rect 64880 315988 64932 315994
rect 64880 315930 64932 315936
rect 64984 315982 65288 316010
rect 65720 315994 65748 320062
rect 66456 318170 66484 320076
rect 66824 320062 66930 320090
rect 66444 318164 66496 318170
rect 66444 318106 66496 318112
rect 65708 315988 65760 315994
rect 64892 3874 64920 315930
rect 64880 3868 64932 3874
rect 64880 3810 64932 3816
rect 64984 3806 65012 315982
rect 65708 315930 65760 315936
rect 66824 313954 66852 320062
rect 67376 318374 67404 320076
rect 67744 318442 67772 320076
rect 67732 318436 67784 318442
rect 67732 318378 67784 318384
rect 67364 318368 67416 318374
rect 67364 318310 67416 318316
rect 68204 318102 68232 320076
rect 68664 318510 68692 320076
rect 69138 320062 69336 320090
rect 68652 318504 68704 318510
rect 68652 318446 68704 318452
rect 68192 318096 68244 318102
rect 68192 318038 68244 318044
rect 69112 315988 69164 315994
rect 69112 315930 69164 315936
rect 66812 313948 66864 313954
rect 66812 313890 66864 313896
rect 66996 313948 67048 313954
rect 66996 313890 67048 313896
rect 67008 309126 67036 313890
rect 66996 309120 67048 309126
rect 66996 309062 67048 309068
rect 66812 299532 66864 299538
rect 66812 299474 66864 299480
rect 66824 294642 66852 299474
rect 66628 294636 66680 294642
rect 66628 294578 66680 294584
rect 66812 294636 66864 294642
rect 66812 294578 66864 294584
rect 66640 282826 66668 294578
rect 66548 282798 66668 282826
rect 66548 280158 66576 282798
rect 66536 280152 66588 280158
rect 66536 280094 66588 280100
rect 66628 270564 66680 270570
rect 66628 270506 66680 270512
rect 66640 263514 66668 270506
rect 66548 263486 66668 263514
rect 66548 260846 66576 263486
rect 66536 260840 66588 260846
rect 66536 260782 66588 260788
rect 66628 251252 66680 251258
rect 66628 251194 66680 251200
rect 66640 244202 66668 251194
rect 66548 244174 66668 244202
rect 66548 241505 66576 244174
rect 66350 241496 66406 241505
rect 66350 241431 66406 241440
rect 66534 241496 66590 241505
rect 66534 241431 66590 241440
rect 66364 231878 66392 241431
rect 66352 231872 66404 231878
rect 66352 231814 66404 231820
rect 66628 231872 66680 231878
rect 66628 231814 66680 231820
rect 66640 224890 66668 231814
rect 66548 224862 66668 224890
rect 66548 222193 66576 224862
rect 66350 222184 66406 222193
rect 66350 222119 66406 222128
rect 66534 222184 66590 222193
rect 66534 222119 66590 222128
rect 66364 212566 66392 222119
rect 66352 212560 66404 212566
rect 66352 212502 66404 212508
rect 66628 212560 66680 212566
rect 66628 212502 66680 212508
rect 66640 205578 66668 212502
rect 66548 205550 66668 205578
rect 66548 202881 66576 205550
rect 66350 202872 66406 202881
rect 66350 202807 66406 202816
rect 66534 202872 66590 202881
rect 66534 202807 66590 202816
rect 66364 193254 66392 202807
rect 66352 193248 66404 193254
rect 66352 193190 66404 193196
rect 66628 193248 66680 193254
rect 66628 193190 66680 193196
rect 66640 186266 66668 193190
rect 66548 186238 66668 186266
rect 66548 183569 66576 186238
rect 66350 183560 66406 183569
rect 66350 183495 66406 183504
rect 66534 183560 66590 183569
rect 66534 183495 66590 183504
rect 66364 173942 66392 183495
rect 66352 173936 66404 173942
rect 66352 173878 66404 173884
rect 66628 173936 66680 173942
rect 66628 173878 66680 173884
rect 66640 166954 66668 173878
rect 66548 166926 66668 166954
rect 66548 164218 66576 166926
rect 66352 164212 66404 164218
rect 66352 164154 66404 164160
rect 66536 164212 66588 164218
rect 66536 164154 66588 164160
rect 66364 154601 66392 164154
rect 66350 154592 66406 154601
rect 66350 154527 66406 154536
rect 66626 154592 66682 154601
rect 66626 154527 66682 154536
rect 66640 147642 66668 154527
rect 66548 147614 66668 147642
rect 66548 140026 66576 147614
rect 66364 139998 66576 140026
rect 66364 135289 66392 139998
rect 66350 135280 66406 135289
rect 66350 135215 66406 135224
rect 66626 135280 66682 135289
rect 66626 135215 66682 135224
rect 66640 128330 66668 135215
rect 66548 128302 66668 128330
rect 66548 120714 66576 128302
rect 66364 120686 66576 120714
rect 66364 115977 66392 120686
rect 66350 115968 66406 115977
rect 66350 115903 66406 115912
rect 66626 115968 66682 115977
rect 66626 115903 66682 115912
rect 66640 109018 66668 115903
rect 66548 108990 66668 109018
rect 66548 101402 66576 108990
rect 66364 101374 66576 101402
rect 66364 96665 66392 101374
rect 66350 96656 66406 96665
rect 66350 96591 66406 96600
rect 66626 96656 66682 96665
rect 66626 96591 66682 96600
rect 66640 89706 66668 96591
rect 66456 89678 66668 89706
rect 66456 86970 66484 89678
rect 66444 86964 66496 86970
rect 66444 86906 66496 86912
rect 66352 77308 66404 77314
rect 66352 77250 66404 77256
rect 66364 77178 66392 77250
rect 66352 77172 66404 77178
rect 66352 77114 66404 77120
rect 66444 70304 66496 70310
rect 66444 70246 66496 70252
rect 66456 60722 66484 70246
rect 66444 60716 66496 60722
rect 66444 60658 66496 60664
rect 66628 60716 66680 60722
rect 66628 60658 66680 60664
rect 66640 57934 66668 60658
rect 66628 57928 66680 57934
rect 66628 57870 66680 57876
rect 66536 48340 66588 48346
rect 66536 48282 66588 48288
rect 66548 41426 66576 48282
rect 66456 41410 66576 41426
rect 66444 41404 66576 41410
rect 66496 41398 66576 41404
rect 66628 41404 66680 41410
rect 66444 41346 66496 41352
rect 66628 41346 66680 41352
rect 66640 38622 66668 41346
rect 66628 38616 66680 38622
rect 66628 38558 66680 38564
rect 66536 29028 66588 29034
rect 66536 28970 66588 28976
rect 66548 22114 66576 28970
rect 66456 22098 66576 22114
rect 66444 22092 66576 22098
rect 66496 22086 66576 22092
rect 66628 22092 66680 22098
rect 66444 22034 66496 22040
rect 66628 22034 66680 22040
rect 66640 19310 66668 22034
rect 66628 19304 66680 19310
rect 66628 19246 66680 19252
rect 66628 9716 66680 9722
rect 66628 9658 66680 9664
rect 66640 3942 66668 9658
rect 69124 4010 69152 315930
rect 69112 4004 69164 4010
rect 69112 3946 69164 3952
rect 66628 3936 66680 3942
rect 66628 3878 66680 3884
rect 67180 3936 67232 3942
rect 67180 3878 67232 3884
rect 64972 3800 65024 3806
rect 64972 3742 65024 3748
rect 63592 3732 63644 3738
rect 63592 3674 63644 3680
rect 62212 3664 62264 3670
rect 62212 3606 62264 3612
rect 62396 3664 62448 3670
rect 62396 3606 62448 3612
rect 65984 3664 66036 3670
rect 65984 3606 66036 3612
rect 62120 3596 62172 3602
rect 62120 3538 62172 3544
rect 61200 3460 61252 3466
rect 61200 3402 61252 3408
rect 60830 3360 60886 3369
rect 60830 3295 60886 3304
rect 61212 480 61240 3402
rect 62408 480 62436 3606
rect 63592 3596 63644 3602
rect 63592 3538 63644 3544
rect 64788 3596 64840 3602
rect 64788 3538 64840 3544
rect 63604 480 63632 3538
rect 64800 480 64828 3538
rect 65996 480 66024 3606
rect 67192 480 67220 3878
rect 68284 3800 68336 3806
rect 68284 3742 68336 3748
rect 68296 480 68324 3742
rect 69308 3641 69336 320062
rect 69400 320062 69598 320090
rect 69400 315994 69428 320062
rect 70044 318306 70072 320076
rect 70518 320062 70624 320090
rect 70032 318300 70084 318306
rect 70032 318242 70084 318248
rect 69388 315988 69440 315994
rect 69388 315930 69440 315936
rect 70596 4282 70624 320062
rect 70964 318782 70992 320076
rect 70952 318776 71004 318782
rect 70952 318718 71004 318724
rect 71332 318646 71360 320076
rect 71792 318714 71820 320076
rect 71884 320062 72266 320090
rect 72344 320062 72726 320090
rect 73186 320062 73292 320090
rect 71780 318708 71832 318714
rect 71780 318650 71832 318656
rect 71320 318640 71372 318646
rect 71320 318582 71372 318588
rect 71884 5234 71912 320062
rect 72344 292670 72372 320062
rect 72332 292664 72384 292670
rect 72332 292606 72384 292612
rect 72240 289876 72292 289882
rect 72240 289818 72292 289824
rect 72252 280158 72280 289818
rect 72240 280152 72292 280158
rect 72240 280094 72292 280100
rect 72240 270564 72292 270570
rect 72240 270506 72292 270512
rect 72252 260846 72280 270506
rect 72240 260840 72292 260846
rect 72240 260782 72292 260788
rect 72240 251252 72292 251258
rect 72240 251194 72292 251200
rect 72252 241505 72280 251194
rect 72054 241496 72110 241505
rect 72054 241431 72110 241440
rect 72238 241496 72294 241505
rect 72238 241431 72294 241440
rect 72068 231878 72096 241431
rect 72056 231872 72108 231878
rect 72056 231814 72108 231820
rect 72240 231872 72292 231878
rect 72240 231814 72292 231820
rect 72252 222193 72280 231814
rect 72054 222184 72110 222193
rect 72054 222119 72110 222128
rect 72238 222184 72294 222193
rect 72238 222119 72294 222128
rect 72068 212566 72096 222119
rect 72056 212560 72108 212566
rect 72056 212502 72108 212508
rect 72240 212560 72292 212566
rect 72240 212502 72292 212508
rect 72252 202881 72280 212502
rect 72054 202872 72110 202881
rect 72054 202807 72110 202816
rect 72238 202872 72294 202881
rect 72238 202807 72294 202816
rect 72068 193254 72096 202807
rect 72056 193248 72108 193254
rect 72056 193190 72108 193196
rect 72240 193248 72292 193254
rect 72240 193190 72292 193196
rect 72252 183569 72280 193190
rect 72054 183560 72110 183569
rect 72054 183495 72110 183504
rect 72238 183560 72294 183569
rect 72238 183495 72294 183504
rect 72068 173942 72096 183495
rect 72056 173936 72108 173942
rect 72056 173878 72108 173884
rect 72240 173936 72292 173942
rect 72240 173878 72292 173884
rect 72252 157434 72280 173878
rect 72160 157406 72280 157434
rect 72160 157298 72188 157406
rect 72160 157270 72280 157298
rect 72252 145081 72280 157270
rect 72238 145072 72294 145081
rect 72238 145007 72294 145016
rect 72238 144936 72294 144945
rect 72238 144871 72294 144880
rect 72252 125769 72280 144871
rect 72238 125760 72294 125769
rect 72238 125695 72294 125704
rect 72238 125624 72294 125633
rect 72238 125559 72294 125568
rect 72252 122806 72280 125559
rect 72240 122800 72292 122806
rect 72240 122742 72292 122748
rect 72240 113212 72292 113218
rect 72240 113154 72292 113160
rect 72252 104836 72280 113154
rect 72252 104808 72372 104836
rect 72344 102134 72372 104808
rect 72332 102128 72384 102134
rect 72332 102070 72384 102076
rect 72240 92540 72292 92546
rect 72240 92482 72292 92488
rect 72252 71074 72280 92482
rect 72160 71046 72280 71074
rect 72160 66230 72188 71046
rect 72148 66224 72200 66230
rect 72148 66166 72200 66172
rect 72424 66224 72476 66230
rect 72424 66166 72476 66172
rect 72436 64870 72464 66166
rect 72424 64864 72476 64870
rect 72424 64806 72476 64812
rect 72424 56568 72476 56574
rect 72424 56510 72476 56516
rect 72436 55214 72464 56510
rect 72424 55208 72476 55214
rect 72424 55150 72476 55156
rect 72332 45688 72384 45694
rect 72332 45630 72384 45636
rect 72344 45558 72372 45630
rect 72332 45552 72384 45558
rect 72332 45494 72384 45500
rect 72148 31748 72200 31754
rect 72148 31690 72200 31696
rect 72160 27606 72188 31690
rect 72148 27600 72200 27606
rect 72148 27542 72200 27548
rect 72332 27532 72384 27538
rect 72332 27474 72384 27480
rect 72344 9722 72372 27474
rect 72056 9716 72108 9722
rect 72056 9658 72108 9664
rect 72332 9716 72384 9722
rect 72332 9658 72384 9664
rect 71872 5228 71924 5234
rect 71872 5170 71924 5176
rect 70584 4276 70636 4282
rect 70584 4218 70636 4224
rect 72068 4010 72096 9658
rect 72148 4140 72200 4146
rect 72148 4082 72200 4088
rect 72056 4004 72108 4010
rect 72056 3946 72108 3952
rect 69294 3632 69350 3641
rect 69294 3567 69350 3576
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 69480 3324 69532 3330
rect 69480 3266 69532 3272
rect 69492 480 69520 3266
rect 70688 480 70716 3334
rect 72160 1986 72188 4082
rect 73068 4004 73120 4010
rect 73068 3946 73120 3952
rect 71884 1958 72188 1986
rect 71884 480 71912 1958
rect 73080 480 73108 3946
rect 73264 3777 73292 320062
rect 73632 317966 73660 320076
rect 73620 317960 73672 317966
rect 73620 317902 73672 317908
rect 74092 317830 74120 320076
rect 74448 318096 74500 318102
rect 74448 318038 74500 318044
rect 74080 317824 74132 317830
rect 74080 317766 74132 317772
rect 74460 309126 74488 318038
rect 74552 318034 74580 320076
rect 74644 320062 75026 320090
rect 75104 320062 75394 320090
rect 75472 320062 75854 320090
rect 74540 318028 74592 318034
rect 74540 317970 74592 317976
rect 74448 309120 74500 309126
rect 74448 309062 74500 309068
rect 74448 299532 74500 299538
rect 74448 299474 74500 299480
rect 74460 298110 74488 299474
rect 74448 298104 74500 298110
rect 74448 298046 74500 298052
rect 74448 280220 74500 280226
rect 74448 280162 74500 280168
rect 74460 278769 74488 280162
rect 74262 278760 74318 278769
rect 74262 278695 74318 278704
rect 74446 278760 74502 278769
rect 74446 278695 74502 278704
rect 74276 269142 74304 278695
rect 74264 269136 74316 269142
rect 74264 269078 74316 269084
rect 74448 269136 74500 269142
rect 74448 269078 74500 269084
rect 74460 259457 74488 269078
rect 74262 259448 74318 259457
rect 74262 259383 74318 259392
rect 74446 259448 74502 259457
rect 74446 259383 74502 259392
rect 74276 249830 74304 259383
rect 74264 249824 74316 249830
rect 74264 249766 74316 249772
rect 74448 249824 74500 249830
rect 74448 249766 74500 249772
rect 74460 240145 74488 249766
rect 74262 240136 74318 240145
rect 74262 240071 74318 240080
rect 74446 240136 74502 240145
rect 74446 240071 74502 240080
rect 74276 230518 74304 240071
rect 74264 230512 74316 230518
rect 74264 230454 74316 230460
rect 74448 230512 74500 230518
rect 74448 230454 74500 230460
rect 74460 220833 74488 230454
rect 74262 220824 74318 220833
rect 74262 220759 74318 220768
rect 74446 220824 74502 220833
rect 74446 220759 74502 220768
rect 74276 211177 74304 220759
rect 74262 211168 74318 211177
rect 74262 211103 74318 211112
rect 74446 211168 74502 211177
rect 74446 211103 74502 211112
rect 74460 201482 74488 211103
rect 74264 201476 74316 201482
rect 74264 201418 74316 201424
rect 74448 201476 74500 201482
rect 74448 201418 74500 201424
rect 74276 191865 74304 201418
rect 74262 191856 74318 191865
rect 74262 191791 74318 191800
rect 74446 191856 74502 191865
rect 74446 191791 74502 191800
rect 74460 182170 74488 191791
rect 74264 182164 74316 182170
rect 74264 182106 74316 182112
rect 74448 182164 74500 182170
rect 74448 182106 74500 182112
rect 74276 172553 74304 182106
rect 74262 172544 74318 172553
rect 74262 172479 74318 172488
rect 74446 172544 74502 172553
rect 74446 172479 74502 172488
rect 74460 162858 74488 172479
rect 74448 162852 74500 162858
rect 74448 162794 74500 162800
rect 74448 153264 74500 153270
rect 74448 153206 74500 153212
rect 74460 145081 74488 153206
rect 74446 145072 74502 145081
rect 74446 145007 74502 145016
rect 74446 144936 74502 144945
rect 74446 144871 74502 144880
rect 74460 143546 74488 144871
rect 74448 143540 74500 143546
rect 74448 143482 74500 143488
rect 74448 133952 74500 133958
rect 74448 133894 74500 133900
rect 74460 125769 74488 133894
rect 74446 125760 74502 125769
rect 74446 125695 74502 125704
rect 74446 125624 74502 125633
rect 74446 125559 74502 125568
rect 74460 104854 74488 125559
rect 74448 104848 74500 104854
rect 74448 104790 74500 104796
rect 74448 95260 74500 95266
rect 74448 95202 74500 95208
rect 74460 66230 74488 95202
rect 74448 66224 74500 66230
rect 74448 66166 74500 66172
rect 74448 56636 74500 56642
rect 74448 56578 74500 56584
rect 74460 46918 74488 56578
rect 74448 46912 74500 46918
rect 74448 46854 74500 46860
rect 74448 37324 74500 37330
rect 74448 37266 74500 37272
rect 74460 27606 74488 37266
rect 74448 27600 74500 27606
rect 74448 27542 74500 27548
rect 74264 9716 74316 9722
rect 74264 9658 74316 9664
rect 73250 3768 73306 3777
rect 73250 3703 73306 3712
rect 74276 480 74304 9658
rect 74644 3913 74672 320062
rect 75104 316010 75132 320062
rect 75184 318300 75236 318306
rect 75184 318242 75236 318248
rect 74736 315982 75132 316010
rect 74736 4049 74764 315982
rect 75000 315920 75052 315926
rect 75000 315862 75052 315868
rect 75012 302394 75040 315862
rect 75000 302388 75052 302394
rect 75000 302330 75052 302336
rect 75000 299532 75052 299538
rect 75000 299474 75052 299480
rect 75012 299402 75040 299474
rect 75000 299396 75052 299402
rect 75000 299338 75052 299344
rect 74908 289876 74960 289882
rect 74908 289818 74960 289824
rect 74920 289746 74948 289818
rect 74908 289740 74960 289746
rect 74908 289682 74960 289688
rect 75000 280220 75052 280226
rect 75000 280162 75052 280168
rect 75012 280106 75040 280162
rect 75012 280078 75132 280106
rect 75104 270552 75132 280078
rect 75012 270524 75132 270552
rect 75012 260846 75040 270524
rect 75000 260840 75052 260846
rect 75000 260782 75052 260788
rect 75000 251252 75052 251258
rect 75000 251194 75052 251200
rect 75012 241505 75040 251194
rect 74814 241496 74870 241505
rect 74814 241431 74870 241440
rect 74998 241496 75054 241505
rect 74998 241431 75054 241440
rect 74828 231878 74856 241431
rect 74816 231872 74868 231878
rect 74816 231814 74868 231820
rect 75000 231872 75052 231878
rect 75000 231814 75052 231820
rect 75012 222193 75040 231814
rect 74814 222184 74870 222193
rect 74814 222119 74870 222128
rect 74998 222184 75054 222193
rect 74998 222119 75054 222128
rect 74828 212566 74856 222119
rect 74816 212560 74868 212566
rect 74816 212502 74868 212508
rect 75000 212560 75052 212566
rect 75000 212502 75052 212508
rect 75012 202881 75040 212502
rect 74814 202872 74870 202881
rect 74814 202807 74870 202816
rect 74998 202872 75054 202881
rect 74998 202807 75054 202816
rect 74828 193254 74856 202807
rect 74816 193248 74868 193254
rect 74816 193190 74868 193196
rect 75000 193248 75052 193254
rect 75000 193190 75052 193196
rect 75012 183569 75040 193190
rect 74814 183560 74870 183569
rect 74814 183495 74870 183504
rect 74998 183560 75054 183569
rect 74998 183495 75054 183504
rect 74828 173942 74856 183495
rect 74816 173936 74868 173942
rect 74816 173878 74868 173884
rect 75000 173936 75052 173942
rect 75000 173878 75052 173884
rect 75012 157434 75040 173878
rect 74920 157406 75040 157434
rect 74920 157298 74948 157406
rect 74920 157270 75040 157298
rect 75012 145081 75040 157270
rect 74998 145072 75054 145081
rect 74998 145007 75054 145016
rect 74998 144936 75054 144945
rect 74998 144871 75054 144880
rect 75012 143546 75040 144871
rect 75000 143540 75052 143546
rect 75000 143482 75052 143488
rect 75000 133952 75052 133958
rect 75000 133894 75052 133900
rect 75012 125769 75040 133894
rect 74998 125760 75054 125769
rect 74998 125695 75054 125704
rect 74998 125624 75054 125633
rect 74998 125559 75054 125568
rect 75012 122806 75040 125559
rect 75000 122800 75052 122806
rect 75000 122742 75052 122748
rect 75000 117292 75052 117298
rect 75000 117234 75052 117240
rect 75012 95418 75040 117234
rect 74920 95390 75040 95418
rect 74920 93922 74948 95390
rect 74920 93894 75040 93922
rect 75012 93838 75040 93894
rect 75000 93832 75052 93838
rect 75000 93774 75052 93780
rect 75000 84312 75052 84318
rect 75000 84254 75052 84260
rect 75012 84182 75040 84254
rect 75000 84176 75052 84182
rect 75000 84118 75052 84124
rect 75000 74588 75052 74594
rect 75000 74530 75052 74536
rect 75012 71126 75040 74530
rect 75000 71120 75052 71126
rect 75000 71062 75052 71068
rect 74816 66292 74868 66298
rect 74816 66234 74868 66240
rect 74828 64870 74856 66234
rect 74816 64864 74868 64870
rect 74816 64806 74868 64812
rect 74908 55276 74960 55282
rect 74908 55218 74960 55224
rect 74920 46918 74948 55218
rect 74908 46912 74960 46918
rect 74908 46854 74960 46860
rect 75092 46912 75144 46918
rect 75092 46854 75144 46860
rect 75104 45558 75132 46854
rect 75092 45552 75144 45558
rect 75092 45494 75144 45500
rect 75092 37256 75144 37262
rect 75092 37198 75144 37204
rect 75104 29782 75132 37198
rect 74816 29776 74868 29782
rect 74816 29718 74868 29724
rect 75092 29776 75144 29782
rect 75092 29718 75144 29724
rect 74828 27606 74856 29718
rect 74816 27600 74868 27606
rect 74816 27542 74868 27548
rect 74908 9716 74960 9722
rect 74908 9658 74960 9664
rect 74722 4040 74778 4049
rect 74722 3975 74778 3984
rect 74630 3904 74686 3913
rect 74630 3839 74686 3848
rect 74920 3262 74948 9658
rect 75196 4146 75224 318242
rect 75472 315926 75500 320062
rect 76300 317898 76328 320076
rect 76288 317892 76340 317898
rect 76288 317834 76340 317840
rect 76760 317762 76788 320076
rect 76748 317756 76800 317762
rect 76748 317698 76800 317704
rect 77220 317626 77248 320076
rect 77312 320062 77694 320090
rect 77772 320062 78154 320090
rect 78232 320062 78614 320090
rect 77208 317620 77260 317626
rect 77208 317562 77260 317568
rect 75460 315920 75512 315926
rect 75460 315862 75512 315868
rect 77208 28892 77260 28898
rect 77208 28834 77260 28840
rect 77220 19242 77248 28834
rect 77208 19236 77260 19242
rect 77208 19178 77260 19184
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 75460 3936 75512 3942
rect 75460 3878 75512 3884
rect 74908 3256 74960 3262
rect 74908 3198 74960 3204
rect 75472 480 75500 3878
rect 76656 3528 76708 3534
rect 76656 3470 76708 3476
rect 76668 480 76696 3470
rect 77312 3194 77340 320062
rect 77772 316010 77800 320062
rect 77944 317620 77996 317626
rect 77944 317562 77996 317568
rect 77404 315982 77800 316010
rect 77300 3188 77352 3194
rect 77300 3130 77352 3136
rect 77404 3058 77432 315982
rect 77576 315920 77628 315926
rect 77576 315862 77628 315868
rect 77588 309126 77616 315862
rect 77576 309120 77628 309126
rect 77576 309062 77628 309068
rect 77576 299532 77628 299538
rect 77576 299474 77628 299480
rect 77588 282946 77616 299474
rect 77576 282940 77628 282946
rect 77576 282882 77628 282888
rect 77576 270564 77628 270570
rect 77576 270506 77628 270512
rect 77588 260846 77616 270506
rect 77576 260840 77628 260846
rect 77576 260782 77628 260788
rect 77576 251252 77628 251258
rect 77576 251194 77628 251200
rect 77588 241482 77616 251194
rect 77588 241454 77708 241482
rect 77680 234666 77708 241454
rect 77668 234660 77720 234666
rect 77668 234602 77720 234608
rect 77576 234592 77628 234598
rect 77576 234534 77628 234540
rect 77588 222193 77616 234534
rect 77574 222184 77630 222193
rect 77574 222119 77630 222128
rect 77758 222184 77814 222193
rect 77758 222119 77814 222128
rect 77772 212566 77800 222119
rect 77576 212560 77628 212566
rect 77576 212502 77628 212508
rect 77760 212560 77812 212566
rect 77760 212502 77812 212508
rect 77588 202858 77616 212502
rect 77588 202830 77708 202858
rect 77680 196042 77708 202830
rect 77668 196036 77720 196042
rect 77668 195978 77720 195984
rect 77576 195968 77628 195974
rect 77576 195910 77628 195916
rect 77588 183546 77616 195910
rect 77496 183518 77616 183546
rect 77496 176730 77524 183518
rect 77484 176724 77536 176730
rect 77484 176666 77536 176672
rect 77576 176656 77628 176662
rect 77576 176598 77628 176604
rect 77588 157434 77616 176598
rect 77496 157406 77616 157434
rect 77496 157298 77524 157406
rect 77496 157270 77616 157298
rect 77588 135386 77616 157270
rect 77576 135380 77628 135386
rect 77576 135322 77628 135328
rect 77576 135244 77628 135250
rect 77576 135186 77628 135192
rect 77588 133906 77616 135186
rect 77588 133890 77708 133906
rect 77588 133884 77720 133890
rect 77588 133878 77668 133884
rect 77668 133826 77720 133832
rect 77852 133884 77904 133890
rect 77852 133826 77904 133832
rect 77680 133795 77708 133826
rect 77864 124273 77892 133826
rect 77482 124264 77538 124273
rect 77482 124199 77538 124208
rect 77850 124264 77906 124273
rect 77850 124199 77906 124208
rect 77496 124166 77524 124199
rect 77484 124160 77536 124166
rect 77484 124102 77536 124108
rect 77576 124160 77628 124166
rect 77576 124102 77628 124108
rect 77588 114510 77616 124102
rect 77576 114504 77628 114510
rect 77576 114446 77628 114452
rect 77576 104916 77628 104922
rect 77576 104858 77628 104864
rect 77588 99498 77616 104858
rect 77588 99470 77708 99498
rect 77680 99226 77708 99470
rect 77588 99198 77708 99226
rect 77588 67726 77616 99198
rect 77576 67720 77628 67726
rect 77576 67662 77628 67668
rect 77484 67652 77536 67658
rect 77484 67594 77536 67600
rect 77496 66230 77524 67594
rect 77484 66224 77536 66230
rect 77484 66166 77536 66172
rect 77484 48408 77536 48414
rect 77484 48350 77536 48356
rect 77496 46918 77524 48350
rect 77484 46912 77536 46918
rect 77484 46854 77536 46860
rect 77760 46912 77812 46918
rect 77760 46854 77812 46860
rect 77772 28898 77800 46854
rect 77760 28892 77812 28898
rect 77760 28834 77812 28840
rect 77760 19236 77812 19242
rect 77760 19178 77812 19184
rect 77772 9722 77800 19178
rect 77484 9716 77536 9722
rect 77484 9658 77536 9664
rect 77760 9716 77812 9722
rect 77760 9658 77812 9664
rect 77496 3262 77524 9658
rect 77956 3874 77984 317562
rect 78232 315926 78260 320062
rect 78968 317694 78996 320076
rect 78956 317688 79008 317694
rect 78956 317630 79008 317636
rect 78220 315920 78272 315926
rect 78220 315862 78272 315868
rect 79060 309194 79088 320198
rect 79324 318436 79376 318442
rect 79324 318378 79376 318384
rect 78864 309188 78916 309194
rect 78864 309130 78916 309136
rect 79048 309188 79100 309194
rect 79048 309130 79100 309136
rect 78876 292618 78904 309130
rect 78784 292590 78904 292618
rect 78784 292482 78812 292590
rect 78784 292454 78904 292482
rect 78876 263650 78904 292454
rect 78784 263622 78904 263650
rect 78784 263514 78812 263622
rect 78784 263486 78904 263514
rect 78876 244338 78904 263486
rect 78784 244310 78904 244338
rect 78784 244202 78812 244310
rect 78784 244174 78904 244202
rect 78876 225026 78904 244174
rect 78784 224998 78904 225026
rect 78784 224890 78812 224998
rect 78784 224862 78904 224890
rect 78876 205714 78904 224862
rect 78784 205686 78904 205714
rect 78784 205578 78812 205686
rect 78784 205550 78904 205578
rect 78876 186402 78904 205550
rect 78784 186374 78904 186402
rect 78784 186266 78812 186374
rect 78784 186238 78904 186266
rect 78876 167006 78904 186238
rect 78864 167000 78916 167006
rect 78864 166942 78916 166948
rect 78864 166864 78916 166870
rect 78864 166806 78916 166812
rect 78876 162858 78904 166806
rect 78864 162852 78916 162858
rect 78864 162794 78916 162800
rect 78864 153264 78916 153270
rect 78864 153206 78916 153212
rect 78876 144922 78904 153206
rect 78784 144894 78904 144922
rect 78784 140078 78812 144894
rect 78772 140072 78824 140078
rect 78772 140014 78824 140020
rect 78864 140004 78916 140010
rect 78864 139946 78916 139952
rect 78876 125769 78904 139946
rect 78862 125760 78918 125769
rect 78862 125695 78918 125704
rect 78770 125624 78826 125633
rect 78770 125559 78772 125568
rect 78824 125559 78826 125568
rect 78772 125530 78824 125536
rect 78864 125452 78916 125458
rect 78864 125394 78916 125400
rect 78876 106457 78904 125394
rect 78862 106448 78918 106457
rect 78862 106383 78918 106392
rect 78770 106312 78826 106321
rect 78770 106247 78826 106256
rect 78784 104854 78812 106247
rect 78772 104848 78824 104854
rect 78772 104790 78824 104796
rect 78956 95260 79008 95266
rect 78956 95202 79008 95208
rect 78968 85610 78996 95202
rect 78772 85604 78824 85610
rect 78772 85546 78824 85552
rect 78956 85604 79008 85610
rect 78956 85546 79008 85552
rect 78784 75954 78812 85546
rect 78772 75948 78824 75954
rect 78772 75890 78824 75896
rect 78864 75948 78916 75954
rect 78864 75890 78916 75896
rect 78876 38622 78904 75890
rect 78864 38616 78916 38622
rect 78864 38558 78916 38564
rect 78864 29028 78916 29034
rect 78864 28970 78916 28976
rect 78876 12458 78904 28970
rect 78784 12430 78904 12458
rect 78784 4078 78812 12430
rect 78772 4072 78824 4078
rect 78772 4014 78824 4020
rect 79048 4072 79100 4078
rect 79048 4014 79100 4020
rect 77944 3868 77996 3874
rect 77944 3810 77996 3816
rect 77484 3256 77536 3262
rect 77484 3198 77536 3204
rect 77852 3256 77904 3262
rect 77852 3198 77904 3204
rect 77392 3052 77444 3058
rect 77392 2994 77444 3000
rect 77864 480 77892 3198
rect 79060 480 79088 4014
rect 79336 4010 79364 318378
rect 79416 317960 79468 317966
rect 79416 317902 79468 317908
rect 79324 4004 79376 4010
rect 79324 3946 79376 3952
rect 79428 3806 79456 317902
rect 79888 317558 79916 320076
rect 80072 320062 80362 320090
rect 80440 320062 80822 320090
rect 80992 320062 81282 320090
rect 79876 317552 79928 317558
rect 79876 317494 79928 317500
rect 79416 3800 79468 3806
rect 79416 3742 79468 3748
rect 80072 2990 80100 320062
rect 80152 315988 80204 315994
rect 80152 315930 80204 315936
rect 80060 2984 80112 2990
rect 80060 2926 80112 2932
rect 80164 2922 80192 315930
rect 80440 301578 80468 320062
rect 80992 315994 81020 320062
rect 81728 317490 81756 320076
rect 81912 320062 82202 320090
rect 82280 320062 82570 320090
rect 83030 320062 83136 320090
rect 81716 317484 81768 317490
rect 81716 317426 81768 317432
rect 80980 315988 81032 315994
rect 80980 315930 81032 315936
rect 81532 315988 81584 315994
rect 81532 315930 81584 315936
rect 80428 301572 80480 301578
rect 80428 301514 80480 301520
rect 80244 296744 80296 296750
rect 80244 296686 80296 296692
rect 80256 288318 80284 296686
rect 80244 288312 80296 288318
rect 80244 288254 80296 288260
rect 80428 288244 80480 288250
rect 80428 288186 80480 288192
rect 80440 263514 80468 288186
rect 80348 263486 80468 263514
rect 80348 260846 80376 263486
rect 80336 260840 80388 260846
rect 80336 260782 80388 260788
rect 80428 260840 80480 260846
rect 80428 260782 80480 260788
rect 80440 244202 80468 260782
rect 80348 244174 80468 244202
rect 80348 231878 80376 244174
rect 80336 231872 80388 231878
rect 80336 231814 80388 231820
rect 80428 231872 80480 231878
rect 80428 231814 80480 231820
rect 80440 224890 80468 231814
rect 80348 224862 80468 224890
rect 80348 212566 80376 224862
rect 80336 212560 80388 212566
rect 80336 212502 80388 212508
rect 80428 212560 80480 212566
rect 80428 212502 80480 212508
rect 80440 205578 80468 212502
rect 80348 205550 80468 205578
rect 80348 202842 80376 205550
rect 80336 202836 80388 202842
rect 80336 202778 80388 202784
rect 80428 202836 80480 202842
rect 80428 202778 80480 202784
rect 80440 186266 80468 202778
rect 80348 186238 80468 186266
rect 80348 183530 80376 186238
rect 80336 183524 80388 183530
rect 80336 183466 80388 183472
rect 80428 183524 80480 183530
rect 80428 183466 80480 183472
rect 80440 166954 80468 183466
rect 80348 166926 80468 166954
rect 80348 157434 80376 166926
rect 80256 157406 80376 157434
rect 80256 157350 80284 157406
rect 80244 157344 80296 157350
rect 80244 157286 80296 157292
rect 80428 157344 80480 157350
rect 80428 157286 80480 157292
rect 80440 154562 80468 157286
rect 80336 154556 80388 154562
rect 80336 154498 80388 154504
rect 80428 154556 80480 154562
rect 80428 154498 80480 154504
rect 80348 138038 80376 154498
rect 80336 138032 80388 138038
rect 80336 137974 80388 137980
rect 80428 137964 80480 137970
rect 80428 137906 80480 137912
rect 80440 128330 80468 137906
rect 80348 128302 80468 128330
rect 80348 118726 80376 128302
rect 80336 118720 80388 118726
rect 80336 118662 80388 118668
rect 80428 118652 80480 118658
rect 80428 118594 80480 118600
rect 80440 109018 80468 118594
rect 80348 108990 80468 109018
rect 80348 100042 80376 108990
rect 80348 100014 80468 100042
rect 80440 89706 80468 100014
rect 80348 89678 80468 89706
rect 80348 70446 80376 89678
rect 80336 70440 80388 70446
rect 80336 70382 80388 70388
rect 80336 70304 80388 70310
rect 80336 70246 80388 70252
rect 80348 60738 80376 70246
rect 80256 60722 80376 60738
rect 80244 60716 80376 60722
rect 80296 60710 80376 60716
rect 80428 60716 80480 60722
rect 80244 60658 80296 60664
rect 80428 60658 80480 60664
rect 80440 51082 80468 60658
rect 80348 51054 80468 51082
rect 80348 41426 80376 51054
rect 80256 41410 80376 41426
rect 80244 41404 80376 41410
rect 80296 41398 80376 41404
rect 80428 41404 80480 41410
rect 80244 41346 80296 41352
rect 80428 41346 80480 41352
rect 80440 31770 80468 41346
rect 80348 31742 80468 31770
rect 80348 22114 80376 31742
rect 80256 22098 80376 22114
rect 80244 22092 80376 22098
rect 80296 22086 80376 22092
rect 80428 22092 80480 22098
rect 80244 22034 80296 22040
rect 80428 22034 80480 22040
rect 80440 12050 80468 22034
rect 80440 12022 80560 12050
rect 80532 11778 80560 12022
rect 80440 11750 80560 11778
rect 80440 4826 80468 11750
rect 80428 4820 80480 4826
rect 80428 4762 80480 4768
rect 80244 4140 80296 4146
rect 80244 4082 80296 4088
rect 80152 2916 80204 2922
rect 80152 2858 80204 2864
rect 80256 480 80284 4082
rect 81440 3732 81492 3738
rect 81440 3674 81492 3680
rect 81452 480 81480 3674
rect 81544 3466 81572 315930
rect 81912 299554 81940 320062
rect 82084 318504 82136 318510
rect 82084 318446 82136 318452
rect 81820 299526 81940 299554
rect 81820 293434 81848 299526
rect 81728 293406 81848 293434
rect 81728 283626 81756 293406
rect 81716 283620 81768 283626
rect 81716 283562 81768 283568
rect 81716 278792 81768 278798
rect 81714 278760 81716 278769
rect 81768 278760 81770 278769
rect 81714 278695 81770 278704
rect 81898 270464 81954 270473
rect 81898 270399 81954 270408
rect 81912 263514 81940 270399
rect 81820 263486 81940 263514
rect 81820 251258 81848 263486
rect 81808 251252 81860 251258
rect 81808 251194 81860 251200
rect 81900 251252 81952 251258
rect 81900 251194 81952 251200
rect 81912 244202 81940 251194
rect 81820 244174 81940 244202
rect 81820 231878 81848 244174
rect 81808 231872 81860 231878
rect 81808 231814 81860 231820
rect 81900 231872 81952 231878
rect 81900 231814 81952 231820
rect 81912 224890 81940 231814
rect 81820 224862 81940 224890
rect 81820 212566 81848 224862
rect 81808 212560 81860 212566
rect 81808 212502 81860 212508
rect 81900 212560 81952 212566
rect 81900 212502 81952 212508
rect 81912 205578 81940 212502
rect 81820 205550 81940 205578
rect 81820 193254 81848 205550
rect 81808 193248 81860 193254
rect 81808 193190 81860 193196
rect 81900 193248 81952 193254
rect 81900 193190 81952 193196
rect 81912 186266 81940 193190
rect 81820 186238 81940 186266
rect 81820 173942 81848 186238
rect 81808 173936 81860 173942
rect 81808 173878 81860 173884
rect 81900 173936 81952 173942
rect 81900 173878 81952 173884
rect 81912 166954 81940 173878
rect 81820 166926 81940 166954
rect 81820 157434 81848 166926
rect 81728 157406 81848 157434
rect 81728 157350 81756 157406
rect 81716 157344 81768 157350
rect 81716 157286 81768 157292
rect 81900 157344 81952 157350
rect 81900 157286 81952 157292
rect 81912 154562 81940 157286
rect 81808 154556 81860 154562
rect 81808 154498 81860 154504
rect 81900 154556 81952 154562
rect 81900 154498 81952 154504
rect 81820 138038 81848 154498
rect 81808 138032 81860 138038
rect 81808 137974 81860 137980
rect 81900 137964 81952 137970
rect 81900 137906 81952 137912
rect 81912 128330 81940 137906
rect 81820 128302 81940 128330
rect 81820 118726 81848 128302
rect 81808 118720 81860 118726
rect 81808 118662 81860 118668
rect 81900 118652 81952 118658
rect 81900 118594 81952 118600
rect 81912 109018 81940 118594
rect 81820 108990 81940 109018
rect 81820 100042 81848 108990
rect 81820 100014 81940 100042
rect 81912 89706 81940 100014
rect 81728 89678 81940 89706
rect 81728 80170 81756 89678
rect 81716 80164 81768 80170
rect 81716 80106 81768 80112
rect 81624 80028 81676 80034
rect 81624 79970 81676 79976
rect 81636 77246 81664 79970
rect 81624 77240 81676 77246
rect 81624 77182 81676 77188
rect 81716 70304 81768 70310
rect 81716 70246 81768 70252
rect 81728 60722 81756 70246
rect 81716 60716 81768 60722
rect 81716 60658 81768 60664
rect 81900 60716 81952 60722
rect 81900 60658 81952 60664
rect 81912 51082 81940 60658
rect 81820 51054 81940 51082
rect 81820 41426 81848 51054
rect 81728 41410 81848 41426
rect 81716 41404 81848 41410
rect 81768 41398 81848 41404
rect 81900 41404 81952 41410
rect 81716 41346 81768 41352
rect 81900 41346 81952 41352
rect 81912 29034 81940 41346
rect 81808 29028 81860 29034
rect 81808 28970 81860 28976
rect 81900 29028 81952 29034
rect 81900 28970 81952 28976
rect 81820 22114 81848 28970
rect 81728 22098 81848 22114
rect 81716 22092 81848 22098
rect 81768 22086 81848 22092
rect 81900 22092 81952 22098
rect 81716 22034 81768 22040
rect 81900 22034 81952 22040
rect 81912 12050 81940 22034
rect 81912 12022 82032 12050
rect 82004 11778 82032 12022
rect 81912 11750 82032 11778
rect 81912 3806 81940 11750
rect 82096 4146 82124 318446
rect 82176 317552 82228 317558
rect 82176 317494 82228 317500
rect 82084 4140 82136 4146
rect 82084 4082 82136 4088
rect 81900 3800 81952 3806
rect 81900 3742 81952 3748
rect 82188 3534 82216 317494
rect 82280 315994 82308 320062
rect 82728 318368 82780 318374
rect 82728 318310 82780 318316
rect 82268 315988 82320 315994
rect 82268 315930 82320 315936
rect 82740 3738 82768 318310
rect 82912 315716 82964 315722
rect 82912 315658 82964 315664
rect 82924 4078 82952 315658
rect 82912 4072 82964 4078
rect 82912 4014 82964 4020
rect 82728 3732 82780 3738
rect 82728 3674 82780 3680
rect 82176 3528 82228 3534
rect 82176 3470 82228 3476
rect 81532 3460 81584 3466
rect 81532 3402 81584 3408
rect 82636 3460 82688 3466
rect 82636 3402 82688 3408
rect 82648 480 82676 3402
rect 83108 2854 83136 320062
rect 83476 317966 83504 320076
rect 83568 320062 83950 320090
rect 83464 317960 83516 317966
rect 83464 317902 83516 317908
rect 83568 315722 83596 320062
rect 84292 315988 84344 315994
rect 84292 315930 84344 315936
rect 83556 315716 83608 315722
rect 83556 315658 83608 315664
rect 83832 4140 83884 4146
rect 83832 4082 83884 4088
rect 83096 2848 83148 2854
rect 83096 2790 83148 2796
rect 83844 480 83872 4082
rect 84304 3670 84332 315930
rect 84292 3664 84344 3670
rect 84292 3606 84344 3612
rect 84396 3602 84424 320076
rect 84488 320062 84870 320090
rect 84488 315994 84516 320062
rect 84844 317824 84896 317830
rect 84844 317766 84896 317772
rect 84476 315988 84528 315994
rect 84476 315930 84528 315936
rect 84856 4146 84884 317766
rect 85316 317626 85344 320076
rect 85488 317960 85540 317966
rect 85488 317902 85540 317908
rect 85304 317620 85356 317626
rect 85304 317562 85356 317568
rect 85500 4146 85528 317902
rect 85580 315988 85632 315994
rect 85580 315930 85632 315936
rect 84844 4140 84896 4146
rect 84844 4082 84896 4088
rect 84936 4140 84988 4146
rect 84936 4082 84988 4088
rect 85488 4140 85540 4146
rect 85488 4082 85540 4088
rect 84384 3596 84436 3602
rect 84384 3538 84436 3544
rect 84948 480 84976 4082
rect 85592 4010 85620 315930
rect 85580 4004 85632 4010
rect 85580 3946 85632 3952
rect 85776 3942 85804 320076
rect 86144 320062 86250 320090
rect 86328 320062 86618 320090
rect 86144 309194 86172 320062
rect 86224 317484 86276 317490
rect 86224 317426 86276 317432
rect 86040 309188 86092 309194
rect 86040 309130 86092 309136
rect 86132 309188 86184 309194
rect 86132 309130 86184 309136
rect 86052 307766 86080 309130
rect 86040 307760 86092 307766
rect 86040 307702 86092 307708
rect 85948 298172 86000 298178
rect 85948 298114 86000 298120
rect 85960 292670 85988 298114
rect 85948 292664 86000 292670
rect 85948 292606 86000 292612
rect 85948 292528 86000 292534
rect 85948 292470 86000 292476
rect 85960 278866 85988 292470
rect 85856 278860 85908 278866
rect 85856 278802 85908 278808
rect 85948 278860 86000 278866
rect 85948 278802 86000 278808
rect 85868 278730 85896 278802
rect 85856 278724 85908 278730
rect 85856 278666 85908 278672
rect 86040 278724 86092 278730
rect 86040 278666 86092 278672
rect 86052 277370 86080 278666
rect 86040 277364 86092 277370
rect 86040 277306 86092 277312
rect 86132 277364 86184 277370
rect 86132 277306 86184 277312
rect 86144 251190 86172 277306
rect 85948 251184 86000 251190
rect 85948 251126 86000 251132
rect 86132 251184 86184 251190
rect 86132 251126 86184 251132
rect 85960 234666 85988 251126
rect 85948 234660 86000 234666
rect 85948 234602 86000 234608
rect 85856 234592 85908 234598
rect 85856 234534 85908 234540
rect 85868 212537 85896 234534
rect 85854 212528 85910 212537
rect 85854 212463 85910 212472
rect 86130 212528 86186 212537
rect 86130 212463 86186 212472
rect 86144 202910 86172 212463
rect 85948 202904 86000 202910
rect 85948 202846 86000 202852
rect 86132 202904 86184 202910
rect 86132 202846 86184 202852
rect 85960 196042 85988 202846
rect 85948 196036 86000 196042
rect 85948 195978 86000 195984
rect 85856 195968 85908 195974
rect 85856 195910 85908 195916
rect 85868 193225 85896 195910
rect 85854 193216 85910 193225
rect 85854 193151 85910 193160
rect 86130 193216 86186 193225
rect 86130 193151 86186 193160
rect 86144 183598 86172 193151
rect 85948 183592 86000 183598
rect 85948 183534 86000 183540
rect 86132 183592 86184 183598
rect 86132 183534 86184 183540
rect 85960 176730 85988 183534
rect 85948 176724 86000 176730
rect 85948 176666 86000 176672
rect 85856 176656 85908 176662
rect 85856 176598 85908 176604
rect 85868 157350 85896 176598
rect 85856 157344 85908 157350
rect 85856 157286 85908 157292
rect 86040 157344 86092 157350
rect 86040 157286 86092 157292
rect 86052 147778 86080 157286
rect 86052 147750 86172 147778
rect 86144 144945 86172 147750
rect 85946 144936 86002 144945
rect 85856 144900 85908 144906
rect 85946 144871 85948 144880
rect 85856 144842 85908 144848
rect 86000 144871 86002 144880
rect 86130 144936 86186 144945
rect 86130 144871 86186 144880
rect 85948 144842 86000 144848
rect 85868 135289 85896 144842
rect 85854 135280 85910 135289
rect 85854 135215 85910 135224
rect 86038 135280 86094 135289
rect 86038 135215 86094 135224
rect 86052 128466 86080 135215
rect 86052 128438 86172 128466
rect 86144 125633 86172 128438
rect 85946 125624 86002 125633
rect 85856 125588 85908 125594
rect 85946 125559 85948 125568
rect 85856 125530 85908 125536
rect 86000 125559 86002 125568
rect 86130 125624 86186 125633
rect 86130 125559 86186 125568
rect 85948 125530 86000 125536
rect 85868 115977 85896 125530
rect 85854 115968 85910 115977
rect 85854 115903 85910 115912
rect 86038 115968 86094 115977
rect 86038 115903 86094 115912
rect 86052 106350 86080 115903
rect 85948 106344 86000 106350
rect 85948 106286 86000 106292
rect 86040 106344 86092 106350
rect 86040 106286 86092 106292
rect 85960 104854 85988 106286
rect 85948 104848 86000 104854
rect 85948 104790 86000 104796
rect 86040 95260 86092 95266
rect 86040 95202 86092 95208
rect 86052 89706 86080 95202
rect 85960 89678 86080 89706
rect 85960 86970 85988 89678
rect 85948 86964 86000 86970
rect 85948 86906 86000 86912
rect 85856 77308 85908 77314
rect 85856 77250 85908 77256
rect 85868 29034 85896 77250
rect 85856 29028 85908 29034
rect 85856 28970 85908 28976
rect 85948 28892 86000 28898
rect 85948 28834 86000 28840
rect 85960 26246 85988 28834
rect 85948 26240 86000 26246
rect 85948 26182 86000 26188
rect 86040 26240 86092 26246
rect 86040 26182 86092 26188
rect 85764 3936 85816 3942
rect 85764 3878 85816 3884
rect 86052 3330 86080 26182
rect 86236 3398 86264 317426
rect 86328 315994 86356 320062
rect 87064 318306 87092 320076
rect 87524 318442 87552 320076
rect 87512 318436 87564 318442
rect 87512 318378 87564 318384
rect 87052 318300 87104 318306
rect 87052 318242 87104 318248
rect 87984 318170 88012 320076
rect 87972 318164 88024 318170
rect 87972 318106 88024 318112
rect 87604 318096 87656 318102
rect 87604 318038 87656 318044
rect 86316 315988 86368 315994
rect 86316 315930 86368 315936
rect 87616 3874 87644 318038
rect 88248 318028 88300 318034
rect 88248 317970 88300 317976
rect 87604 3868 87656 3874
rect 87604 3810 87656 3816
rect 88260 3602 88288 317970
rect 88444 317490 88472 320076
rect 88904 317558 88932 320076
rect 88892 317552 88944 317558
rect 88892 317494 88944 317500
rect 88432 317484 88484 317490
rect 88432 317426 88484 317432
rect 88996 316010 89024 320198
rect 89824 318102 89852 320076
rect 90192 318510 90220 320076
rect 90180 318504 90232 318510
rect 90180 318446 90232 318452
rect 90652 318374 90680 320076
rect 90640 318368 90692 318374
rect 90640 318310 90692 318316
rect 89812 318096 89864 318102
rect 89812 318038 89864 318044
rect 89628 317892 89680 317898
rect 89628 317834 89680 317840
rect 88444 315982 89024 316010
rect 87328 3596 87380 3602
rect 87328 3538 87380 3544
rect 88248 3596 88300 3602
rect 88248 3538 88300 3544
rect 86224 3392 86276 3398
rect 86224 3334 86276 3340
rect 86040 3324 86092 3330
rect 86040 3266 86092 3272
rect 86132 3052 86184 3058
rect 86132 2994 86184 3000
rect 86144 480 86172 2994
rect 87340 480 87368 3538
rect 88444 3262 88472 315982
rect 89640 4146 89668 317834
rect 91008 317620 91060 317626
rect 91008 317562 91060 317568
rect 90364 317484 90416 317490
rect 90364 317426 90416 317432
rect 90376 4826 90404 317426
rect 90364 4820 90416 4826
rect 90364 4762 90416 4768
rect 88524 4140 88576 4146
rect 88524 4082 88576 4088
rect 89628 4140 89680 4146
rect 89628 4082 89680 4088
rect 88432 3256 88484 3262
rect 88432 3198 88484 3204
rect 88536 480 88564 4082
rect 89720 3868 89772 3874
rect 89720 3810 89772 3816
rect 89732 480 89760 3810
rect 91020 626 91048 317562
rect 91112 317490 91140 320076
rect 91572 317830 91600 320076
rect 92032 317966 92060 320076
rect 92506 320062 92704 320090
rect 92020 317960 92072 317966
rect 92020 317902 92072 317908
rect 91560 317824 91612 317830
rect 91560 317766 91612 317772
rect 92388 317552 92440 317558
rect 92388 317494 92440 317500
rect 91100 317484 91152 317490
rect 91100 317426 91152 317432
rect 90928 598 91048 626
rect 92400 610 92428 317494
rect 92572 315988 92624 315994
rect 92572 315930 92624 315936
rect 92584 3874 92612 315930
rect 92572 3868 92624 3874
rect 92572 3810 92624 3816
rect 92676 3058 92704 320062
rect 92952 318034 92980 320076
rect 92940 318028 92992 318034
rect 92940 317970 92992 317976
rect 93412 317898 93440 320076
rect 93504 320062 93794 320090
rect 93400 317892 93452 317898
rect 93400 317834 93452 317840
rect 93504 315994 93532 320062
rect 94240 317626 94268 320076
rect 94228 317620 94280 317626
rect 94228 317562 94280 317568
rect 94700 317558 94728 320076
rect 94688 317552 94740 317558
rect 94688 317494 94740 317500
rect 95160 317490 95188 320076
rect 95344 320062 95634 320090
rect 95804 320062 96094 320090
rect 93768 317484 93820 317490
rect 93768 317426 93820 317432
rect 95148 317484 95200 317490
rect 95148 317426 95200 317432
rect 93492 315988 93544 315994
rect 93492 315930 93544 315936
rect 93780 4146 93808 317426
rect 93308 4140 93360 4146
rect 93308 4082 93360 4088
rect 93768 4140 93820 4146
rect 93768 4082 93820 4088
rect 92664 3052 92716 3058
rect 92664 2994 92716 3000
rect 92112 604 92164 610
rect 90928 480 90956 598
rect 92112 546 92164 552
rect 92388 604 92440 610
rect 92388 546 92440 552
rect 92124 480 92152 546
rect 93320 480 93348 4082
rect 95344 3874 95372 320062
rect 95804 316010 95832 320062
rect 95436 315982 95832 316010
rect 95436 309126 95464 315982
rect 95424 309120 95476 309126
rect 95424 309062 95476 309068
rect 95700 299532 95752 299538
rect 95700 299474 95752 299480
rect 95712 285002 95740 299474
rect 95620 284974 95740 285002
rect 95620 280158 95648 284974
rect 95608 280152 95660 280158
rect 95608 280094 95660 280100
rect 95700 270564 95752 270570
rect 95700 270506 95752 270512
rect 95712 263514 95740 270506
rect 95620 263486 95740 263514
rect 95620 260846 95648 263486
rect 95608 260840 95660 260846
rect 95608 260782 95660 260788
rect 95700 251252 95752 251258
rect 95700 251194 95752 251200
rect 95712 244202 95740 251194
rect 95620 244174 95740 244202
rect 95620 241505 95648 244174
rect 95422 241496 95478 241505
rect 95422 241431 95478 241440
rect 95606 241496 95662 241505
rect 95606 241431 95662 241440
rect 95436 231878 95464 241431
rect 95424 231872 95476 231878
rect 95424 231814 95476 231820
rect 95700 231872 95752 231878
rect 95700 231814 95752 231820
rect 95712 224890 95740 231814
rect 95620 224862 95740 224890
rect 95620 222193 95648 224862
rect 95422 222184 95478 222193
rect 95422 222119 95478 222128
rect 95606 222184 95662 222193
rect 95606 222119 95662 222128
rect 95436 212566 95464 222119
rect 95424 212560 95476 212566
rect 95424 212502 95476 212508
rect 95700 212560 95752 212566
rect 95700 212502 95752 212508
rect 95712 205578 95740 212502
rect 95620 205550 95740 205578
rect 95620 202881 95648 205550
rect 95422 202872 95478 202881
rect 95422 202807 95478 202816
rect 95606 202872 95662 202881
rect 95606 202807 95662 202816
rect 95436 193254 95464 202807
rect 95424 193248 95476 193254
rect 95424 193190 95476 193196
rect 95700 193248 95752 193254
rect 95700 193190 95752 193196
rect 95712 186266 95740 193190
rect 95620 186238 95740 186266
rect 95620 183569 95648 186238
rect 95422 183560 95478 183569
rect 95422 183495 95478 183504
rect 95606 183560 95662 183569
rect 95606 183495 95662 183504
rect 95436 173942 95464 183495
rect 95424 173936 95476 173942
rect 95424 173878 95476 173884
rect 95700 173936 95752 173942
rect 95700 173878 95752 173884
rect 95712 166954 95740 173878
rect 95620 166926 95740 166954
rect 95620 164218 95648 166926
rect 95424 164212 95476 164218
rect 95424 164154 95476 164160
rect 95608 164212 95660 164218
rect 95608 164154 95660 164160
rect 95436 154601 95464 164154
rect 95422 154592 95478 154601
rect 95422 154527 95478 154536
rect 95698 154592 95754 154601
rect 95698 154527 95754 154536
rect 95712 147642 95740 154527
rect 95620 147614 95740 147642
rect 95620 140026 95648 147614
rect 95436 139998 95648 140026
rect 95436 135289 95464 139998
rect 95422 135280 95478 135289
rect 95422 135215 95478 135224
rect 95698 135280 95754 135289
rect 95698 135215 95754 135224
rect 95712 128330 95740 135215
rect 95620 128302 95740 128330
rect 95620 120714 95648 128302
rect 95436 120686 95648 120714
rect 95436 115977 95464 120686
rect 95422 115968 95478 115977
rect 95422 115903 95478 115912
rect 95698 115968 95754 115977
rect 95698 115903 95754 115912
rect 95712 109018 95740 115903
rect 95620 108990 95740 109018
rect 95620 101402 95648 108990
rect 95436 101374 95648 101402
rect 95436 96665 95464 101374
rect 95422 96656 95478 96665
rect 95422 96591 95478 96600
rect 95698 96656 95754 96665
rect 95698 96591 95754 96600
rect 95712 89706 95740 96591
rect 95528 89678 95740 89706
rect 95528 86970 95556 89678
rect 95516 86964 95568 86970
rect 95516 86906 95568 86912
rect 95424 77308 95476 77314
rect 95424 77250 95476 77256
rect 95436 77178 95464 77250
rect 95424 77172 95476 77178
rect 95424 77114 95476 77120
rect 95516 70304 95568 70310
rect 95516 70246 95568 70252
rect 95528 60722 95556 70246
rect 95516 60716 95568 60722
rect 95516 60658 95568 60664
rect 95700 60716 95752 60722
rect 95700 60658 95752 60664
rect 95712 57934 95740 60658
rect 95700 57928 95752 57934
rect 95700 57870 95752 57876
rect 95608 48340 95660 48346
rect 95608 48282 95660 48288
rect 95620 41426 95648 48282
rect 95528 41410 95648 41426
rect 95516 41404 95648 41410
rect 95568 41398 95648 41404
rect 95700 41404 95752 41410
rect 95516 41346 95568 41352
rect 95700 41346 95752 41352
rect 95712 38622 95740 41346
rect 95700 38616 95752 38622
rect 95700 38558 95752 38564
rect 95608 29028 95660 29034
rect 95608 28970 95660 28976
rect 95620 22114 95648 28970
rect 95528 22098 95648 22114
rect 95516 22092 95648 22098
rect 95568 22086 95648 22092
rect 95700 22092 95752 22098
rect 95516 22034 95568 22040
rect 95700 22034 95752 22040
rect 95712 19310 95740 22034
rect 95700 19304 95752 19310
rect 95700 19246 95752 19252
rect 95700 9716 95752 9722
rect 95700 9658 95752 9664
rect 94504 3868 94556 3874
rect 94504 3810 94556 3816
rect 95332 3868 95384 3874
rect 95332 3810 95384 3816
rect 94516 480 94544 3810
rect 95712 2854 95740 9658
rect 96540 4146 96568 320076
rect 97000 317490 97028 320076
rect 97460 317558 97488 320076
rect 97448 317552 97500 317558
rect 97448 317494 97500 317500
rect 96988 317484 97040 317490
rect 96988 317426 97040 317432
rect 97724 317484 97776 317490
rect 97724 317426 97776 317432
rect 96528 4140 96580 4146
rect 96528 4082 96580 4088
rect 96896 4140 96948 4146
rect 96896 4082 96948 4088
rect 95424 2848 95476 2854
rect 95424 2790 95476 2796
rect 95700 2848 95752 2854
rect 95700 2790 95752 2796
rect 95436 610 95464 2790
rect 95424 604 95476 610
rect 95424 546 95476 552
rect 95700 604 95752 610
rect 95700 546 95752 552
rect 95712 480 95740 546
rect 96908 480 96936 4082
rect 97736 3346 97764 317426
rect 97828 3466 97856 320076
rect 98288 317898 98316 320076
rect 98748 318102 98776 320076
rect 98736 318096 98788 318102
rect 98736 318038 98788 318044
rect 98276 317892 98328 317898
rect 98276 317834 98328 317840
rect 99208 317762 99236 320076
rect 99668 318714 99696 320076
rect 99656 318708 99708 318714
rect 99656 318650 99708 318656
rect 100116 317892 100168 317898
rect 100116 317834 100168 317840
rect 99196 317756 99248 317762
rect 99196 317698 99248 317704
rect 100024 317756 100076 317762
rect 100024 317698 100076 317704
rect 97908 317552 97960 317558
rect 97908 317494 97960 317500
rect 97920 4146 97948 317494
rect 100036 4146 100064 317698
rect 97908 4140 97960 4146
rect 97908 4082 97960 4088
rect 99288 4140 99340 4146
rect 99288 4082 99340 4088
rect 100024 4140 100076 4146
rect 100024 4082 100076 4088
rect 97816 3460 97868 3466
rect 97816 3402 97868 3408
rect 97736 3318 98132 3346
rect 98104 480 98132 3318
rect 99300 480 99328 4082
rect 100128 3534 100156 317834
rect 100496 317540 100524 320198
rect 100588 317694 100616 320076
rect 101048 317762 101076 320076
rect 101784 318050 101812 320198
rect 101890 320062 102088 320090
rect 101784 318022 101996 318050
rect 101036 317756 101088 317762
rect 101036 317698 101088 317704
rect 100576 317688 100628 317694
rect 100576 317630 100628 317636
rect 100496 317512 100708 317540
rect 100680 3602 100708 317512
rect 100668 3596 100720 3602
rect 100668 3538 100720 3544
rect 101968 3534 101996 318022
rect 100116 3528 100168 3534
rect 100116 3470 100168 3476
rect 101588 3528 101640 3534
rect 101588 3470 101640 3476
rect 101956 3528 102008 3534
rect 101956 3470 102008 3476
rect 100484 3460 100536 3466
rect 100484 3402 100536 3408
rect 100496 480 100524 3402
rect 101600 480 101628 3470
rect 102060 3466 102088 320062
rect 102336 317626 102364 320076
rect 102796 318102 102824 320076
rect 103270 320062 103468 320090
rect 102416 318096 102468 318102
rect 102416 318038 102468 318044
rect 102784 318096 102836 318102
rect 102784 318038 102836 318044
rect 103336 318096 103388 318102
rect 103336 318038 103388 318044
rect 102324 317620 102376 317626
rect 102324 317562 102376 317568
rect 102048 3460 102100 3466
rect 102048 3402 102100 3408
rect 102428 3346 102456 318038
rect 102784 317756 102836 317762
rect 102784 317698 102836 317704
rect 102796 3670 102824 317698
rect 102784 3664 102836 3670
rect 102784 3606 102836 3612
rect 102428 3318 102824 3346
rect 102796 480 102824 3318
rect 103348 3194 103376 318038
rect 103440 3262 103468 320062
rect 103716 317490 103744 320076
rect 104544 318050 104572 320198
rect 104650 320062 104848 320090
rect 104544 318022 104664 318050
rect 104164 317688 104216 317694
rect 104164 317630 104216 317636
rect 103704 317484 103756 317490
rect 103704 317426 103756 317432
rect 103980 4140 104032 4146
rect 103980 4082 104032 4088
rect 103428 3256 103480 3262
rect 103428 3198 103480 3204
rect 103336 3188 103388 3194
rect 103336 3130 103388 3136
rect 103992 480 104020 4082
rect 104176 3126 104204 317630
rect 104256 317620 104308 317626
rect 104256 317562 104308 317568
rect 104268 3398 104296 317562
rect 104636 4146 104664 318022
rect 104716 317484 104768 317490
rect 104716 317426 104768 317432
rect 104624 4140 104676 4146
rect 104624 4082 104676 4088
rect 104728 3738 104756 317426
rect 104820 4078 104848 320062
rect 105004 318102 105032 320076
rect 105478 320062 105860 320090
rect 105938 320062 106228 320090
rect 105176 318708 105228 318714
rect 105176 318650 105228 318656
rect 104992 318096 105044 318102
rect 104992 318038 105044 318044
rect 104808 4072 104860 4078
rect 104808 4014 104860 4020
rect 104716 3732 104768 3738
rect 104716 3674 104768 3680
rect 104256 3392 104308 3398
rect 104256 3334 104308 3340
rect 104164 3120 104216 3126
rect 104164 3062 104216 3068
rect 105188 480 105216 318650
rect 105728 318096 105780 318102
rect 105728 318038 105780 318044
rect 105740 316418 105768 318038
rect 105832 316554 105860 320062
rect 105832 316526 106136 316554
rect 105740 316390 106044 316418
rect 106016 3330 106044 316390
rect 106108 4010 106136 316526
rect 106096 4004 106148 4010
rect 106096 3946 106148 3952
rect 106200 3874 106228 320062
rect 106384 317626 106412 320076
rect 106844 317762 106872 320076
rect 107304 318306 107332 320076
rect 107292 318300 107344 318306
rect 107292 318242 107344 318248
rect 107764 318102 107792 320076
rect 107752 318096 107804 318102
rect 107752 318038 107804 318044
rect 108224 317762 108252 320076
rect 108592 318442 108620 320076
rect 108580 318436 108632 318442
rect 108580 318378 108632 318384
rect 108856 318096 108908 318102
rect 108856 318038 108908 318044
rect 106832 317756 106884 317762
rect 106832 317698 106884 317704
rect 107476 317756 107528 317762
rect 107476 317698 107528 317704
rect 108212 317756 108264 317762
rect 108212 317698 108264 317704
rect 106372 317620 106424 317626
rect 106372 317562 106424 317568
rect 106188 3868 106240 3874
rect 106188 3810 106240 3816
rect 107488 3806 107516 317698
rect 107568 317620 107620 317626
rect 107568 317562 107620 317568
rect 107580 3942 107608 317562
rect 107568 3936 107620 3942
rect 107568 3878 107620 3884
rect 107476 3800 107528 3806
rect 107476 3742 107528 3748
rect 108764 3664 108816 3670
rect 108764 3606 108816 3612
rect 106372 3596 106424 3602
rect 106372 3538 106424 3544
rect 106004 3324 106056 3330
rect 106004 3266 106056 3272
rect 106384 480 106412 3538
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 107580 480 107608 3062
rect 108776 480 108804 3606
rect 108868 2854 108896 318038
rect 108948 317756 109000 317762
rect 108948 317698 109000 317704
rect 108960 3738 108988 317698
rect 109052 317490 109080 320076
rect 109512 317558 109540 320076
rect 109986 320062 110276 320090
rect 109500 317552 109552 317558
rect 109500 317494 109552 317500
rect 110144 317552 110196 317558
rect 110144 317494 110196 317500
rect 109040 317484 109092 317490
rect 109040 317426 109092 317432
rect 108948 3732 109000 3738
rect 108948 3674 109000 3680
rect 110156 3670 110184 317494
rect 110144 3664 110196 3670
rect 110144 3606 110196 3612
rect 110248 3602 110276 320062
rect 110432 318034 110460 320076
rect 110420 318028 110472 318034
rect 110420 317970 110472 317976
rect 110892 317490 110920 320076
rect 111366 320062 111748 320090
rect 110328 317484 110380 317490
rect 110328 317426 110380 317432
rect 110880 317484 110932 317490
rect 110880 317426 110932 317432
rect 111616 317484 111668 317490
rect 111616 317426 111668 317432
rect 110236 3596 110288 3602
rect 110236 3538 110288 3544
rect 109960 3528 110012 3534
rect 109960 3470 110012 3476
rect 108856 2848 108908 2854
rect 108856 2790 108908 2796
rect 109972 480 110000 3470
rect 110340 3126 110368 317426
rect 111156 3460 111208 3466
rect 111156 3402 111208 3408
rect 110328 3120 110380 3126
rect 110328 3062 110380 3068
rect 111168 480 111196 3402
rect 111628 2922 111656 317426
rect 111720 3534 111748 320062
rect 111812 318578 111840 320076
rect 111800 318572 111852 318578
rect 111800 318514 111852 318520
rect 112272 317490 112300 320076
rect 112654 320062 113036 320090
rect 113008 317642 113036 320062
rect 113100 317830 113128 320076
rect 113088 317824 113140 317830
rect 113088 317766 113140 317772
rect 113008 317614 113128 317642
rect 112260 317484 112312 317490
rect 112260 317426 112312 317432
rect 112996 317484 113048 317490
rect 112996 317426 113048 317432
rect 111708 3528 111760 3534
rect 111708 3470 111760 3476
rect 113008 3466 113036 317426
rect 112996 3460 113048 3466
rect 112996 3402 113048 3408
rect 112352 3392 112404 3398
rect 112352 3334 112404 3340
rect 111616 2916 111668 2922
rect 111616 2858 111668 2864
rect 112364 480 112392 3334
rect 113100 2990 113128 317614
rect 113560 317490 113588 320076
rect 114034 320062 114324 320090
rect 113548 317484 113600 317490
rect 113548 317426 113600 317432
rect 114296 3194 114324 320062
rect 114376 317484 114428 317490
rect 114376 317426 114428 317432
rect 113548 3188 113600 3194
rect 113548 3130 113600 3136
rect 114284 3188 114336 3194
rect 114284 3130 114336 3136
rect 113088 2984 113140 2990
rect 113088 2926 113140 2932
rect 113560 480 113588 3130
rect 114388 3058 114416 317426
rect 114480 3369 114508 320076
rect 114940 317490 114968 320076
rect 115414 320062 115796 320090
rect 114928 317484 114980 317490
rect 114928 317426 114980 317432
rect 114466 3360 114522 3369
rect 114466 3295 114522 3304
rect 114744 3256 114796 3262
rect 114744 3198 114796 3204
rect 114376 3052 114428 3058
rect 114376 2994 114428 3000
rect 114756 480 114784 3198
rect 115768 2961 115796 320062
rect 115860 318782 115888 320076
rect 115848 318776 115900 318782
rect 115848 318718 115900 318724
rect 116228 317490 116256 320076
rect 116702 320062 117084 320090
rect 115848 317484 115900 317490
rect 115848 317426 115900 317432
rect 116216 317484 116268 317490
rect 116216 317426 116268 317432
rect 116952 317484 117004 317490
rect 116952 317426 117004 317432
rect 115860 3262 115888 317426
rect 116964 315874 116992 317426
rect 117056 316010 117084 320062
rect 117148 318714 117176 320076
rect 117622 320062 117912 320090
rect 118082 320062 118464 320090
rect 117136 318708 117188 318714
rect 117136 318650 117188 318656
rect 117056 315982 117268 316010
rect 116964 315846 117176 315874
rect 117148 6882 117176 315846
rect 116964 6854 117176 6882
rect 116964 3330 116992 6854
rect 117240 4146 117268 315982
rect 117884 315926 117912 320062
rect 118436 316010 118464 320062
rect 118528 318646 118556 320076
rect 118516 318640 118568 318646
rect 118516 318582 118568 318588
rect 118988 317490 119016 320076
rect 119448 317694 119476 320076
rect 119830 320062 120028 320090
rect 119436 317688 119488 317694
rect 119436 317630 119488 317636
rect 118976 317484 119028 317490
rect 118976 317426 119028 317432
rect 119896 317484 119948 317490
rect 119896 317426 119948 317432
rect 118436 315982 118648 316010
rect 117872 315920 117924 315926
rect 117872 315862 117924 315868
rect 118516 315920 118568 315926
rect 118516 315862 118568 315868
rect 117136 4140 117188 4146
rect 117136 4082 117188 4088
rect 117228 4140 117280 4146
rect 117228 4082 117280 4088
rect 115940 3324 115992 3330
rect 115940 3266 115992 3272
rect 116952 3324 117004 3330
rect 116952 3266 117004 3272
rect 115848 3256 115900 3262
rect 115848 3198 115900 3204
rect 115754 2952 115810 2961
rect 115754 2887 115810 2896
rect 115952 480 115980 3266
rect 117148 480 117176 4082
rect 118528 4078 118556 315862
rect 118240 4072 118292 4078
rect 118240 4014 118292 4020
rect 118516 4072 118568 4078
rect 118516 4014 118568 4020
rect 118252 480 118280 4014
rect 118620 3097 118648 315982
rect 119908 4214 119936 317426
rect 119896 4208 119948 4214
rect 119896 4150 119948 4156
rect 120000 3505 120028 320062
rect 120276 317490 120304 320076
rect 120736 318102 120764 320076
rect 121210 320062 121408 320090
rect 120724 318096 120776 318102
rect 120724 318038 120776 318044
rect 120264 317484 120316 317490
rect 120264 317426 120316 317432
rect 121276 317484 121328 317490
rect 121276 317426 121328 317432
rect 121288 4010 121316 317426
rect 120632 4004 120684 4010
rect 120632 3946 120684 3952
rect 121276 4004 121328 4010
rect 121276 3946 121328 3952
rect 119986 3496 120042 3505
rect 119986 3431 120042 3440
rect 119436 3392 119488 3398
rect 119436 3334 119488 3340
rect 118606 3088 118662 3097
rect 118606 3023 118662 3032
rect 119448 480 119476 3334
rect 120644 480 120672 3946
rect 121380 3641 121408 320062
rect 121656 317490 121684 320076
rect 122116 318170 122144 320076
rect 122590 320062 122788 320090
rect 122104 318164 122156 318170
rect 122104 318106 122156 318112
rect 121644 317484 121696 317490
rect 121644 317426 121696 317432
rect 122656 317484 122708 317490
rect 122656 317426 122708 317432
rect 122668 6050 122696 317426
rect 122656 6044 122708 6050
rect 122656 5986 122708 5992
rect 122760 3874 122788 320062
rect 123036 317490 123064 320076
rect 123496 317626 123524 320076
rect 123878 320062 124076 320090
rect 123484 317620 123536 317626
rect 123484 317562 123536 317568
rect 123024 317484 123076 317490
rect 123024 317426 123076 317432
rect 123944 317484 123996 317490
rect 123944 317426 123996 317432
rect 123956 6118 123984 317426
rect 123944 6112 123996 6118
rect 123944 6054 123996 6060
rect 121828 3868 121880 3874
rect 121828 3810 121880 3816
rect 122748 3868 122800 3874
rect 122748 3810 122800 3816
rect 121366 3632 121422 3641
rect 121366 3567 121422 3576
rect 121840 480 121868 3810
rect 123024 3732 123076 3738
rect 123024 3674 123076 3680
rect 123036 480 123064 3674
rect 124048 3233 124076 320062
rect 124128 317620 124180 317626
rect 124128 317562 124180 317568
rect 124140 3738 124168 317562
rect 124324 317490 124352 320076
rect 124784 318510 124812 320076
rect 125258 320062 125548 320090
rect 124772 318504 124824 318510
rect 124772 318446 124824 318452
rect 124312 317484 124364 317490
rect 124312 317426 124364 317432
rect 125416 317484 125468 317490
rect 125416 317426 125468 317432
rect 124496 307896 124548 307902
rect 124416 307844 124496 307850
rect 124416 307838 124548 307844
rect 124416 307822 124536 307838
rect 124416 307766 124444 307822
rect 124404 307760 124456 307766
rect 124404 307702 124456 307708
rect 124220 298240 124272 298246
rect 124220 298182 124272 298188
rect 124232 298110 124260 298182
rect 124220 298104 124272 298110
rect 124220 298046 124272 298052
rect 124404 292460 124456 292466
rect 124404 292402 124456 292408
rect 124416 283014 124444 292402
rect 124404 283008 124456 283014
rect 124404 282950 124456 282956
rect 124404 282872 124456 282878
rect 124404 282814 124456 282820
rect 124416 280158 124444 282814
rect 124404 280152 124456 280158
rect 124404 280094 124456 280100
rect 124404 273964 124456 273970
rect 124404 273906 124456 273912
rect 124416 269090 124444 273906
rect 124324 269062 124444 269090
rect 124324 263634 124352 269062
rect 124312 263628 124364 263634
rect 124312 263570 124364 263576
rect 124312 259480 124364 259486
rect 124312 259422 124364 259428
rect 124324 253978 124352 259422
rect 124312 253972 124364 253978
rect 124312 253914 124364 253920
rect 124404 253836 124456 253842
rect 124404 253778 124456 253784
rect 124416 244390 124444 253778
rect 124404 244384 124456 244390
rect 124404 244326 124456 244332
rect 124312 244248 124364 244254
rect 124312 244190 124364 244196
rect 124324 234666 124352 244190
rect 124312 234660 124364 234666
rect 124312 234602 124364 234608
rect 124404 234524 124456 234530
rect 124404 234466 124456 234472
rect 124416 231826 124444 234466
rect 124324 231798 124444 231826
rect 124324 225010 124352 231798
rect 124312 225004 124364 225010
rect 124312 224946 124364 224952
rect 124312 222216 124364 222222
rect 124312 222158 124364 222164
rect 124324 215354 124352 222158
rect 124312 215348 124364 215354
rect 124312 215290 124364 215296
rect 124404 215212 124456 215218
rect 124404 215154 124456 215160
rect 124416 212514 124444 215154
rect 124324 212486 124444 212514
rect 124324 205698 124352 212486
rect 124312 205692 124364 205698
rect 124312 205634 124364 205640
rect 124312 202904 124364 202910
rect 124312 202846 124364 202852
rect 124324 196042 124352 202846
rect 124312 196036 124364 196042
rect 124312 195978 124364 195984
rect 124404 195900 124456 195906
rect 124404 195842 124456 195848
rect 124416 193202 124444 195842
rect 124324 193174 124444 193202
rect 124324 186386 124352 193174
rect 124312 186380 124364 186386
rect 124312 186322 124364 186328
rect 124312 183592 124364 183598
rect 124312 183534 124364 183540
rect 124324 176730 124352 183534
rect 124312 176724 124364 176730
rect 124312 176666 124364 176672
rect 124404 176588 124456 176594
rect 124404 176530 124456 176536
rect 124416 173890 124444 176530
rect 124324 173862 124444 173890
rect 124324 167074 124352 173862
rect 124312 167068 124364 167074
rect 124312 167010 124364 167016
rect 124312 164280 124364 164286
rect 124312 164222 124364 164228
rect 124324 157418 124352 164222
rect 124312 157412 124364 157418
rect 124312 157354 124364 157360
rect 124404 157276 124456 157282
rect 124404 157218 124456 157224
rect 124416 154562 124444 157218
rect 124404 154556 124456 154562
rect 124404 154498 124456 154504
rect 124588 154556 124640 154562
rect 124588 154498 124640 154504
rect 124600 144945 124628 154498
rect 124310 144936 124366 144945
rect 124310 144871 124366 144880
rect 124586 144936 124642 144945
rect 124586 144871 124642 144880
rect 124324 138038 124352 144871
rect 124312 138032 124364 138038
rect 124312 137974 124364 137980
rect 124404 137964 124456 137970
rect 124404 137906 124456 137912
rect 124416 135250 124444 137906
rect 124404 135244 124456 135250
rect 124404 135186 124456 135192
rect 124588 135244 124640 135250
rect 124588 135186 124640 135192
rect 124600 125633 124628 135186
rect 124310 125624 124366 125633
rect 124310 125559 124366 125568
rect 124586 125624 124642 125633
rect 124586 125559 124642 125568
rect 124324 118726 124352 125559
rect 124312 118720 124364 118726
rect 124312 118662 124364 118668
rect 124404 118652 124456 118658
rect 124404 118594 124456 118600
rect 124416 115938 124444 118594
rect 124404 115932 124456 115938
rect 124404 115874 124456 115880
rect 124588 115932 124640 115938
rect 124588 115874 124640 115880
rect 124600 106321 124628 115874
rect 124310 106312 124366 106321
rect 124310 106247 124366 106256
rect 124586 106312 124642 106321
rect 124586 106247 124642 106256
rect 124324 99414 124352 106247
rect 124312 99408 124364 99414
rect 124312 99350 124364 99356
rect 124404 99340 124456 99346
rect 124404 99282 124456 99288
rect 124416 96626 124444 99282
rect 124404 96620 124456 96626
rect 124404 96562 124456 96568
rect 124588 96620 124640 96626
rect 124588 96562 124640 96568
rect 124600 87009 124628 96562
rect 124310 87000 124366 87009
rect 124310 86935 124366 86944
rect 124586 87000 124642 87009
rect 124586 86935 124642 86944
rect 124324 80102 124352 86935
rect 124312 80096 124364 80102
rect 124312 80038 124364 80044
rect 124404 79960 124456 79966
rect 124404 79902 124456 79908
rect 124416 66298 124444 79902
rect 124404 66292 124456 66298
rect 124404 66234 124456 66240
rect 124588 66292 124640 66298
rect 124588 66234 124640 66240
rect 124600 60654 124628 66234
rect 124404 60648 124456 60654
rect 124404 60590 124456 60596
rect 124588 60648 124640 60654
rect 124588 60590 124640 60596
rect 124416 56574 124444 60590
rect 124404 56568 124456 56574
rect 124404 56510 124456 56516
rect 124496 46980 124548 46986
rect 124496 46922 124548 46928
rect 124508 42129 124536 46922
rect 124494 42120 124550 42129
rect 124494 42055 124550 42064
rect 124402 32464 124458 32473
rect 124402 32399 124458 32408
rect 124416 27674 124444 32399
rect 124404 27668 124456 27674
rect 124404 27610 124456 27616
rect 124588 27668 124640 27674
rect 124588 27610 124640 27616
rect 124600 18018 124628 27610
rect 124404 18012 124456 18018
rect 124404 17954 124456 17960
rect 124588 18012 124640 18018
rect 124588 17954 124640 17960
rect 124416 13122 124444 17954
rect 124404 13116 124456 13122
rect 124404 13058 124456 13064
rect 125324 13116 125376 13122
rect 125324 13058 125376 13064
rect 125336 6746 125364 13058
rect 125428 6866 125456 317426
rect 125416 6860 125468 6866
rect 125416 6802 125468 6808
rect 125336 6718 125456 6746
rect 124220 3936 124272 3942
rect 124220 3878 124272 3884
rect 124128 3732 124180 3738
rect 124128 3674 124180 3680
rect 124034 3224 124090 3233
rect 124034 3159 124090 3168
rect 124232 480 124260 3878
rect 125428 480 125456 6718
rect 125520 3942 125548 320062
rect 125704 317490 125732 320076
rect 126164 318374 126192 320076
rect 126152 318368 126204 318374
rect 126152 318310 126204 318316
rect 125692 317484 125744 317490
rect 125692 317426 125744 317432
rect 126624 317422 126652 320076
rect 127084 317898 127112 320076
rect 127452 318306 127480 320076
rect 127440 318300 127492 318306
rect 127440 318242 127492 318248
rect 127624 318028 127676 318034
rect 127624 317970 127676 317976
rect 127072 317892 127124 317898
rect 127072 317834 127124 317840
rect 126888 317484 126940 317490
rect 126888 317426 126940 317432
rect 126612 317416 126664 317422
rect 126612 317358 126664 317364
rect 126900 6798 126928 317426
rect 126888 6792 126940 6798
rect 126888 6734 126940 6740
rect 125508 3936 125560 3942
rect 125508 3878 125560 3884
rect 127636 3738 127664 317970
rect 127912 317830 127940 320076
rect 128268 317892 128320 317898
rect 128268 317834 128320 317840
rect 127900 317824 127952 317830
rect 127900 317766 127952 317772
rect 128280 6730 128308 317834
rect 128372 315450 128400 320076
rect 128636 318436 128688 318442
rect 128636 318378 128688 318384
rect 128360 315444 128412 315450
rect 128360 315386 128412 315392
rect 128268 6724 128320 6730
rect 128268 6666 128320 6672
rect 127624 3732 127676 3738
rect 127624 3674 127676 3680
rect 127808 3392 127860 3398
rect 127808 3334 127860 3340
rect 126612 2848 126664 2854
rect 126612 2790 126664 2796
rect 126624 480 126652 2790
rect 127820 480 127848 3334
rect 128648 610 128676 318378
rect 128832 317490 128860 320076
rect 129292 317898 129320 320076
rect 129280 317892 129332 317898
rect 129280 317834 129332 317840
rect 129752 317490 129780 320076
rect 130212 318442 130240 320076
rect 130200 318436 130252 318442
rect 130200 318378 130252 318384
rect 130672 317966 130700 320076
rect 130948 320062 131054 320090
rect 130660 317960 130712 317966
rect 130660 317902 130712 317908
rect 130384 317552 130436 317558
rect 130384 317494 130436 317500
rect 128820 317484 128872 317490
rect 128820 317426 128872 317432
rect 129648 317484 129700 317490
rect 129648 317426 129700 317432
rect 129740 317484 129792 317490
rect 129740 317426 129792 317432
rect 129556 315444 129608 315450
rect 129556 315386 129608 315392
rect 129568 6662 129596 315386
rect 129556 6656 129608 6662
rect 129556 6598 129608 6604
rect 129660 2854 129688 317426
rect 130396 3670 130424 317494
rect 130948 6526 130976 320062
rect 131500 317490 131528 320076
rect 131960 317694 131988 320076
rect 132328 320062 132434 320090
rect 131948 317688 132000 317694
rect 131948 317630 132000 317636
rect 131028 317484 131080 317490
rect 131028 317426 131080 317432
rect 131488 317484 131540 317490
rect 131488 317426 131540 317432
rect 131040 6594 131068 317426
rect 131028 6588 131080 6594
rect 131028 6530 131080 6536
rect 130936 6520 130988 6526
rect 130936 6462 130988 6468
rect 132328 6458 132356 320062
rect 132880 317490 132908 320076
rect 133144 318572 133196 318578
rect 133144 318514 133196 318520
rect 132408 317484 132460 317490
rect 132408 317426 132460 317432
rect 132868 317484 132920 317490
rect 132868 317426 132920 317432
rect 132316 6452 132368 6458
rect 132316 6394 132368 6400
rect 131396 3800 131448 3806
rect 131396 3742 131448 3748
rect 130384 3664 130436 3670
rect 130384 3606 130436 3612
rect 130200 3120 130252 3126
rect 130200 3062 130252 3068
rect 129556 2848 129608 2854
rect 129554 2816 129556 2825
rect 129648 2848 129700 2854
rect 129608 2816 129610 2825
rect 129648 2790 129700 2796
rect 129554 2751 129610 2760
rect 128636 604 128688 610
rect 128636 546 128688 552
rect 129004 604 129056 610
rect 129004 546 129056 552
rect 129016 480 129044 546
rect 130212 480 130240 3062
rect 131408 480 131436 3742
rect 132420 3670 132448 317426
rect 133156 3670 133184 318514
rect 133340 317558 133368 320076
rect 133708 320062 133814 320090
rect 133328 317552 133380 317558
rect 133328 317494 133380 317500
rect 133708 6390 133736 320062
rect 134260 318578 134288 320076
rect 134248 318572 134300 318578
rect 134248 318514 134300 318520
rect 134720 317966 134748 320076
rect 135102 320062 135208 320090
rect 135562 320062 135944 320090
rect 134616 317960 134668 317966
rect 134614 317928 134616 317937
rect 134708 317960 134760 317966
rect 134668 317928 134670 317937
rect 134708 317902 134760 317908
rect 134614 317863 134670 317872
rect 133788 317484 133840 317490
rect 133788 317426 133840 317432
rect 133696 6384 133748 6390
rect 133696 6326 133748 6332
rect 133800 6202 133828 317426
rect 135180 311982 135208 320062
rect 135916 317422 135944 320062
rect 136008 319054 136036 320076
rect 135996 319048 136048 319054
rect 135996 318990 136048 318996
rect 136468 318209 136496 320076
rect 136652 320062 136942 320090
rect 137402 320062 137600 320090
rect 136548 319048 136600 319054
rect 136548 318990 136600 318996
rect 136454 318200 136510 318209
rect 136454 318135 136510 318144
rect 135904 317416 135956 317422
rect 135904 317358 135956 317364
rect 135168 311976 135220 311982
rect 135168 311918 135220 311924
rect 135076 309188 135128 309194
rect 135076 309130 135128 309136
rect 135088 309074 135116 309130
rect 134996 309046 135116 309074
rect 134996 302258 135024 309046
rect 134984 302252 135036 302258
rect 134984 302194 135036 302200
rect 134984 299532 135036 299538
rect 134984 299474 135036 299480
rect 134996 292618 135024 299474
rect 134996 292590 135208 292618
rect 135180 289814 135208 292590
rect 135168 289808 135220 289814
rect 135168 289750 135220 289756
rect 134892 280220 134944 280226
rect 134892 280162 134944 280168
rect 134904 280106 134932 280162
rect 134982 280120 135038 280129
rect 134904 280078 134982 280106
rect 134982 280055 135038 280064
rect 134982 270600 135038 270609
rect 134982 270535 135038 270544
rect 134996 270502 135024 270535
rect 134984 270496 135036 270502
rect 134984 270438 135036 270444
rect 134892 260908 134944 260914
rect 134892 260850 134944 260856
rect 134904 260794 134932 260850
rect 134982 260808 135038 260817
rect 134904 260766 134982 260794
rect 134982 260743 135038 260752
rect 134982 251288 135038 251297
rect 134982 251223 135038 251232
rect 134996 251190 135024 251223
rect 134984 251184 135036 251190
rect 134984 251126 135036 251132
rect 134892 241528 134944 241534
rect 134892 241470 134944 241476
rect 134904 234666 134932 241470
rect 134892 234660 134944 234666
rect 134892 234602 134944 234608
rect 134984 234524 135036 234530
rect 134984 234466 135036 234472
rect 134996 231826 135024 234466
rect 134904 231798 135024 231826
rect 134904 225010 134932 231798
rect 134892 225004 134944 225010
rect 134892 224946 134944 224952
rect 134892 222216 134944 222222
rect 134892 222158 134944 222164
rect 134904 215354 134932 222158
rect 134892 215348 134944 215354
rect 134892 215290 134944 215296
rect 134984 215212 135036 215218
rect 134984 215154 135036 215160
rect 134996 212514 135024 215154
rect 134904 212486 135024 212514
rect 134904 205698 134932 212486
rect 134892 205692 134944 205698
rect 134892 205634 134944 205640
rect 134892 202904 134944 202910
rect 134892 202846 134944 202852
rect 134904 196042 134932 202846
rect 134892 196036 134944 196042
rect 134892 195978 134944 195984
rect 134984 195900 135036 195906
rect 134984 195842 135036 195848
rect 134996 193225 135024 195842
rect 134798 193216 134854 193225
rect 134798 193151 134854 193160
rect 134982 193216 135038 193225
rect 134982 193151 135038 193160
rect 134812 183598 134840 193151
rect 134800 183592 134852 183598
rect 134800 183534 134852 183540
rect 135076 183592 135128 183598
rect 135076 183534 135128 183540
rect 135088 176798 135116 183534
rect 135076 176792 135128 176798
rect 135076 176734 135128 176740
rect 134984 176588 135036 176594
rect 134984 176530 135036 176536
rect 134996 173913 135024 176530
rect 134798 173904 134854 173913
rect 134798 173839 134854 173848
rect 134982 173904 135038 173913
rect 134982 173839 135038 173848
rect 134812 167006 134840 173839
rect 134800 167000 134852 167006
rect 134800 166942 134852 166948
rect 134984 167000 135036 167006
rect 134984 166942 135036 166948
rect 134996 164234 135024 166942
rect 134996 164206 135116 164234
rect 135088 157486 135116 164206
rect 135076 157480 135128 157486
rect 135076 157422 135128 157428
rect 135076 154624 135128 154630
rect 135076 154566 135128 154572
rect 135088 147694 135116 154566
rect 135076 147688 135128 147694
rect 135076 147630 135128 147636
rect 135076 144968 135128 144974
rect 135076 144910 135128 144916
rect 135088 138106 135116 144910
rect 135076 138100 135128 138106
rect 135076 138042 135128 138048
rect 134984 137964 135036 137970
rect 134984 137906 135036 137912
rect 134996 128382 135024 137906
rect 134984 128376 135036 128382
rect 134984 128318 135036 128324
rect 135076 128308 135128 128314
rect 135076 128250 135128 128256
rect 135088 124166 135116 128250
rect 135076 124160 135128 124166
rect 135076 124102 135128 124108
rect 134984 114572 135036 114578
rect 134984 114514 135036 114520
rect 134996 109070 135024 114514
rect 134984 109064 135036 109070
rect 134984 109006 135036 109012
rect 135076 108996 135128 109002
rect 135076 108938 135128 108944
rect 135088 104854 135116 108938
rect 135076 104848 135128 104854
rect 135076 104790 135128 104796
rect 134984 89684 135036 89690
rect 134984 89626 135036 89632
rect 134996 86986 135024 89626
rect 134996 86958 135116 86986
rect 135088 82142 135116 86958
rect 134708 82136 134760 82142
rect 134708 82078 134760 82084
rect 135076 82136 135128 82142
rect 135076 82078 135128 82084
rect 134720 77353 134748 82078
rect 134706 77344 134762 77353
rect 134706 77279 134762 77288
rect 134890 77344 134946 77353
rect 134946 77302 135024 77330
rect 134890 77279 134946 77288
rect 134996 70514 135024 77302
rect 134984 70508 135036 70514
rect 134984 70450 135036 70456
rect 134892 70372 134944 70378
rect 134892 70314 134944 70320
rect 134904 67833 134932 70314
rect 134890 67824 134946 67833
rect 134890 67759 134946 67768
rect 134890 67688 134946 67697
rect 134890 67623 134946 67632
rect 134904 66230 134932 67623
rect 134892 66224 134944 66230
rect 134892 66166 134944 66172
rect 135076 66224 135128 66230
rect 135076 66166 135128 66172
rect 135088 61441 135116 66166
rect 135074 61432 135130 61441
rect 135074 61367 135130 61376
rect 134982 48376 135038 48385
rect 134904 48334 134982 48362
rect 134904 46918 134932 48334
rect 134982 48311 135038 48320
rect 134892 46912 134944 46918
rect 134892 46854 134944 46860
rect 135076 46912 135128 46918
rect 135076 46854 135128 46860
rect 135088 42129 135116 46854
rect 135074 42120 135130 42129
rect 135074 42055 135130 42064
rect 134982 29064 135038 29073
rect 134904 29022 134982 29050
rect 134904 27606 134932 29022
rect 134982 28999 135038 29008
rect 134892 27600 134944 27606
rect 134892 27542 134944 27548
rect 134984 18012 135036 18018
rect 134984 17954 135036 17960
rect 134996 12510 135024 17954
rect 134984 12504 135036 12510
rect 134984 12446 135036 12452
rect 134892 12436 134944 12442
rect 134892 12378 134944 12384
rect 134904 6322 134932 12378
rect 134892 6316 134944 6322
rect 134892 6258 134944 6264
rect 133708 6174 133828 6202
rect 132408 3664 132460 3670
rect 132408 3606 132460 3612
rect 133144 3664 133196 3670
rect 133144 3606 133196 3612
rect 132592 3596 132644 3602
rect 132592 3538 132644 3544
rect 132604 480 132632 3538
rect 133708 3466 133736 6174
rect 136560 4214 136588 318990
rect 136652 307086 136680 320062
rect 137572 316010 137600 320062
rect 137848 316146 137876 320076
rect 138112 318776 138164 318782
rect 138112 318718 138164 318724
rect 137926 317928 137982 317937
rect 137926 317863 137982 317872
rect 137940 317626 137968 317863
rect 138124 317778 138152 318718
rect 138032 317750 138152 317778
rect 138032 317694 138060 317750
rect 138020 317688 138072 317694
rect 138020 317630 138072 317636
rect 137928 317620 137980 317626
rect 137928 317562 137980 317568
rect 138308 317558 138336 320076
rect 138296 317552 138348 317558
rect 138296 317494 138348 317500
rect 138676 317490 138704 320076
rect 138664 317484 138716 317490
rect 138664 317426 138716 317432
rect 137848 316118 137968 316146
rect 137572 315982 137876 316010
rect 137744 311908 137796 311914
rect 137744 311850 137796 311856
rect 136640 307080 136692 307086
rect 136640 307022 136692 307028
rect 137756 8226 137784 311850
rect 137744 8220 137796 8226
rect 137744 8162 137796 8168
rect 137848 4282 137876 315982
rect 137940 311914 137968 316118
rect 137928 311908 137980 311914
rect 137928 311850 137980 311856
rect 137928 307080 137980 307086
rect 137928 307022 137980 307028
rect 137836 4276 137888 4282
rect 137836 4218 137888 4224
rect 136548 4208 136600 4214
rect 136548 4150 136600 4156
rect 133788 3732 133840 3738
rect 133788 3674 133840 3680
rect 133696 3460 133748 3466
rect 133696 3402 133748 3408
rect 133800 480 133828 3674
rect 137284 3664 137336 3670
rect 137284 3606 137336 3612
rect 136088 3528 136140 3534
rect 136088 3470 136140 3476
rect 134892 2916 134944 2922
rect 134892 2858 134944 2864
rect 133972 2848 134024 2854
rect 133970 2816 133972 2825
rect 134024 2816 134026 2825
rect 133970 2751 134026 2760
rect 134904 480 134932 2858
rect 136100 480 136128 3470
rect 137296 480 137324 3606
rect 137940 3534 137968 307022
rect 139136 8158 139164 320076
rect 139412 320062 139610 320090
rect 139308 317552 139360 317558
rect 139308 317494 139360 317500
rect 139216 317484 139268 317490
rect 139216 317426 139268 317432
rect 139124 8152 139176 8158
rect 139124 8094 139176 8100
rect 139228 4350 139256 317426
rect 139216 4344 139268 4350
rect 139216 4286 139268 4292
rect 137928 3528 137980 3534
rect 137928 3470 137980 3476
rect 138480 3120 138532 3126
rect 138480 3062 138532 3068
rect 138492 480 138520 3062
rect 139320 2922 139348 317494
rect 139412 307086 139440 320062
rect 140056 317490 140084 320076
rect 140044 317484 140096 317490
rect 140044 317426 140096 317432
rect 139400 307080 139452 307086
rect 139400 307022 139452 307028
rect 140516 8090 140544 320076
rect 140884 320062 140990 320090
rect 140780 317688 140832 317694
rect 140780 317630 140832 317636
rect 140596 317484 140648 317490
rect 140596 317426 140648 317432
rect 140504 8084 140556 8090
rect 140504 8026 140556 8032
rect 140608 4418 140636 317426
rect 140792 311846 140820 317630
rect 140780 311840 140832 311846
rect 140780 311782 140832 311788
rect 140884 307086 140912 320062
rect 141436 317490 141464 320076
rect 141424 317484 141476 317490
rect 141424 317426 141476 317432
rect 140964 311840 141016 311846
rect 140964 311782 141016 311788
rect 140688 307080 140740 307086
rect 140688 307022 140740 307028
rect 140872 307080 140924 307086
rect 140872 307022 140924 307028
rect 140596 4412 140648 4418
rect 140596 4354 140648 4360
rect 140700 4049 140728 307022
rect 140976 296750 141004 311782
rect 140780 296744 140832 296750
rect 140780 296686 140832 296692
rect 140964 296744 141016 296750
rect 140964 296686 141016 296692
rect 140792 292482 140820 296686
rect 140792 292454 140912 292482
rect 140884 282962 140912 292454
rect 140884 282934 141004 282962
rect 140976 263634 141004 282934
rect 140780 263628 140832 263634
rect 140780 263570 140832 263576
rect 140964 263628 141016 263634
rect 140964 263570 141016 263576
rect 140792 263514 140820 263570
rect 140792 263486 140912 263514
rect 140884 253994 140912 263486
rect 140884 253966 141004 253994
rect 140976 244322 141004 253966
rect 140780 244316 140832 244322
rect 140780 244258 140832 244264
rect 140964 244316 141016 244322
rect 140964 244258 141016 244264
rect 140792 244202 140820 244258
rect 140792 244174 140912 244202
rect 140884 234682 140912 244174
rect 140884 234654 141004 234682
rect 140976 225010 141004 234654
rect 140780 225004 140832 225010
rect 140780 224946 140832 224952
rect 140964 225004 141016 225010
rect 140964 224946 141016 224952
rect 140792 224890 140820 224946
rect 140792 224862 140912 224890
rect 140884 215370 140912 224862
rect 140884 215342 141004 215370
rect 140976 205698 141004 215342
rect 140780 205692 140832 205698
rect 140780 205634 140832 205640
rect 140964 205692 141016 205698
rect 140964 205634 141016 205640
rect 140792 205578 140820 205634
rect 140792 205550 140912 205578
rect 140884 196058 140912 205550
rect 140884 196030 141004 196058
rect 140976 186386 141004 196030
rect 140780 186380 140832 186386
rect 140780 186322 140832 186328
rect 140964 186380 141016 186386
rect 140964 186322 141016 186328
rect 140792 186266 140820 186322
rect 140792 186238 140912 186266
rect 140884 183569 140912 186238
rect 140870 183560 140926 183569
rect 140870 183495 140926 183504
rect 141146 183560 141202 183569
rect 141146 183495 141202 183504
rect 141160 173942 141188 183495
rect 140964 173936 141016 173942
rect 140964 173878 141016 173884
rect 141148 173936 141200 173942
rect 141148 173878 141200 173884
rect 140976 167074 141004 173878
rect 140780 167068 140832 167074
rect 140780 167010 140832 167016
rect 140964 167068 141016 167074
rect 140964 167010 141016 167016
rect 140792 166954 140820 167010
rect 140792 166926 140912 166954
rect 140884 164218 140912 166926
rect 140872 164212 140924 164218
rect 140872 164154 140924 164160
rect 140872 157344 140924 157350
rect 140872 157286 140924 157292
rect 140884 154578 140912 157286
rect 140884 154550 141004 154578
rect 140976 147694 141004 154550
rect 140780 147688 140832 147694
rect 140964 147688 141016 147694
rect 140832 147636 140912 147642
rect 140780 147630 140912 147636
rect 140964 147630 141016 147636
rect 140792 147614 140912 147630
rect 140884 144906 140912 147614
rect 140872 144900 140924 144906
rect 140872 144842 140924 144848
rect 140872 137964 140924 137970
rect 140872 137906 140924 137912
rect 140884 135266 140912 137906
rect 140884 135238 141004 135266
rect 140976 128382 141004 135238
rect 140780 128376 140832 128382
rect 140964 128376 141016 128382
rect 140832 128324 140912 128330
rect 140780 128318 140912 128324
rect 140964 128318 141016 128324
rect 140792 128302 140912 128318
rect 140884 125594 140912 128302
rect 140872 125588 140924 125594
rect 140872 125530 140924 125536
rect 140872 118652 140924 118658
rect 140872 118594 140924 118600
rect 140884 115954 140912 118594
rect 140884 115926 141004 115954
rect 140976 109070 141004 115926
rect 140780 109064 140832 109070
rect 140964 109064 141016 109070
rect 140832 109012 140912 109018
rect 140780 109006 140912 109012
rect 140964 109006 141016 109012
rect 140792 108990 140912 109006
rect 140884 106282 140912 108990
rect 140872 106276 140924 106282
rect 140872 106218 140924 106224
rect 140872 99340 140924 99346
rect 140872 99282 140924 99288
rect 140884 96642 140912 99282
rect 140884 96614 141004 96642
rect 140976 89758 141004 96614
rect 140780 89752 140832 89758
rect 140964 89752 141016 89758
rect 140832 89700 140912 89706
rect 140780 89694 140912 89700
rect 140964 89694 141016 89700
rect 140792 89678 140912 89694
rect 140884 86970 140912 89678
rect 140872 86964 140924 86970
rect 140872 86906 140924 86912
rect 140964 77308 141016 77314
rect 140964 77250 141016 77256
rect 140976 77178 141004 77250
rect 140964 77172 141016 77178
rect 140964 77114 141016 77120
rect 140872 67652 140924 67658
rect 140872 67594 140924 67600
rect 140884 60738 140912 67594
rect 140884 60710 141004 60738
rect 140976 57934 141004 60710
rect 140964 57928 141016 57934
rect 140964 57870 141016 57876
rect 140872 51060 140924 51066
rect 140872 51002 140924 51008
rect 140884 41426 140912 51002
rect 140884 41398 141004 41426
rect 140976 38622 141004 41398
rect 140964 38616 141016 38622
rect 140964 38558 141016 38564
rect 140872 31748 140924 31754
rect 140872 31690 140924 31696
rect 140884 22114 140912 31690
rect 140884 22086 141004 22114
rect 140976 12458 141004 22086
rect 140792 12430 141004 12458
rect 140792 9654 140820 12430
rect 140780 9648 140832 9654
rect 140780 9590 140832 9596
rect 141896 8022 141924 320076
rect 142264 317558 142292 320076
rect 142252 317552 142304 317558
rect 142252 317494 142304 317500
rect 142724 317490 142752 320076
rect 143198 320062 143304 320090
rect 141976 317484 142028 317490
rect 141976 317426 142028 317432
rect 142712 317484 142764 317490
rect 142712 317426 142764 317432
rect 141884 8016 141936 8022
rect 141884 7958 141936 7964
rect 141988 4486 142016 317426
rect 142068 307080 142120 307086
rect 142068 307022 142120 307028
rect 141976 4480 142028 4486
rect 141976 4422 142028 4428
rect 140686 4040 140742 4049
rect 140686 3975 140742 3984
rect 142080 3913 142108 307022
rect 143276 7954 143304 320062
rect 143448 317552 143500 317558
rect 143448 317494 143500 317500
rect 143356 317484 143408 317490
rect 143356 317426 143408 317432
rect 143264 7948 143316 7954
rect 143264 7890 143316 7896
rect 143368 4554 143396 317426
rect 143356 4548 143408 4554
rect 143356 4490 143408 4496
rect 142066 3904 142122 3913
rect 142066 3839 142122 3848
rect 143460 3777 143488 317494
rect 143644 307086 143672 320076
rect 144104 317490 144132 320076
rect 144578 320062 144684 320090
rect 144092 317484 144144 317490
rect 144092 317426 144144 317432
rect 143632 307080 143684 307086
rect 143632 307022 143684 307028
rect 144656 7886 144684 320062
rect 145024 318646 145052 320076
rect 145012 318640 145064 318646
rect 145012 318582 145064 318588
rect 145484 317490 145512 320076
rect 145958 320062 146156 320090
rect 145656 318844 145708 318850
rect 145656 318786 145708 318792
rect 145564 317688 145616 317694
rect 145564 317630 145616 317636
rect 144736 317484 144788 317490
rect 144736 317426 144788 317432
rect 145472 317484 145524 317490
rect 145472 317426 145524 317432
rect 144644 7880 144696 7886
rect 144644 7822 144696 7828
rect 144748 4622 144776 317426
rect 144828 307080 144880 307086
rect 144828 307022 144880 307028
rect 144736 4616 144788 4622
rect 144736 4558 144788 4564
rect 143446 3768 143502 3777
rect 143446 3703 143502 3712
rect 144840 3369 144868 307022
rect 144458 3360 144514 3369
rect 144458 3295 144514 3304
rect 144826 3360 144882 3369
rect 144826 3295 144882 3304
rect 143264 3188 143316 3194
rect 143264 3130 143316 3136
rect 142068 3052 142120 3058
rect 142068 2994 142120 3000
rect 139676 2984 139728 2990
rect 139676 2926 139728 2932
rect 139308 2916 139360 2922
rect 139308 2858 139360 2864
rect 139688 480 139716 2926
rect 140872 604 140924 610
rect 140872 546 140924 552
rect 140884 480 140912 546
rect 142080 480 142108 2994
rect 143276 480 143304 3130
rect 144472 480 144500 3295
rect 145576 2922 145604 317630
rect 145668 7834 145696 318786
rect 145668 7806 145880 7834
rect 145852 3330 145880 7806
rect 146128 7750 146156 320062
rect 146312 317490 146340 320076
rect 146772 317966 146800 320076
rect 147246 320062 147444 320090
rect 146760 317960 146812 317966
rect 146760 317902 146812 317908
rect 146208 317484 146260 317490
rect 146208 317426 146260 317432
rect 146300 317484 146352 317490
rect 146300 317426 146352 317432
rect 146116 7744 146168 7750
rect 146116 7686 146168 7692
rect 146220 4690 146248 317426
rect 147416 7614 147444 320062
rect 147692 317966 147720 320076
rect 147588 317960 147640 317966
rect 147588 317902 147640 317908
rect 147680 317960 147732 317966
rect 147680 317902 147732 317908
rect 147496 317484 147548 317490
rect 147496 317426 147548 317432
rect 147508 7818 147536 317426
rect 147496 7812 147548 7818
rect 147496 7754 147548 7760
rect 147404 7608 147456 7614
rect 147404 7550 147456 7556
rect 147600 4758 147628 317902
rect 148152 317490 148180 320076
rect 148612 318782 148640 320076
rect 148600 318776 148652 318782
rect 148600 318718 148652 318724
rect 148876 317960 148928 317966
rect 148876 317902 148928 317908
rect 148416 317824 148468 317830
rect 148416 317766 148468 317772
rect 148324 317620 148376 317626
rect 148324 317562 148376 317568
rect 148140 317484 148192 317490
rect 148140 317426 148192 317432
rect 147588 4752 147640 4758
rect 147588 4694 147640 4700
rect 146208 4684 146260 4690
rect 146208 4626 146260 4632
rect 148336 4146 148364 317562
rect 148324 4140 148376 4146
rect 148324 4082 148376 4088
rect 145840 3324 145892 3330
rect 145840 3266 145892 3272
rect 148048 3324 148100 3330
rect 148048 3266 148100 3272
rect 145656 3256 145708 3262
rect 145656 3198 145708 3204
rect 145564 2916 145616 2922
rect 145564 2858 145616 2864
rect 145668 480 145696 3198
rect 146850 2952 146906 2961
rect 146850 2887 146906 2896
rect 146864 480 146892 2887
rect 148060 480 148088 3266
rect 148428 2854 148456 317766
rect 148888 7682 148916 317902
rect 149072 317830 149100 320076
rect 149060 317824 149112 317830
rect 149060 317766 149112 317772
rect 149532 317490 149560 320076
rect 149900 318714 149928 320076
rect 150360 318782 150388 320076
rect 150348 318776 150400 318782
rect 150348 318718 150400 318724
rect 149888 318708 149940 318714
rect 149888 318650 149940 318656
rect 149702 318472 149758 318481
rect 149702 318407 149758 318416
rect 149716 318209 149744 318407
rect 149702 318200 149758 318209
rect 149702 318135 149758 318144
rect 150820 317490 150848 320076
rect 151294 320062 151584 320090
rect 151084 317552 151136 317558
rect 151084 317494 151136 317500
rect 148968 317484 149020 317490
rect 148968 317426 149020 317432
rect 149520 317484 149572 317490
rect 149520 317426 149572 317432
rect 150164 317484 150216 317490
rect 150164 317426 150216 317432
rect 150808 317484 150860 317490
rect 150808 317426 150860 317432
rect 148876 7676 148928 7682
rect 148876 7618 148928 7624
rect 148980 5506 149008 317426
rect 150176 311794 150204 317426
rect 150176 311766 150296 311794
rect 150268 302274 150296 311766
rect 150268 302246 150388 302274
rect 150360 282946 150388 302246
rect 150164 282940 150216 282946
rect 150164 282882 150216 282888
rect 150348 282940 150400 282946
rect 150348 282882 150400 282888
rect 150176 282826 150204 282882
rect 150176 282798 150296 282826
rect 150268 273306 150296 282798
rect 150268 273278 150388 273306
rect 150360 263634 150388 273278
rect 150164 263628 150216 263634
rect 150164 263570 150216 263576
rect 150348 263628 150400 263634
rect 150348 263570 150400 263576
rect 150176 263514 150204 263570
rect 150176 263486 150296 263514
rect 150268 253994 150296 263486
rect 150268 253966 150388 253994
rect 150360 244322 150388 253966
rect 150164 244316 150216 244322
rect 150164 244258 150216 244264
rect 150348 244316 150400 244322
rect 150348 244258 150400 244264
rect 150176 244202 150204 244258
rect 150176 244174 150296 244202
rect 150268 234682 150296 244174
rect 150268 234654 150388 234682
rect 150360 225010 150388 234654
rect 150164 225004 150216 225010
rect 150164 224946 150216 224952
rect 150348 225004 150400 225010
rect 150348 224946 150400 224952
rect 150176 224890 150204 224946
rect 150176 224862 150296 224890
rect 150268 215370 150296 224862
rect 150268 215342 150388 215370
rect 150360 205698 150388 215342
rect 150164 205692 150216 205698
rect 150164 205634 150216 205640
rect 150348 205692 150400 205698
rect 150348 205634 150400 205640
rect 150176 205578 150204 205634
rect 150176 205550 150296 205578
rect 150268 196058 150296 205550
rect 150268 196030 150388 196058
rect 150360 186386 150388 196030
rect 150164 186380 150216 186386
rect 150164 186322 150216 186328
rect 150348 186380 150400 186386
rect 150348 186322 150400 186328
rect 150176 186266 150204 186322
rect 150176 186238 150296 186266
rect 150268 183569 150296 186238
rect 150070 183560 150126 183569
rect 150070 183495 150126 183504
rect 150254 183560 150310 183569
rect 150254 183495 150310 183504
rect 150084 173942 150112 183495
rect 150072 173936 150124 173942
rect 150072 173878 150124 173884
rect 150348 173936 150400 173942
rect 150348 173878 150400 173884
rect 150360 167074 150388 173878
rect 150164 167068 150216 167074
rect 150164 167010 150216 167016
rect 150348 167068 150400 167074
rect 150348 167010 150400 167016
rect 150176 166954 150204 167010
rect 150176 166926 150296 166954
rect 150268 164218 150296 166926
rect 150256 164212 150308 164218
rect 150256 164154 150308 164160
rect 150256 157344 150308 157350
rect 150256 157286 150308 157292
rect 150268 154578 150296 157286
rect 150268 154550 150388 154578
rect 150360 147694 150388 154550
rect 150164 147688 150216 147694
rect 150348 147688 150400 147694
rect 150216 147636 150296 147642
rect 150164 147630 150296 147636
rect 150348 147630 150400 147636
rect 150176 147614 150296 147630
rect 150268 144906 150296 147614
rect 150256 144900 150308 144906
rect 150256 144842 150308 144848
rect 150256 137964 150308 137970
rect 150256 137906 150308 137912
rect 150268 135266 150296 137906
rect 150268 135238 150388 135266
rect 150360 128382 150388 135238
rect 150164 128376 150216 128382
rect 150348 128376 150400 128382
rect 150216 128324 150296 128330
rect 150164 128318 150296 128324
rect 150348 128318 150400 128324
rect 150176 128302 150296 128318
rect 150268 125594 150296 128302
rect 150256 125588 150308 125594
rect 150256 125530 150308 125536
rect 150256 118652 150308 118658
rect 150256 118594 150308 118600
rect 150268 115954 150296 118594
rect 150268 115926 150388 115954
rect 150360 109070 150388 115926
rect 150164 109064 150216 109070
rect 150348 109064 150400 109070
rect 150216 109012 150296 109018
rect 150164 109006 150296 109012
rect 150348 109006 150400 109012
rect 150176 108990 150296 109006
rect 150268 106282 150296 108990
rect 150256 106276 150308 106282
rect 150256 106218 150308 106224
rect 150256 99340 150308 99346
rect 150256 99282 150308 99288
rect 150268 96642 150296 99282
rect 150268 96614 150388 96642
rect 150360 89758 150388 96614
rect 150164 89752 150216 89758
rect 150348 89752 150400 89758
rect 150216 89700 150296 89706
rect 150164 89694 150296 89700
rect 150348 89694 150400 89700
rect 150176 89678 150296 89694
rect 150268 86970 150296 89678
rect 150256 86964 150308 86970
rect 150256 86906 150308 86912
rect 150348 77308 150400 77314
rect 150348 77250 150400 77256
rect 150360 77217 150388 77250
rect 150162 77208 150218 77217
rect 150162 77143 150218 77152
rect 150346 77208 150402 77217
rect 150346 77143 150402 77152
rect 150176 70446 150204 77143
rect 150164 70440 150216 70446
rect 150164 70382 150216 70388
rect 150256 70372 150308 70378
rect 150256 70314 150308 70320
rect 150268 60738 150296 70314
rect 150268 60710 150388 60738
rect 150360 57934 150388 60710
rect 150348 57928 150400 57934
rect 150348 57870 150400 57876
rect 150256 48340 150308 48346
rect 150256 48282 150308 48288
rect 150268 41426 150296 48282
rect 150268 41398 150388 41426
rect 150360 38622 150388 41398
rect 150348 38616 150400 38622
rect 150348 38558 150400 38564
rect 150256 29028 150308 29034
rect 150256 28970 150308 28976
rect 150268 22114 150296 28970
rect 150268 22086 150388 22114
rect 150360 12458 150388 22086
rect 150176 12430 150388 12458
rect 148968 5500 149020 5506
rect 148968 5442 149020 5448
rect 150176 5438 150204 12430
rect 150164 5432 150216 5438
rect 150164 5374 150216 5380
rect 151096 3738 151124 317494
rect 151556 8770 151584 320062
rect 151648 320062 151754 320090
rect 151648 8906 151676 320062
rect 152200 317490 152228 320076
rect 152674 320062 153056 320090
rect 152292 317762 152504 317778
rect 152280 317756 152504 317762
rect 152332 317750 152504 317756
rect 152280 317698 152332 317704
rect 151728 317484 151780 317490
rect 151728 317426 151780 317432
rect 152188 317484 152240 317490
rect 152188 317426 152240 317432
rect 151636 8900 151688 8906
rect 151636 8842 151688 8848
rect 151544 8764 151596 8770
rect 151544 8706 151596 8712
rect 151740 5370 151768 317426
rect 151728 5364 151780 5370
rect 151728 5306 151780 5312
rect 152476 4146 152504 317750
rect 152556 317688 152608 317694
rect 152556 317630 152608 317636
rect 151544 4140 151596 4146
rect 151544 4082 151596 4088
rect 152464 4140 152516 4146
rect 152464 4082 152516 4088
rect 150440 3732 150492 3738
rect 150440 3674 150492 3680
rect 151084 3732 151136 3738
rect 151084 3674 151136 3680
rect 149244 3052 149296 3058
rect 149244 2994 149296 3000
rect 148416 2848 148468 2854
rect 148416 2790 148468 2796
rect 149256 480 149284 2994
rect 150452 480 150480 3674
rect 151556 480 151584 4082
rect 152568 3262 152596 317630
rect 153028 8838 153056 320062
rect 153120 317898 153148 320076
rect 153108 317892 153160 317898
rect 153108 317834 153160 317840
rect 153488 317490 153516 320076
rect 153962 320062 154344 320090
rect 153844 318096 153896 318102
rect 153844 318038 153896 318044
rect 153108 317484 153160 317490
rect 153108 317426 153160 317432
rect 153476 317484 153528 317490
rect 153476 317426 153528 317432
rect 153016 8832 153068 8838
rect 153016 8774 153068 8780
rect 153120 5302 153148 317426
rect 153108 5296 153160 5302
rect 153108 5238 153160 5244
rect 153856 4078 153884 318038
rect 154316 9654 154344 320062
rect 154304 9648 154356 9654
rect 154304 9590 154356 9596
rect 154408 9586 154436 320076
rect 154868 317490 154896 320076
rect 155328 318102 155356 320076
rect 155788 318646 155816 320076
rect 155776 318640 155828 318646
rect 155776 318582 155828 318588
rect 155316 318096 155368 318102
rect 155316 318038 155368 318044
rect 155776 318096 155828 318102
rect 155776 318038 155828 318044
rect 155224 317824 155276 317830
rect 155224 317766 155276 317772
rect 154488 317484 154540 317490
rect 154488 317426 154540 317432
rect 154856 317484 154908 317490
rect 154856 317426 154908 317432
rect 154396 9580 154448 9586
rect 154396 9522 154448 9528
rect 154500 5234 154528 317426
rect 154488 5228 154540 5234
rect 154488 5170 154540 5176
rect 155236 4146 155264 317766
rect 155788 9518 155816 318038
rect 156248 317558 156276 320076
rect 156708 317626 156736 320076
rect 157090 320062 157196 320090
rect 156604 317620 156656 317626
rect 156604 317562 156656 317568
rect 156696 317620 156748 317626
rect 156696 317562 156748 317568
rect 157064 317620 157116 317626
rect 157064 317562 157116 317568
rect 156236 317552 156288 317558
rect 156236 317494 156288 317500
rect 155868 317484 155920 317490
rect 155868 317426 155920 317432
rect 155776 9512 155828 9518
rect 155776 9454 155828 9460
rect 155880 5166 155908 317426
rect 155868 5160 155920 5166
rect 155868 5102 155920 5108
rect 155132 4140 155184 4146
rect 155132 4082 155184 4088
rect 155224 4140 155276 4146
rect 155224 4082 155276 4088
rect 153844 4072 153896 4078
rect 153844 4014 153896 4020
rect 152556 3256 152608 3262
rect 152556 3198 152608 3204
rect 152740 3188 152792 3194
rect 152740 3130 152792 3136
rect 152752 480 152780 3130
rect 153934 3088 153990 3097
rect 153934 3023 153990 3032
rect 153948 480 153976 3023
rect 155144 480 155172 4082
rect 156328 3324 156380 3330
rect 156328 3266 156380 3272
rect 156340 480 156368 3266
rect 156616 2854 156644 317562
rect 157076 9450 157104 317562
rect 157064 9444 157116 9450
rect 157064 9386 157116 9392
rect 157168 9382 157196 320062
rect 157536 317626 157564 320076
rect 157890 318200 157946 318209
rect 157890 318135 157946 318144
rect 157524 317620 157576 317626
rect 157524 317562 157576 317568
rect 157248 317552 157300 317558
rect 157248 317494 157300 317500
rect 157156 9376 157208 9382
rect 157156 9318 157208 9324
rect 157260 5098 157288 317494
rect 157904 311794 157932 318135
rect 157996 317490 158024 320076
rect 157984 317484 158036 317490
rect 157984 317426 158036 317432
rect 157904 311766 158024 311794
rect 157248 5092 157300 5098
rect 157248 5034 157300 5040
rect 157996 3738 158024 311766
rect 158456 9314 158484 320076
rect 158916 317626 158944 320076
rect 158628 317620 158680 317626
rect 158628 317562 158680 317568
rect 158904 317620 158956 317626
rect 158904 317562 158956 317568
rect 158536 317484 158588 317490
rect 158536 317426 158588 317432
rect 158444 9308 158496 9314
rect 158444 9250 158496 9256
rect 158548 6254 158576 317426
rect 158536 6248 158588 6254
rect 158536 6190 158588 6196
rect 158640 5030 158668 317562
rect 159376 317490 159404 320076
rect 159456 317756 159508 317762
rect 159456 317698 159508 317704
rect 159364 317484 159416 317490
rect 159364 317426 159416 317432
rect 159364 317348 159416 317354
rect 159364 317290 159416 317296
rect 158628 5024 158680 5030
rect 158628 4966 158680 4972
rect 157984 3732 158036 3738
rect 157984 3674 158036 3680
rect 158718 3496 158774 3505
rect 158718 3431 158774 3440
rect 157524 3188 157576 3194
rect 157524 3130 157576 3136
rect 156604 2848 156656 2854
rect 156604 2790 156656 2796
rect 157536 480 157564 3130
rect 158732 480 158760 3431
rect 159376 3097 159404 317290
rect 159468 3874 159496 317698
rect 159836 9246 159864 320076
rect 160008 317620 160060 317626
rect 160008 317562 160060 317568
rect 159916 317484 159968 317490
rect 159916 317426 159968 317432
rect 159824 9240 159876 9246
rect 159824 9182 159876 9188
rect 159928 6186 159956 317426
rect 159916 6180 159968 6186
rect 159916 6122 159968 6128
rect 160020 4962 160048 317562
rect 160296 317558 160324 320076
rect 160376 317756 160428 317762
rect 160376 317698 160428 317704
rect 160284 317552 160336 317558
rect 160284 317494 160336 317500
rect 160388 12442 160416 317698
rect 160756 317490 160784 320076
rect 161138 320062 161244 320090
rect 160744 317484 160796 317490
rect 160744 317426 160796 317432
rect 160744 309188 160796 309194
rect 160744 309130 160796 309136
rect 160756 202881 160784 309130
rect 160558 202872 160614 202881
rect 160558 202807 160614 202816
rect 160742 202872 160798 202881
rect 160742 202807 160798 202816
rect 160572 193254 160600 202807
rect 160560 193248 160612 193254
rect 160560 193190 160612 193196
rect 160744 193248 160796 193254
rect 160744 193190 160796 193196
rect 160756 86902 160784 193190
rect 160744 86896 160796 86902
rect 160744 86838 160796 86844
rect 160744 77308 160796 77314
rect 160744 77250 160796 77256
rect 160756 28914 160784 77250
rect 160664 28886 160784 28914
rect 160664 19378 160692 28886
rect 160652 19372 160704 19378
rect 160652 19314 160704 19320
rect 160744 19372 160796 19378
rect 160744 19314 160796 19320
rect 160376 12436 160428 12442
rect 160376 12378 160428 12384
rect 160008 4956 160060 4962
rect 160008 4898 160060 4904
rect 159916 4004 159968 4010
rect 159916 3946 159968 3952
rect 159456 3868 159508 3874
rect 159456 3810 159508 3816
rect 159362 3088 159418 3097
rect 159362 3023 159418 3032
rect 159928 480 159956 3946
rect 160756 3126 160784 19314
rect 161112 12436 161164 12442
rect 161112 12378 161164 12384
rect 160744 3120 160796 3126
rect 160744 3062 160796 3068
rect 161124 480 161152 12378
rect 161216 9178 161244 320062
rect 161388 317552 161440 317558
rect 161388 317494 161440 317500
rect 161296 317484 161348 317490
rect 161296 317426 161348 317432
rect 161204 9172 161256 9178
rect 161204 9114 161256 9120
rect 161308 7002 161336 317426
rect 161296 6996 161348 7002
rect 161296 6938 161348 6944
rect 161400 4894 161428 317494
rect 161584 317490 161612 320076
rect 162044 317558 162072 320076
rect 162124 318708 162176 318714
rect 162124 318650 162176 318656
rect 162032 317552 162084 317558
rect 162032 317494 162084 317500
rect 161572 317484 161624 317490
rect 161572 317426 161624 317432
rect 161388 4888 161440 4894
rect 161388 4830 161440 4836
rect 162136 3505 162164 318650
rect 162504 317762 162532 320076
rect 162492 317756 162544 317762
rect 162492 317698 162544 317704
rect 162676 317552 162728 317558
rect 162676 317494 162728 317500
rect 162688 9110 162716 317494
rect 162964 317490 162992 320076
rect 163424 317558 163452 320076
rect 163884 318714 163912 320076
rect 163872 318708 163924 318714
rect 163872 318650 163924 318656
rect 164344 317558 164372 320076
rect 163412 317552 163464 317558
rect 163412 317494 163464 317500
rect 164056 317552 164108 317558
rect 164056 317494 164108 317500
rect 164332 317552 164384 317558
rect 164332 317494 164384 317500
rect 162768 317484 162820 317490
rect 162768 317426 162820 317432
rect 162952 317484 163004 317490
rect 162952 317426 163004 317432
rect 162676 9104 162728 9110
rect 162676 9046 162728 9052
rect 162780 4826 162808 317426
rect 164068 9042 164096 317494
rect 164712 317490 164740 320076
rect 165172 318374 165200 320076
rect 164884 318368 164936 318374
rect 164884 318310 164936 318316
rect 165160 318368 165212 318374
rect 165160 318310 165212 318316
rect 164148 317484 164200 317490
rect 164148 317426 164200 317432
rect 164700 317484 164752 317490
rect 164700 317426 164752 317432
rect 164056 9036 164108 9042
rect 164056 8978 164108 8984
rect 163504 6044 163556 6050
rect 163504 5986 163556 5992
rect 162768 4820 162820 4826
rect 162768 4762 162820 4768
rect 162306 3632 162362 3641
rect 162306 3567 162362 3576
rect 162122 3496 162178 3505
rect 162122 3431 162178 3440
rect 162320 480 162348 3567
rect 162766 3496 162822 3505
rect 162766 3431 162822 3440
rect 162780 3097 162808 3431
rect 162766 3088 162822 3097
rect 162766 3023 162822 3032
rect 163516 480 163544 5986
rect 164160 5137 164188 317426
rect 164146 5128 164202 5137
rect 164146 5063 164202 5072
rect 164700 3868 164752 3874
rect 164700 3810 164752 3816
rect 164712 480 164740 3810
rect 164896 3126 164924 318310
rect 165528 317552 165580 317558
rect 165528 317494 165580 317500
rect 165436 317484 165488 317490
rect 165436 317426 165488 317432
rect 165448 8974 165476 317426
rect 165436 8968 165488 8974
rect 165436 8910 165488 8916
rect 165540 5001 165568 317494
rect 165632 317490 165660 320076
rect 166092 317626 166120 320076
rect 166356 318300 166408 318306
rect 166356 318242 166408 318248
rect 166264 318028 166316 318034
rect 166264 317970 166316 317976
rect 166080 317620 166132 317626
rect 166080 317562 166132 317568
rect 165620 317484 165672 317490
rect 165620 317426 165672 317432
rect 165526 4992 165582 5001
rect 165526 4927 165582 4936
rect 166276 3874 166304 317970
rect 166264 3868 166316 3874
rect 166264 3810 166316 3816
rect 166368 3398 166396 318242
rect 166552 317558 166580 320076
rect 167012 318170 167040 320076
rect 167000 318164 167052 318170
rect 167000 318106 167052 318112
rect 167472 318102 167500 320076
rect 167644 318436 167696 318442
rect 167644 318378 167696 318384
rect 167460 318096 167512 318102
rect 167460 318038 167512 318044
rect 166816 317620 166868 317626
rect 166816 317562 166868 317568
rect 166540 317552 166592 317558
rect 166540 317494 166592 317500
rect 166828 8362 166856 317562
rect 166908 317484 166960 317490
rect 166908 317426 166960 317432
rect 166816 8356 166868 8362
rect 166816 8298 166868 8304
rect 166920 4865 166948 317426
rect 167092 6112 167144 6118
rect 167092 6054 167144 6060
rect 166906 4856 166962 4865
rect 166906 4791 166962 4800
rect 166356 3392 166408 3398
rect 166356 3334 166408 3340
rect 164884 3120 164936 3126
rect 164884 3062 164936 3068
rect 165896 2916 165948 2922
rect 165896 2858 165948 2864
rect 165908 480 165936 2858
rect 167104 480 167132 6054
rect 167656 4010 167684 318378
rect 167932 318034 167960 320076
rect 168116 320062 168314 320090
rect 167920 318028 167972 318034
rect 167920 317970 167972 317976
rect 168116 13870 168144 320062
rect 168288 318164 168340 318170
rect 168288 318106 168340 318112
rect 168196 318096 168248 318102
rect 168196 318038 168248 318044
rect 168104 13864 168156 13870
rect 168104 13806 168156 13812
rect 168208 8430 168236 318038
rect 168196 8424 168248 8430
rect 168196 8366 168248 8372
rect 168300 5545 168328 318106
rect 168760 318102 168788 320076
rect 169024 318572 169076 318578
rect 169024 318514 169076 318520
rect 168748 318096 168800 318102
rect 168748 318038 168800 318044
rect 168286 5536 168342 5545
rect 168286 5471 168342 5480
rect 169036 4010 169064 318514
rect 169220 318034 169248 320076
rect 169576 318096 169628 318102
rect 169576 318038 169628 318044
rect 169208 318028 169260 318034
rect 169208 317970 169260 317976
rect 169588 8498 169616 318038
rect 169576 8492 169628 8498
rect 169576 8434 169628 8440
rect 169680 5409 169708 320076
rect 170140 317966 170168 320076
rect 170600 318510 170628 320076
rect 170968 320062 171074 320090
rect 170588 318504 170640 318510
rect 170588 318446 170640 318452
rect 170128 317960 170180 317966
rect 170128 317902 170180 317908
rect 170968 14006 170996 320062
rect 171048 317960 171100 317966
rect 171048 317902 171100 317908
rect 170956 14000 171008 14006
rect 170956 13942 171008 13948
rect 171060 8566 171088 317902
rect 171520 317490 171548 320076
rect 171980 318442 172008 320076
rect 172362 320062 172468 320090
rect 171968 318436 172020 318442
rect 171968 318378 172020 318384
rect 171784 317688 171836 317694
rect 171784 317630 171836 317636
rect 171508 317484 171560 317490
rect 171508 317426 171560 317432
rect 171048 8560 171100 8566
rect 171048 8502 171100 8508
rect 170588 6860 170640 6866
rect 170588 6802 170640 6808
rect 169666 5400 169722 5409
rect 169666 5335 169722 5344
rect 167644 4004 167696 4010
rect 167644 3946 167696 3952
rect 169024 4004 169076 4010
rect 169024 3946 169076 3952
rect 168196 3936 168248 3942
rect 168196 3878 168248 3884
rect 169944 3936 169996 3942
rect 169944 3878 169996 3884
rect 168208 480 168236 3878
rect 169956 3806 169984 3878
rect 169944 3800 169996 3806
rect 169944 3742 169996 3748
rect 169390 3224 169446 3233
rect 169390 3159 169446 3168
rect 169404 480 169432 3159
rect 170600 480 170628 6802
rect 171796 3097 171824 317630
rect 172336 317484 172388 317490
rect 172336 317426 172388 317432
rect 172348 13938 172376 317426
rect 172336 13932 172388 13938
rect 172336 13874 172388 13880
rect 172440 5574 172468 320062
rect 172808 317966 172836 320076
rect 172796 317960 172848 317966
rect 172796 317902 172848 317908
rect 173268 317830 173296 320076
rect 173742 320062 173848 320090
rect 173716 317960 173768 317966
rect 173716 317902 173768 317908
rect 173164 317824 173216 317830
rect 173164 317766 173216 317772
rect 173256 317824 173308 317830
rect 173256 317766 173308 317772
rect 172428 5568 172480 5574
rect 172428 5510 172480 5516
rect 172334 4856 172390 4865
rect 172518 4856 172574 4865
rect 172390 4814 172518 4842
rect 172334 4791 172390 4800
rect 172518 4791 172574 4800
rect 172980 3936 173032 3942
rect 172980 3878 173032 3884
rect 171782 3088 171838 3097
rect 171782 3023 171838 3032
rect 171784 2984 171836 2990
rect 171784 2926 171836 2932
rect 171796 480 171824 2926
rect 172992 480 173020 3878
rect 173176 2990 173204 317766
rect 173728 14074 173756 317902
rect 173716 14068 173768 14074
rect 173716 14010 173768 14016
rect 173820 5642 173848 320062
rect 174188 317966 174216 320076
rect 174648 318374 174676 320076
rect 175122 320062 175228 320090
rect 174636 318368 174688 318374
rect 174636 318310 174688 318316
rect 174176 317960 174228 317966
rect 174176 317902 174228 317908
rect 175096 317960 175148 317966
rect 175096 317902 175148 317908
rect 175108 14142 175136 317902
rect 175096 14136 175148 14142
rect 175096 14078 175148 14084
rect 174176 6792 174228 6798
rect 174176 6734 174228 6740
rect 173808 5636 173860 5642
rect 173808 5578 173860 5584
rect 173164 2984 173216 2990
rect 173164 2926 173216 2932
rect 174188 480 174216 6734
rect 175200 5710 175228 320062
rect 175568 317490 175596 320076
rect 175832 318776 175884 318782
rect 175832 318718 175884 318724
rect 175844 318186 175872 318718
rect 175936 318306 175964 320076
rect 176410 320062 176608 320090
rect 175924 318300 175976 318306
rect 175924 318242 175976 318248
rect 175844 318158 175964 318186
rect 175556 317484 175608 317490
rect 175556 317426 175608 317432
rect 175936 6118 175964 318158
rect 176016 317892 176068 317898
rect 176016 317834 176068 317840
rect 175924 6112 175976 6118
rect 175924 6054 175976 6060
rect 175188 5704 175240 5710
rect 175188 5646 175240 5652
rect 176028 3738 176056 317834
rect 176476 317484 176528 317490
rect 176476 317426 176528 317432
rect 176488 14210 176516 317426
rect 176476 14204 176528 14210
rect 176476 14146 176528 14152
rect 176580 5778 176608 320062
rect 176856 317966 176884 320076
rect 177316 318578 177344 320076
rect 177790 320062 177988 320090
rect 177304 318572 177356 318578
rect 177304 318514 177356 318520
rect 176844 317960 176896 317966
rect 176844 317902 176896 317908
rect 177856 317960 177908 317966
rect 177856 317902 177908 317908
rect 177868 9722 177896 317902
rect 177856 9716 177908 9722
rect 177856 9658 177908 9664
rect 177764 6724 177816 6730
rect 177764 6666 177816 6672
rect 176568 5772 176620 5778
rect 176568 5714 176620 5720
rect 176566 4312 176622 4321
rect 176566 4247 176622 4256
rect 176750 4312 176806 4321
rect 176750 4247 176806 4256
rect 176474 4176 176530 4185
rect 176474 4111 176530 4120
rect 176488 4010 176516 4111
rect 176476 4004 176528 4010
rect 176476 3946 176528 3952
rect 176580 3874 176608 4247
rect 176764 3874 176792 4247
rect 176842 4176 176898 4185
rect 176842 4111 176898 4120
rect 176856 3942 176884 4111
rect 176844 3936 176896 3942
rect 176844 3878 176896 3884
rect 176568 3868 176620 3874
rect 176568 3810 176620 3816
rect 176752 3868 176804 3874
rect 176752 3810 176804 3816
rect 176016 3732 176068 3738
rect 176016 3674 176068 3680
rect 176936 3732 176988 3738
rect 176936 3674 176988 3680
rect 176948 3618 176976 3674
rect 176672 3590 176976 3618
rect 176672 3262 176700 3590
rect 176660 3256 176712 3262
rect 176660 3198 176712 3204
rect 175372 3120 175424 3126
rect 175372 3062 175424 3068
rect 176750 3088 176806 3097
rect 175384 480 175412 3062
rect 176568 3052 176620 3058
rect 176750 3023 176806 3032
rect 176568 2994 176620 3000
rect 176580 480 176608 2994
rect 176764 2990 176792 3023
rect 176752 2984 176804 2990
rect 176752 2926 176804 2932
rect 177776 480 177804 6666
rect 177960 5846 177988 320062
rect 178236 317966 178264 320076
rect 178592 318640 178644 318646
rect 178592 318582 178644 318588
rect 178604 318050 178632 318582
rect 178696 318209 178724 320076
rect 179170 320062 179368 320090
rect 178682 318200 178738 318209
rect 178682 318135 178738 318144
rect 178604 318022 178724 318050
rect 178224 317960 178276 317966
rect 178224 317902 178276 317908
rect 177948 5840 178000 5846
rect 177948 5782 178000 5788
rect 178696 4185 178724 318022
rect 179236 317960 179288 317966
rect 179236 317902 179288 317908
rect 179248 9790 179276 317902
rect 179236 9784 179288 9790
rect 179236 9726 179288 9732
rect 179340 5914 179368 320062
rect 179524 317966 179552 320076
rect 179512 317960 179564 317966
rect 179512 317902 179564 317908
rect 179984 317490 180012 320076
rect 180458 320062 180748 320090
rect 180616 317960 180668 317966
rect 180616 317902 180668 317908
rect 180064 317756 180116 317762
rect 180064 317698 180116 317704
rect 179972 317484 180024 317490
rect 179972 317426 180024 317432
rect 179328 5908 179380 5914
rect 179328 5850 179380 5856
rect 178682 4176 178738 4185
rect 178682 4111 178738 4120
rect 180076 3398 180104 317698
rect 180524 317484 180576 317490
rect 180524 317426 180576 317432
rect 180536 15570 180564 317426
rect 180524 15564 180576 15570
rect 180524 15506 180576 15512
rect 180628 9858 180656 317902
rect 180616 9852 180668 9858
rect 180616 9794 180668 9800
rect 180720 5982 180748 320062
rect 180904 317830 180932 320076
rect 181364 318073 181392 320076
rect 181838 320062 182128 320090
rect 181350 318064 181406 318073
rect 181350 317999 181406 318008
rect 180892 317824 180944 317830
rect 180892 317766 180944 317772
rect 181996 317824 182048 317830
rect 181996 317766 182048 317772
rect 182008 9926 182036 317766
rect 181996 9920 182048 9926
rect 181996 9862 182048 9868
rect 181352 6656 181404 6662
rect 181352 6598 181404 6604
rect 180708 5976 180760 5982
rect 180708 5918 180760 5924
rect 180706 4856 180762 4865
rect 180706 4791 180762 4800
rect 180720 4593 180748 4791
rect 180706 4584 180762 4593
rect 180706 4519 180762 4528
rect 178960 3392 179012 3398
rect 178960 3334 179012 3340
rect 180064 3392 180116 3398
rect 180064 3334 180116 3340
rect 178972 480 179000 3334
rect 180156 2780 180208 2786
rect 180156 2722 180208 2728
rect 180168 480 180196 2722
rect 181364 480 181392 6598
rect 182100 6050 182128 320062
rect 182284 318034 182312 320076
rect 182272 318028 182324 318034
rect 182272 317970 182324 317976
rect 182744 317626 182772 320076
rect 183218 320062 183508 320090
rect 183376 318028 183428 318034
rect 183376 317970 183428 317976
rect 182824 317688 182876 317694
rect 182824 317630 182876 317636
rect 182732 317620 182784 317626
rect 182732 317562 182784 317568
rect 182088 6044 182140 6050
rect 182088 5986 182140 5992
rect 182086 4856 182142 4865
rect 182086 4791 182142 4800
rect 182100 4593 182128 4791
rect 182086 4584 182142 4593
rect 182086 4519 182142 4528
rect 181534 4176 181590 4185
rect 181534 4111 181590 4120
rect 181548 3806 181576 4111
rect 182548 4004 182600 4010
rect 182548 3946 182600 3952
rect 181536 3800 181588 3806
rect 181536 3742 181588 3748
rect 182560 480 182588 3946
rect 182836 3398 182864 317630
rect 183388 9994 183416 317970
rect 183376 9988 183428 9994
rect 183376 9930 183428 9936
rect 183480 6118 183508 320062
rect 183572 318034 183600 320076
rect 184046 320062 184336 320090
rect 184506 320062 184888 320090
rect 183560 318028 183612 318034
rect 183560 317970 183612 317976
rect 184308 317966 184336 320062
rect 184756 318028 184808 318034
rect 184756 317970 184808 317976
rect 184204 317960 184256 317966
rect 184204 317902 184256 317908
rect 184296 317960 184348 317966
rect 184296 317902 184348 317908
rect 183468 6112 183520 6118
rect 183468 6054 183520 6060
rect 184216 3738 184244 317902
rect 184768 10062 184796 317970
rect 184756 10056 184808 10062
rect 184756 9998 184808 10004
rect 184860 6866 184888 320062
rect 184952 318034 184980 320076
rect 184940 318028 184992 318034
rect 184940 317970 184992 317976
rect 185412 317830 185440 320076
rect 185886 320062 186268 320090
rect 186136 318028 186188 318034
rect 186136 317970 186188 317976
rect 185584 317892 185636 317898
rect 185584 317834 185636 317840
rect 185400 317824 185452 317830
rect 185400 317766 185452 317772
rect 184848 6860 184900 6866
rect 184848 6802 184900 6808
rect 184848 6588 184900 6594
rect 184848 6530 184900 6536
rect 183744 3732 183796 3738
rect 183744 3674 183796 3680
rect 184204 3732 184256 3738
rect 184204 3674 184256 3680
rect 182824 3392 182876 3398
rect 182824 3334 182876 3340
rect 183756 480 183784 3674
rect 184860 480 184888 6530
rect 185596 3806 185624 317834
rect 186148 10130 186176 317970
rect 186136 10124 186188 10130
rect 186136 10066 186188 10072
rect 186240 6798 186268 320062
rect 186332 318034 186360 320076
rect 186792 318646 186820 320076
rect 186780 318640 186832 318646
rect 186780 318582 186832 318588
rect 186320 318028 186372 318034
rect 186320 317970 186372 317976
rect 187160 317966 187188 320076
rect 187528 320062 187634 320090
rect 187424 318028 187476 318034
rect 187424 317970 187476 317976
rect 187148 317960 187200 317966
rect 187148 317902 187200 317908
rect 187436 10198 187464 317970
rect 187528 10266 187556 320062
rect 187608 317960 187660 317966
rect 187608 317902 187660 317908
rect 187516 10260 187568 10266
rect 187516 10202 187568 10208
rect 187424 10192 187476 10198
rect 187424 10134 187476 10140
rect 186228 6792 186280 6798
rect 186228 6734 186280 6740
rect 187620 6730 187648 317902
rect 188080 317762 188108 320076
rect 188540 318034 188568 320076
rect 188908 320062 189014 320090
rect 189474 320062 189856 320090
rect 188528 318028 188580 318034
rect 188528 317970 188580 317976
rect 188068 317756 188120 317762
rect 188068 317698 188120 317704
rect 188908 11014 188936 320062
rect 189080 318572 189132 318578
rect 189080 318514 189132 318520
rect 188988 318028 189040 318034
rect 188988 317970 189040 317976
rect 188896 11008 188948 11014
rect 188896 10950 188948 10956
rect 187608 6724 187660 6730
rect 187608 6666 187660 6672
rect 189000 6662 189028 317970
rect 189092 317694 189120 318514
rect 189828 317914 189856 320062
rect 189920 318034 189948 320076
rect 190288 320062 190394 320090
rect 189908 318028 189960 318034
rect 189908 317970 189960 317976
rect 189828 317886 190224 317914
rect 189724 317824 189776 317830
rect 189724 317766 189776 317772
rect 189080 317688 189132 317694
rect 189080 317630 189132 317636
rect 188988 6656 189040 6662
rect 188988 6598 189040 6604
rect 188436 6520 188488 6526
rect 188436 6462 188488 6468
rect 185584 3800 185636 3806
rect 185584 3742 185636 3748
rect 186412 3596 186464 3602
rect 186412 3538 186464 3544
rect 187240 3596 187292 3602
rect 187240 3538 187292 3544
rect 186424 3482 186452 3538
rect 186332 3454 186452 3482
rect 186136 3392 186188 3398
rect 186136 3334 186188 3340
rect 186044 3256 186096 3262
rect 186148 3233 186176 3334
rect 186332 3330 186360 3454
rect 186320 3324 186372 3330
rect 186320 3266 186372 3272
rect 186412 3324 186464 3330
rect 186412 3266 186464 3272
rect 186424 3233 186452 3266
rect 186044 3198 186096 3204
rect 186134 3224 186190 3233
rect 186056 480 186084 3198
rect 186134 3159 186190 3168
rect 186410 3224 186466 3233
rect 186410 3159 186466 3168
rect 187252 480 187280 3538
rect 188448 480 188476 6462
rect 189736 3670 189764 317766
rect 189816 317688 189868 317694
rect 189816 317630 189868 317636
rect 189828 3942 189856 317630
rect 190196 12510 190224 317886
rect 190184 12504 190236 12510
rect 190184 12446 190236 12452
rect 190288 10946 190316 320062
rect 190368 318028 190420 318034
rect 190368 317970 190420 317976
rect 190276 10940 190328 10946
rect 190276 10882 190328 10888
rect 190380 6594 190408 317970
rect 190748 317694 190776 320076
rect 191208 318034 191236 320076
rect 191576 320062 191682 320090
rect 191196 318028 191248 318034
rect 191196 317970 191248 317976
rect 190736 317688 190788 317694
rect 190736 317630 190788 317636
rect 191576 10878 191604 320062
rect 192128 318034 192156 320076
rect 191656 318028 191708 318034
rect 191656 317970 191708 317976
rect 192116 318028 192168 318034
rect 192116 317970 192168 317976
rect 191564 10872 191616 10878
rect 191564 10814 191616 10820
rect 190368 6588 190420 6594
rect 190368 6530 190420 6536
rect 191668 5273 191696 317970
rect 192588 317966 192616 320076
rect 192944 318028 192996 318034
rect 192944 317970 192996 317976
rect 192576 317960 192628 317966
rect 192576 317902 192628 317908
rect 191748 317688 191800 317694
rect 191748 317630 191800 317636
rect 191654 5264 191710 5273
rect 191654 5199 191710 5208
rect 190828 4004 190880 4010
rect 190828 3946 190880 3952
rect 189816 3936 189868 3942
rect 189816 3878 189868 3884
rect 190460 3800 190512 3806
rect 190288 3748 190460 3754
rect 190288 3742 190512 3748
rect 190288 3726 190500 3742
rect 190288 3670 190316 3726
rect 189632 3664 189684 3670
rect 189632 3606 189684 3612
rect 189724 3664 189776 3670
rect 189724 3606 189776 3612
rect 190276 3664 190328 3670
rect 190276 3606 190328 3612
rect 189644 480 189672 3606
rect 190840 480 190868 3946
rect 191760 3806 191788 317630
rect 192956 12578 192984 317970
rect 192944 12572 192996 12578
rect 192944 12514 192996 12520
rect 193048 10810 193076 320076
rect 193508 318578 193536 320076
rect 193864 318640 193916 318646
rect 193864 318582 193916 318588
rect 193496 318572 193548 318578
rect 193496 318514 193548 318520
rect 193128 317960 193180 317966
rect 193128 317902 193180 317908
rect 193036 10804 193088 10810
rect 193036 10746 193088 10752
rect 193140 6526 193168 317902
rect 193128 6520 193180 6526
rect 193128 6462 193180 6468
rect 192024 6452 192076 6458
rect 192024 6394 192076 6400
rect 191748 3800 191800 3806
rect 191748 3742 191800 3748
rect 192036 480 192064 6394
rect 193220 4072 193272 4078
rect 193220 4014 193272 4020
rect 193232 480 193260 4014
rect 193876 3874 193904 318582
rect 193968 318034 193996 320076
rect 194350 320062 194456 320090
rect 193956 318028 194008 318034
rect 193956 317970 194008 317976
rect 194428 10742 194456 320062
rect 194796 318034 194824 320076
rect 194508 318028 194560 318034
rect 194508 317970 194560 317976
rect 194784 318028 194836 318034
rect 194784 317970 194836 317976
rect 194416 10736 194468 10742
rect 194416 10678 194468 10684
rect 194520 6458 194548 317970
rect 195256 317966 195284 320076
rect 195730 320062 195836 320090
rect 195704 318028 195756 318034
rect 195704 317970 195756 317976
rect 195244 317960 195296 317966
rect 195244 317902 195296 317908
rect 195716 12646 195744 317970
rect 195704 12640 195756 12646
rect 195704 12582 195756 12588
rect 195808 10674 195836 320062
rect 196176 317966 196204 320076
rect 196636 318034 196664 320076
rect 196624 318028 196676 318034
rect 196624 317970 196676 317976
rect 195888 317960 195940 317966
rect 195888 317902 195940 317908
rect 196164 317960 196216 317966
rect 196164 317902 196216 317908
rect 195796 10668 195848 10674
rect 195796 10610 195848 10616
rect 194508 6452 194560 6458
rect 194508 6394 194560 6400
rect 195900 6390 195928 317902
rect 197096 10606 197124 320076
rect 197556 318034 197584 320076
rect 197176 318028 197228 318034
rect 197176 317970 197228 317976
rect 197544 318028 197596 318034
rect 197544 317970 197596 317976
rect 197084 10600 197136 10606
rect 197084 10542 197136 10548
rect 197188 6769 197216 317970
rect 197268 317960 197320 317966
rect 197268 317902 197320 317908
rect 197174 6760 197230 6769
rect 197174 6695 197230 6704
rect 195612 6384 195664 6390
rect 195612 6326 195664 6332
rect 195888 6384 195940 6390
rect 195888 6326 195940 6332
rect 193864 3868 193916 3874
rect 193864 3810 193916 3816
rect 194416 3664 194468 3670
rect 194416 3606 194468 3612
rect 194428 480 194456 3606
rect 195624 480 195652 6326
rect 197280 3670 197308 317902
rect 198016 317490 198044 320076
rect 198398 320062 198596 320090
rect 198464 318028 198516 318034
rect 198464 317970 198516 317976
rect 198004 317484 198056 317490
rect 198004 317426 198056 317432
rect 198476 12714 198504 317970
rect 198464 12708 198516 12714
rect 198464 12650 198516 12656
rect 198568 10538 198596 320062
rect 198844 318646 198872 320076
rect 198832 318640 198884 318646
rect 198832 318582 198884 318588
rect 199304 318034 199332 320076
rect 199778 320062 199976 320090
rect 199292 318028 199344 318034
rect 199292 317970 199344 317976
rect 198648 317484 198700 317490
rect 198648 317426 198700 317432
rect 198556 10532 198608 10538
rect 198556 10474 198608 10480
rect 198660 6633 198688 317426
rect 199948 10470 199976 320062
rect 200224 318034 200252 320076
rect 200028 318028 200080 318034
rect 200028 317970 200080 317976
rect 200212 318028 200264 318034
rect 200212 317970 200264 317976
rect 199936 10464 199988 10470
rect 199936 10406 199988 10412
rect 198646 6624 198702 6633
rect 198646 6559 198702 6568
rect 200040 6322 200068 317970
rect 200684 317966 200712 320076
rect 201158 320062 201356 320090
rect 201224 318028 201276 318034
rect 201224 317970 201276 317976
rect 200672 317960 200724 317966
rect 200672 317902 200724 317908
rect 201236 12782 201264 317970
rect 201224 12776 201276 12782
rect 201224 12718 201276 12724
rect 201328 10402 201356 320062
rect 201604 318034 201632 320076
rect 201592 318028 201644 318034
rect 201592 317970 201644 317976
rect 201408 317960 201460 317966
rect 201408 317902 201460 317908
rect 201316 10396 201368 10402
rect 201316 10338 201368 10344
rect 201420 6497 201448 317902
rect 201972 317490 202000 320076
rect 202446 320062 202736 320090
rect 202604 318028 202656 318034
rect 202604 317970 202656 317976
rect 201960 317484 202012 317490
rect 201960 317426 202012 317432
rect 202616 12850 202644 317970
rect 202604 12844 202656 12850
rect 202604 12786 202656 12792
rect 202708 10334 202736 320062
rect 202892 318034 202920 320076
rect 202880 318028 202932 318034
rect 202880 317970 202932 317976
rect 203352 317966 203380 320076
rect 203826 320062 204116 320090
rect 203984 318028 204036 318034
rect 203984 317970 204036 317976
rect 203340 317960 203392 317966
rect 203340 317902 203392 317908
rect 202788 317484 202840 317490
rect 202788 317426 202840 317432
rect 202696 10328 202748 10334
rect 202696 10270 202748 10276
rect 202800 6934 202828 317426
rect 203996 12918 204024 317970
rect 203984 12912 204036 12918
rect 203984 12854 204036 12860
rect 204088 10849 204116 320062
rect 204168 317960 204220 317966
rect 204168 317902 204220 317908
rect 204074 10840 204130 10849
rect 204074 10775 204130 10784
rect 202788 6928 202840 6934
rect 202788 6870 202840 6876
rect 201406 6488 201462 6497
rect 201406 6423 201462 6432
rect 204180 6361 204208 317902
rect 204272 317558 204300 320076
rect 204732 317694 204760 320076
rect 205206 320062 205496 320090
rect 205364 318028 205416 318034
rect 205364 317970 205416 317976
rect 204720 317688 204772 317694
rect 204720 317630 204772 317636
rect 204260 317552 204312 317558
rect 204260 317494 204312 317500
rect 205376 12986 205404 317970
rect 205364 12980 205416 12986
rect 205364 12922 205416 12928
rect 205468 10713 205496 320062
rect 205560 318034 205588 320076
rect 206020 318034 206048 320076
rect 206494 320062 206784 320090
rect 205548 318028 205600 318034
rect 205548 317970 205600 317976
rect 206008 318028 206060 318034
rect 206008 317970 206060 317976
rect 205548 317688 205600 317694
rect 205548 317630 205600 317636
rect 205454 10704 205510 10713
rect 205454 10639 205510 10648
rect 204166 6352 204222 6361
rect 199200 6316 199252 6322
rect 199200 6258 199252 6264
rect 200028 6316 200080 6322
rect 204166 6287 204222 6296
rect 200028 6258 200080 6264
rect 197268 3664 197320 3670
rect 197268 3606 197320 3612
rect 196808 3596 196860 3602
rect 196808 3538 196860 3544
rect 196820 480 196848 3538
rect 198004 2848 198056 2854
rect 198004 2790 198056 2796
rect 198016 480 198044 2790
rect 199212 480 199240 6258
rect 205454 4856 205510 4865
rect 205454 4791 205510 4800
rect 205468 4593 205496 4791
rect 205454 4584 205510 4593
rect 205454 4519 205510 4528
rect 205560 4282 205588 317630
rect 206756 8634 206784 320062
rect 206836 318028 206888 318034
rect 206836 317970 206888 317976
rect 206744 8628 206796 8634
rect 206744 8570 206796 8576
rect 206284 8220 206336 8226
rect 206284 8162 206336 8168
rect 205088 4276 205140 4282
rect 205088 4218 205140 4224
rect 205548 4276 205600 4282
rect 205548 4218 205600 4224
rect 201500 4208 201552 4214
rect 201500 4150 201552 4156
rect 200396 3732 200448 3738
rect 200396 3674 200448 3680
rect 200408 480 200436 3674
rect 201512 480 201540 4150
rect 203892 3528 203944 3534
rect 203892 3470 203944 3476
rect 202696 2916 202748 2922
rect 202696 2858 202748 2864
rect 202708 480 202736 2858
rect 203904 480 203932 3470
rect 205100 480 205128 4218
rect 206296 480 206324 8162
rect 206848 6225 206876 317970
rect 206834 6216 206890 6225
rect 206834 6151 206890 6160
rect 206940 3670 206968 320076
rect 207400 318034 207428 320076
rect 207388 318028 207440 318034
rect 207388 317970 207440 317976
rect 207860 317966 207888 320076
rect 208228 320062 208334 320090
rect 208124 318028 208176 318034
rect 208124 317970 208176 317976
rect 207848 317960 207900 317966
rect 207848 317902 207900 317908
rect 208136 14278 208164 317970
rect 208124 14272 208176 14278
rect 208124 14214 208176 14220
rect 208228 13054 208256 320062
rect 208780 318034 208808 320076
rect 209254 320062 209544 320090
rect 209622 320062 209728 320090
rect 208768 318028 208820 318034
rect 208768 317970 208820 317976
rect 208308 317960 208360 317966
rect 208308 317902 208360 317908
rect 208216 13048 208268 13054
rect 208216 12990 208268 12996
rect 208320 10577 208348 317902
rect 208306 10568 208362 10577
rect 208306 10503 208362 10512
rect 209516 10441 209544 320062
rect 209596 318028 209648 318034
rect 209596 317970 209648 317976
rect 209502 10432 209558 10441
rect 209502 10367 209558 10376
rect 209608 4350 209636 317970
rect 208676 4344 208728 4350
rect 208676 4286 208728 4292
rect 209596 4344 209648 4350
rect 209596 4286 209648 4292
rect 206928 3664 206980 3670
rect 206928 3606 206980 3612
rect 207480 3460 207532 3466
rect 207480 3402 207532 3408
rect 207492 480 207520 3402
rect 208688 480 208716 4286
rect 209700 3602 209728 320062
rect 210068 318034 210096 320076
rect 210896 318050 210924 320198
rect 210988 318782 211016 320076
rect 210976 318776 211028 318782
rect 210976 318718 211028 318724
rect 210056 318028 210108 318034
rect 210896 318022 211016 318050
rect 211448 318034 211476 320076
rect 211922 320062 212304 320090
rect 210056 317970 210108 317976
rect 210988 10305 211016 318022
rect 211068 318028 211120 318034
rect 211068 317970 211120 317976
rect 211436 318028 211488 318034
rect 211436 317970 211488 317976
rect 210974 10296 211030 10305
rect 210974 10231 211030 10240
rect 209872 8152 209924 8158
rect 209872 8094 209924 8100
rect 209688 3596 209740 3602
rect 209688 3538 209740 3544
rect 209884 480 209912 8094
rect 211080 7070 211108 317970
rect 212276 14346 212304 320062
rect 212264 14340 212316 14346
rect 212264 14282 212316 14288
rect 212368 13802 212396 320076
rect 212448 318028 212500 318034
rect 212448 317970 212500 317976
rect 212356 13796 212408 13802
rect 212356 13738 212408 13744
rect 212460 7138 212488 317970
rect 212828 317966 212856 320076
rect 213196 318034 213224 320076
rect 213184 318028 213236 318034
rect 213184 317970 213236 317976
rect 212816 317960 212868 317966
rect 212816 317902 212868 317908
rect 213656 15638 213684 320076
rect 214116 318034 214144 320076
rect 214944 318050 214972 320198
rect 215050 320062 215248 320090
rect 213736 318028 213788 318034
rect 213736 317970 213788 317976
rect 214104 318028 214156 318034
rect 214944 318022 215064 318050
rect 214104 317970 214156 317976
rect 213644 15632 213696 15638
rect 213644 15574 213696 15580
rect 213748 14414 213776 317970
rect 213828 317960 213880 317966
rect 213828 317902 213880 317908
rect 213736 14408 213788 14414
rect 213736 14350 213788 14356
rect 213460 8084 213512 8090
rect 213460 8026 213512 8032
rect 212448 7132 212500 7138
rect 212448 7074 212500 7080
rect 211068 7064 211120 7070
rect 211068 7006 211120 7012
rect 212446 4856 212502 4865
rect 212446 4791 212502 4800
rect 212460 4593 212488 4791
rect 212446 4584 212502 4593
rect 212446 4519 212502 4528
rect 212264 4412 212316 4418
rect 212264 4354 212316 4360
rect 211066 4040 211122 4049
rect 211066 3975 211122 3984
rect 211080 480 211108 3975
rect 212276 480 212304 4354
rect 213472 480 213500 8026
rect 213840 7206 213868 317902
rect 215036 15162 215064 318022
rect 215116 318028 215168 318034
rect 215116 317970 215168 317976
rect 215024 15156 215076 15162
rect 215024 15098 215076 15104
rect 215128 7274 215156 317970
rect 215116 7268 215168 7274
rect 215116 7210 215168 7216
rect 213828 7200 213880 7206
rect 213828 7142 213880 7148
rect 214654 3904 214710 3913
rect 214654 3839 214710 3848
rect 214668 480 214696 3839
rect 215220 3534 215248 320062
rect 215496 317966 215524 320076
rect 215956 318034 215984 320076
rect 215944 318028 215996 318034
rect 215944 317970 215996 317976
rect 215484 317960 215536 317966
rect 215484 317902 215536 317908
rect 216416 13734 216444 320076
rect 216784 318034 216812 320076
rect 216496 318028 216548 318034
rect 216496 317970 216548 317976
rect 216772 318028 216824 318034
rect 216772 317970 216824 317976
rect 216404 13728 216456 13734
rect 216404 13670 216456 13676
rect 216508 11150 216536 317970
rect 217244 317966 217272 320076
rect 217704 318782 217732 320076
rect 217692 318776 217744 318782
rect 217692 318718 217744 318724
rect 217968 318028 218020 318034
rect 217968 317970 218020 317976
rect 216588 317960 216640 317966
rect 216588 317902 216640 317908
rect 217232 317960 217284 317966
rect 217232 317902 217284 317908
rect 217876 317960 217928 317966
rect 217876 317902 217928 317908
rect 216496 11144 216548 11150
rect 216496 11086 216548 11092
rect 216600 7342 216628 317902
rect 217888 11218 217916 317902
rect 217876 11212 217928 11218
rect 217876 11154 217928 11160
rect 217048 8016 217100 8022
rect 217048 7958 217100 7964
rect 216588 7336 216640 7342
rect 216588 7278 216640 7284
rect 215852 4480 215904 4486
rect 215852 4422 215904 4428
rect 215208 3528 215260 3534
rect 215208 3470 215260 3476
rect 215864 480 215892 4422
rect 217060 480 217088 7958
rect 217980 7410 218008 317970
rect 218164 317966 218192 320076
rect 218152 317960 218204 317966
rect 218152 317902 218204 317908
rect 218624 317626 218652 320076
rect 219098 320062 219204 320090
rect 218612 317620 218664 317626
rect 218612 317562 218664 317568
rect 219176 15706 219204 320062
rect 219348 317960 219400 317966
rect 219348 317902 219400 317908
rect 219256 317620 219308 317626
rect 219256 317562 219308 317568
rect 219164 15700 219216 15706
rect 219164 15642 219216 15648
rect 219268 11286 219296 317562
rect 219256 11280 219308 11286
rect 219256 11222 219308 11228
rect 219360 7478 219388 317902
rect 219544 317626 219572 320076
rect 220004 317966 220032 320076
rect 220478 320062 220584 320090
rect 219992 317960 220044 317966
rect 219992 317902 220044 317908
rect 219532 317620 219584 317626
rect 219532 317562 219584 317568
rect 220556 13666 220584 320062
rect 220832 317966 220860 320076
rect 220636 317960 220688 317966
rect 220636 317902 220688 317908
rect 220820 317960 220872 317966
rect 220820 317902 220872 317908
rect 220544 13660 220596 13666
rect 220544 13602 220596 13608
rect 220648 11354 220676 317902
rect 221292 317626 221320 320076
rect 221766 320062 222148 320090
rect 222016 317960 222068 317966
rect 222016 317902 222068 317908
rect 220728 317620 220780 317626
rect 220728 317562 220780 317568
rect 221280 317620 221332 317626
rect 221280 317562 221332 317568
rect 221924 317620 221976 317626
rect 221924 317562 221976 317568
rect 220636 11348 220688 11354
rect 220636 11290 220688 11296
rect 220544 7948 220596 7954
rect 220544 7890 220596 7896
rect 219348 7472 219400 7478
rect 219348 7414 219400 7420
rect 217968 7404 218020 7410
rect 217968 7346 218020 7352
rect 219348 4548 219400 4554
rect 219348 4490 219400 4496
rect 218150 3768 218206 3777
rect 218150 3703 218206 3712
rect 218164 480 218192 3703
rect 219360 480 219388 4490
rect 220556 480 220584 7890
rect 220740 7546 220768 317562
rect 221936 11422 221964 317562
rect 221924 11416 221976 11422
rect 221924 11358 221976 11364
rect 222028 8294 222056 317902
rect 222016 8288 222068 8294
rect 222016 8230 222068 8236
rect 220728 7540 220780 7546
rect 220728 7482 220780 7488
rect 222120 3466 222148 320062
rect 222212 317626 222240 320076
rect 222672 317966 222700 320076
rect 223146 320062 223344 320090
rect 222660 317960 222712 317966
rect 222660 317902 222712 317908
rect 222200 317620 222252 317626
rect 222200 317562 222252 317568
rect 223316 15094 223344 320062
rect 223592 317966 223620 320076
rect 223396 317960 223448 317966
rect 223396 317902 223448 317908
rect 223580 317960 223632 317966
rect 223580 317902 223632 317908
rect 223304 15088 223356 15094
rect 223304 15030 223356 15036
rect 223408 11490 223436 317902
rect 223488 317620 223540 317626
rect 223488 317562 223540 317568
rect 223396 11484 223448 11490
rect 223396 11426 223448 11432
rect 223500 8226 223528 317562
rect 224052 317558 224080 320076
rect 224420 317626 224448 320076
rect 224788 320062 224894 320090
rect 224408 317620 224460 317626
rect 224408 317562 224460 317568
rect 224040 317552 224092 317558
rect 224040 317494 224092 317500
rect 224684 317552 224736 317558
rect 224684 317494 224736 317500
rect 224696 11558 224724 317494
rect 224684 11552 224736 11558
rect 224684 11494 224736 11500
rect 223488 8220 223540 8226
rect 223488 8162 223540 8168
rect 224788 8090 224816 320062
rect 225340 317966 225368 320076
rect 225814 320062 226104 320090
rect 224868 317960 224920 317966
rect 224868 317902 224920 317908
rect 225328 317960 225380 317966
rect 225328 317902 225380 317908
rect 224880 8158 224908 317902
rect 226076 15026 226104 320062
rect 226156 317960 226208 317966
rect 226156 317902 226208 317908
rect 226064 15020 226116 15026
rect 226064 14962 226116 14968
rect 226168 11626 226196 317902
rect 226156 11620 226208 11626
rect 226156 11562 226208 11568
rect 224868 8152 224920 8158
rect 224868 8094 224920 8100
rect 224776 8084 224828 8090
rect 224776 8026 224828 8032
rect 226260 8022 226288 320076
rect 226720 317966 226748 320076
rect 227194 320062 227484 320090
rect 226708 317960 226760 317966
rect 226708 317902 226760 317908
rect 227456 15774 227484 320062
rect 227536 317960 227588 317966
rect 227536 317902 227588 317908
rect 227444 15768 227496 15774
rect 227444 15710 227496 15716
rect 227548 11694 227576 317902
rect 227536 11688 227588 11694
rect 227536 11630 227588 11636
rect 226248 8016 226300 8022
rect 226248 7958 226300 7964
rect 227640 7954 227668 320076
rect 228008 317966 228036 320076
rect 228482 320062 228864 320090
rect 228942 320062 229048 320090
rect 227996 317960 228048 317966
rect 227996 317902 228048 317908
rect 228836 14958 228864 320062
rect 228916 317960 228968 317966
rect 228916 317902 228968 317908
rect 228824 14952 228876 14958
rect 228824 14894 228876 14900
rect 228928 12442 228956 317902
rect 228916 12436 228968 12442
rect 228916 12378 228968 12384
rect 227628 7948 227680 7954
rect 227628 7890 227680 7896
rect 229020 7886 229048 320062
rect 229388 317626 229416 320076
rect 229376 317620 229428 317626
rect 229376 317562 229428 317568
rect 229848 317558 229876 320076
rect 230204 317620 230256 317626
rect 230204 317562 230256 317568
rect 229836 317552 229888 317558
rect 229836 317494 229888 317500
rect 230216 12374 230244 317562
rect 230204 12368 230256 12374
rect 230204 12310 230256 12316
rect 224132 7880 224184 7886
rect 224132 7822 224184 7828
rect 229008 7880 229060 7886
rect 229008 7822 229060 7828
rect 222936 4616 222988 4622
rect 222936 4558 222988 4564
rect 222108 3460 222160 3466
rect 222108 3402 222160 3408
rect 221738 3360 221794 3369
rect 221738 3295 221794 3304
rect 221752 480 221780 3295
rect 222948 480 222976 4558
rect 224144 480 224172 7822
rect 230308 7818 230336 320076
rect 230768 317626 230796 320076
rect 231242 320062 231624 320090
rect 231702 320062 231808 320090
rect 230756 317620 230808 317626
rect 230756 317562 230808 317568
rect 230388 317552 230440 317558
rect 230388 317494 230440 317500
rect 228916 7812 228968 7818
rect 228916 7754 228968 7760
rect 230296 7812 230348 7818
rect 230296 7754 230348 7760
rect 227720 7744 227772 7750
rect 227720 7686 227772 7692
rect 226524 4684 226576 4690
rect 226524 4626 226576 4632
rect 225328 2984 225380 2990
rect 225328 2926 225380 2932
rect 225340 480 225368 2926
rect 226536 480 226564 4626
rect 227732 480 227760 7686
rect 228928 480 228956 7754
rect 230112 4752 230164 4758
rect 230112 4694 230164 4700
rect 230124 480 230152 4694
rect 230400 4049 230428 317494
rect 231596 14890 231624 320062
rect 231676 317620 231728 317626
rect 231676 317562 231728 317568
rect 231584 14884 231636 14890
rect 231584 14826 231636 14832
rect 231688 12306 231716 317562
rect 231676 12300 231728 12306
rect 231676 12242 231728 12248
rect 231780 7750 231808 320062
rect 232056 317626 232084 320076
rect 232044 317620 232096 317626
rect 232044 317562 232096 317568
rect 232516 317558 232544 320076
rect 232990 320062 233096 320090
rect 232964 317620 233016 317626
rect 232964 317562 233016 317568
rect 232504 317552 232556 317558
rect 232504 317494 232556 317500
rect 232976 12238 233004 317562
rect 232964 12232 233016 12238
rect 232964 12174 233016 12180
rect 231768 7744 231820 7750
rect 231768 7686 231820 7692
rect 233068 7682 233096 320062
rect 233436 317626 233464 320076
rect 234264 318050 234292 320198
rect 234370 320062 234568 320090
rect 234264 318022 234384 318050
rect 233424 317620 233476 317626
rect 233424 317562 233476 317568
rect 233148 317552 233200 317558
rect 233148 317494 233200 317500
rect 232504 7676 232556 7682
rect 232504 7618 232556 7624
rect 233056 7676 233108 7682
rect 233056 7618 233108 7624
rect 231308 7608 231360 7614
rect 231308 7550 231360 7556
rect 230386 4040 230442 4049
rect 230386 3975 230442 3984
rect 231320 480 231348 7550
rect 231766 4584 231822 4593
rect 231766 4519 231822 4528
rect 231780 4185 231808 4519
rect 231766 4176 231822 4185
rect 231766 4111 231822 4120
rect 232516 480 232544 7618
rect 233160 3913 233188 317494
rect 234356 14822 234384 318022
rect 234436 317620 234488 317626
rect 234436 317562 234488 317568
rect 234344 14816 234396 14822
rect 234344 14758 234396 14764
rect 234448 12170 234476 317562
rect 234436 12164 234488 12170
rect 234436 12106 234488 12112
rect 234540 7614 234568 320062
rect 234816 317626 234844 320076
rect 234804 317620 234856 317626
rect 234804 317562 234856 317568
rect 235276 317558 235304 320076
rect 235658 320062 235856 320090
rect 235724 317620 235776 317626
rect 235724 317562 235776 317568
rect 235264 317552 235316 317558
rect 235264 317494 235316 317500
rect 235736 12102 235764 317562
rect 235724 12096 235776 12102
rect 235724 12038 235776 12044
rect 235828 8265 235856 320062
rect 236104 317626 236132 320076
rect 236092 317620 236144 317626
rect 236092 317562 236144 317568
rect 236564 317558 236592 320076
rect 237038 320062 237328 320090
rect 237196 317620 237248 317626
rect 237196 317562 237248 317568
rect 235908 317552 235960 317558
rect 235908 317494 235960 317500
rect 236552 317552 236604 317558
rect 236552 317494 236604 317500
rect 237104 317552 237156 317558
rect 237104 317494 237156 317500
rect 235814 8256 235870 8265
rect 235814 8191 235870 8200
rect 234528 7608 234580 7614
rect 234528 7550 234580 7556
rect 233700 5500 233752 5506
rect 233700 5442 233752 5448
rect 233146 3904 233202 3913
rect 233146 3839 233202 3848
rect 233712 480 233740 5442
rect 234526 4584 234582 4593
rect 234582 4542 234752 4570
rect 234526 4519 234582 4528
rect 234724 4457 234752 4542
rect 234710 4448 234766 4457
rect 234710 4383 234766 4392
rect 235920 3777 235948 317494
rect 237116 14754 237144 317494
rect 237104 14748 237156 14754
rect 237104 14690 237156 14696
rect 237208 12034 237236 317562
rect 237196 12028 237248 12034
rect 237196 11970 237248 11976
rect 237300 8129 237328 320062
rect 237484 317626 237512 320076
rect 237472 317620 237524 317626
rect 237472 317562 237524 317568
rect 237944 317558 237972 320076
rect 238418 320062 238616 320090
rect 238484 317620 238536 317626
rect 238484 317562 238536 317568
rect 237932 317552 237984 317558
rect 237932 317494 237984 317500
rect 238496 11966 238524 317562
rect 238484 11960 238536 11966
rect 238484 11902 238536 11908
rect 237286 8120 237342 8129
rect 237286 8055 237342 8064
rect 238588 7993 238616 320062
rect 238864 317626 238892 320076
rect 238852 317620 238904 317626
rect 238852 317562 238904 317568
rect 239232 317558 239260 320076
rect 239706 320062 240088 320090
rect 239956 317620 240008 317626
rect 239956 317562 240008 317568
rect 238668 317552 238720 317558
rect 238668 317494 238720 317500
rect 239220 317552 239272 317558
rect 239220 317494 239272 317500
rect 239864 317552 239916 317558
rect 239864 317494 239916 317500
rect 238574 7984 238630 7993
rect 238574 7919 238630 7928
rect 237196 5432 237248 5438
rect 237196 5374 237248 5380
rect 235906 3768 235962 3777
rect 235906 3703 235962 3712
rect 234802 3496 234858 3505
rect 234802 3431 234858 3440
rect 234816 480 234844 3431
rect 236000 3120 236052 3126
rect 236000 3062 236052 3068
rect 236012 480 236040 3062
rect 237208 480 237236 5374
rect 238680 3641 238708 317494
rect 239876 14686 239904 317494
rect 239864 14680 239916 14686
rect 239864 14622 239916 14628
rect 239968 11898 239996 317562
rect 239956 11892 240008 11898
rect 239956 11834 240008 11840
rect 240060 7857 240088 320062
rect 240152 317626 240180 320076
rect 240140 317620 240192 317626
rect 240140 317562 240192 317568
rect 240612 317558 240640 320076
rect 241086 320062 241376 320090
rect 241244 317620 241296 317626
rect 241244 317562 241296 317568
rect 240600 317552 240652 317558
rect 240600 317494 240652 317500
rect 241256 11830 241284 317562
rect 241244 11824 241296 11830
rect 241244 11766 241296 11772
rect 240046 7848 240102 7857
rect 240046 7783 240102 7792
rect 241348 7721 241376 320062
rect 241532 317558 241560 320076
rect 241992 317626 242020 320076
rect 242466 320062 242572 320090
rect 241980 317620 242032 317626
rect 241980 317562 242032 317568
rect 241428 317552 241480 317558
rect 241428 317494 241480 317500
rect 241520 317552 241572 317558
rect 241520 317494 241572 317500
rect 241334 7712 241390 7721
rect 241334 7647 241390 7656
rect 240784 5364 240836 5370
rect 240784 5306 240836 5312
rect 238390 3632 238446 3641
rect 238390 3567 238446 3576
rect 238666 3632 238722 3641
rect 238666 3567 238722 3576
rect 238404 480 238432 3567
rect 239588 3052 239640 3058
rect 239588 2994 239640 3000
rect 239600 480 239628 2994
rect 240796 480 240824 5306
rect 241440 3505 241468 317494
rect 242544 15842 242572 320062
rect 242624 317620 242676 317626
rect 242624 317562 242676 317568
rect 242532 15836 242584 15842
rect 242532 15778 242584 15784
rect 242636 14618 242664 317562
rect 242716 317552 242768 317558
rect 242716 317494 242768 317500
rect 242624 14612 242676 14618
rect 242624 14554 242676 14560
rect 242728 11762 242756 317494
rect 242716 11756 242768 11762
rect 242716 11698 242768 11704
rect 241980 8764 242032 8770
rect 241980 8706 242032 8712
rect 241426 3496 241482 3505
rect 241426 3431 241482 3440
rect 241992 480 242020 8706
rect 242820 7585 242848 320076
rect 243280 317626 243308 320076
rect 243754 320062 244044 320090
rect 243268 317620 243320 317626
rect 243268 317562 243320 317568
rect 244016 16590 244044 320062
rect 244108 320062 244214 320090
rect 244004 16584 244056 16590
rect 244004 16526 244056 16532
rect 244108 14550 244136 320062
rect 244188 317620 244240 317626
rect 244188 317562 244240 317568
rect 244096 14544 244148 14550
rect 244096 14486 244148 14492
rect 244200 12209 244228 317562
rect 244660 317558 244688 320076
rect 245134 320062 245424 320090
rect 244648 317552 244700 317558
rect 244648 317494 244700 317500
rect 245396 16522 245424 320062
rect 245488 320062 245594 320090
rect 245384 16516 245436 16522
rect 245384 16458 245436 16464
rect 245488 14482 245516 320062
rect 246040 317626 246068 320076
rect 246514 320062 246804 320090
rect 246304 318708 246356 318714
rect 246304 318650 246356 318656
rect 246028 317620 246080 317626
rect 246028 317562 246080 317568
rect 245568 317552 245620 317558
rect 245568 317494 245620 317500
rect 245476 14476 245528 14482
rect 245476 14418 245528 14424
rect 244186 12200 244242 12209
rect 244186 12135 244242 12144
rect 245580 12073 245608 317494
rect 245566 12064 245622 12073
rect 245566 11999 245622 12008
rect 243176 8900 243228 8906
rect 243176 8842 243228 8848
rect 242806 7576 242862 7585
rect 242806 7511 242862 7520
rect 243188 480 243216 8842
rect 245568 8832 245620 8838
rect 245568 8774 245620 8780
rect 244372 5296 244424 5302
rect 244372 5238 244424 5244
rect 244094 4448 244150 4457
rect 244278 4448 244334 4457
rect 244150 4406 244278 4434
rect 244094 4383 244150 4392
rect 244278 4383 244334 4392
rect 244384 480 244412 5238
rect 245580 480 245608 8774
rect 246316 2922 246344 318650
rect 246776 16386 246804 320062
rect 246868 16454 246896 320076
rect 247328 317626 247356 320076
rect 247802 320062 248184 320090
rect 248262 320062 248368 320090
rect 246948 317620 247000 317626
rect 246948 317562 247000 317568
rect 247316 317620 247368 317626
rect 247316 317562 247368 317568
rect 246856 16448 246908 16454
rect 246856 16390 246908 16396
rect 246764 16380 246816 16386
rect 246764 16322 246816 16328
rect 246960 11937 246988 317562
rect 248156 16318 248184 320062
rect 248236 317620 248288 317626
rect 248236 317562 248288 317568
rect 248144 16312 248196 16318
rect 248144 16254 248196 16260
rect 246946 11928 247002 11937
rect 246946 11863 247002 11872
rect 248248 11801 248276 317562
rect 248234 11792 248290 11801
rect 248234 11727 248290 11736
rect 248340 8702 248368 320062
rect 248708 318170 248736 320076
rect 249182 320062 249564 320090
rect 249642 320062 249748 320090
rect 248696 318164 248748 318170
rect 248696 318106 248748 318112
rect 249536 16250 249564 320062
rect 249616 318164 249668 318170
rect 249616 318106 249668 318112
rect 249524 16244 249576 16250
rect 249524 16186 249576 16192
rect 249628 11665 249656 318106
rect 249614 11656 249670 11665
rect 249614 11591 249670 11600
rect 249156 9648 249208 9654
rect 249156 9590 249208 9596
rect 248328 8696 248380 8702
rect 248328 8638 248380 8644
rect 247960 5228 248012 5234
rect 247960 5170 248012 5176
rect 246764 3188 246816 3194
rect 246764 3130 246816 3136
rect 246304 2916 246356 2922
rect 246304 2858 246356 2864
rect 246776 480 246804 3130
rect 247972 480 248000 5170
rect 249168 480 249196 9590
rect 249720 8770 249748 320062
rect 250088 318170 250116 320076
rect 250076 318164 250128 318170
rect 250076 318106 250128 318112
rect 250824 318050 250852 320198
rect 250930 320062 251128 320090
rect 250996 318164 251048 318170
rect 250996 318106 251048 318112
rect 250824 318022 250944 318050
rect 250444 317824 250496 317830
rect 250444 317766 250496 317772
rect 250352 9580 250404 9586
rect 250352 9522 250404 9528
rect 249708 8764 249760 8770
rect 249708 8706 249760 8712
rect 250364 480 250392 9522
rect 250456 3058 250484 317766
rect 250916 16182 250944 318022
rect 250904 16176 250956 16182
rect 250904 16118 250956 16124
rect 251008 15065 251036 318106
rect 250994 15056 251050 15065
rect 250994 14991 251050 15000
rect 251100 8838 251128 320062
rect 251376 318170 251404 320076
rect 251850 320062 252140 320090
rect 252310 320062 252508 320090
rect 251364 318164 251416 318170
rect 251364 318106 251416 318112
rect 252112 318050 252140 320062
rect 252376 318164 252428 318170
rect 252376 318106 252428 318112
rect 252112 318022 252324 318050
rect 252296 16114 252324 318022
rect 252284 16108 252336 16114
rect 252284 16050 252336 16056
rect 252388 14929 252416 318106
rect 252374 14920 252430 14929
rect 252374 14855 252430 14864
rect 252480 8906 252508 320062
rect 252756 318170 252784 320076
rect 252744 318164 252796 318170
rect 252744 318106 252796 318112
rect 253216 317898 253244 320076
rect 253690 320062 253796 320090
rect 253664 318164 253716 318170
rect 253664 318106 253716 318112
rect 253112 317892 253164 317898
rect 253112 317834 253164 317840
rect 253204 317892 253256 317898
rect 253204 317834 253256 317840
rect 253124 317778 253152 317834
rect 253124 317750 253244 317778
rect 252652 9512 252704 9518
rect 252652 9454 252704 9460
rect 252468 8900 252520 8906
rect 252468 8842 252520 8848
rect 251088 8832 251140 8838
rect 251088 8774 251140 8780
rect 251456 5160 251508 5166
rect 251456 5102 251508 5108
rect 250444 3052 250496 3058
rect 250444 2994 250496 3000
rect 251468 480 251496 5102
rect 252664 480 252692 9454
rect 253216 3194 253244 317750
rect 253296 317756 253348 317762
rect 253296 317698 253348 317704
rect 253204 3188 253256 3194
rect 253204 3130 253256 3136
rect 253308 2990 253336 317698
rect 253676 14793 253704 318106
rect 253662 14784 253718 14793
rect 253662 14719 253718 14728
rect 253768 9654 253796 320062
rect 254044 318170 254072 320076
rect 254032 318164 254084 318170
rect 254032 318106 254084 318112
rect 254504 317898 254532 320076
rect 254978 320062 255176 320090
rect 255044 318164 255096 318170
rect 255044 318106 255096 318112
rect 253848 317892 253900 317898
rect 253848 317834 253900 317840
rect 254492 317892 254544 317898
rect 254492 317834 254544 317840
rect 253756 9648 253808 9654
rect 253756 9590 253808 9596
rect 253860 4418 253888 317834
rect 255056 14657 255084 318106
rect 255042 14648 255098 14657
rect 255042 14583 255098 14592
rect 255148 9586 255176 320062
rect 255424 318170 255452 320076
rect 255412 318164 255464 318170
rect 255412 318106 255464 318112
rect 255884 317898 255912 320076
rect 256358 320062 256556 320090
rect 256424 318164 256476 318170
rect 256424 318106 256476 318112
rect 255228 317892 255280 317898
rect 255228 317834 255280 317840
rect 255872 317892 255924 317898
rect 255872 317834 255924 317840
rect 255136 9580 255188 9586
rect 255136 9522 255188 9528
rect 255044 5092 255096 5098
rect 255044 5034 255096 5040
rect 253848 4412 253900 4418
rect 253848 4354 253900 4360
rect 253848 3256 253900 3262
rect 253848 3198 253900 3204
rect 253296 2984 253348 2990
rect 253296 2926 253348 2932
rect 253860 480 253888 3198
rect 255056 480 255084 5034
rect 255240 4486 255268 317834
rect 255964 317620 256016 317626
rect 255964 317562 256016 317568
rect 255228 4480 255280 4486
rect 255228 4422 255280 4428
rect 255976 3262 256004 317562
rect 256436 13598 256464 318106
rect 256424 13592 256476 13598
rect 256424 13534 256476 13540
rect 256528 9518 256556 320062
rect 256804 318170 256832 320076
rect 256792 318164 256844 318170
rect 256792 318106 256844 318112
rect 257264 317898 257292 320076
rect 257738 320062 257936 320090
rect 257804 318164 257856 318170
rect 257804 318106 257856 318112
rect 256608 317892 256660 317898
rect 256608 317834 256660 317840
rect 257252 317892 257304 317898
rect 257252 317834 257304 317840
rect 256516 9512 256568 9518
rect 256516 9454 256568 9460
rect 256240 9444 256292 9450
rect 256240 9386 256292 9392
rect 255964 3256 256016 3262
rect 255964 3198 256016 3204
rect 256252 480 256280 9386
rect 256620 4554 256648 317834
rect 257816 13530 257844 318106
rect 257804 13524 257856 13530
rect 257804 13466 257856 13472
rect 257908 9450 257936 320062
rect 258092 318170 258120 320076
rect 258080 318164 258132 318170
rect 258080 318106 258132 318112
rect 258552 317898 258580 320076
rect 259026 320062 259316 320090
rect 259184 318164 259236 318170
rect 259184 318106 259236 318112
rect 257988 317892 258040 317898
rect 257988 317834 258040 317840
rect 258540 317892 258592 317898
rect 258540 317834 258592 317840
rect 257896 9444 257948 9450
rect 257896 9386 257948 9392
rect 257436 9376 257488 9382
rect 257436 9318 257488 9324
rect 256608 4548 256660 4554
rect 256608 4490 256660 4496
rect 257448 480 257476 9318
rect 258000 4622 258028 317834
rect 259196 13462 259224 318106
rect 259184 13456 259236 13462
rect 259184 13398 259236 13404
rect 259288 9382 259316 320062
rect 259368 317892 259420 317898
rect 259368 317834 259420 317840
rect 259276 9376 259328 9382
rect 259276 9318 259328 9324
rect 258632 5024 258684 5030
rect 258632 4966 258684 4972
rect 257988 4616 258040 4622
rect 257988 4558 258040 4564
rect 258644 480 258672 4966
rect 259380 4690 259408 317834
rect 259472 317558 259500 320076
rect 259932 318170 259960 320076
rect 260406 320062 260696 320090
rect 259920 318164 259972 318170
rect 259920 318106 259972 318112
rect 259460 317552 259512 317558
rect 259460 317494 259512 317500
rect 260564 317552 260616 317558
rect 260564 317494 260616 317500
rect 260576 13394 260604 317494
rect 260564 13388 260616 13394
rect 260564 13330 260616 13336
rect 260668 9625 260696 320062
rect 260748 318164 260800 318170
rect 260748 318106 260800 318112
rect 260654 9616 260710 9625
rect 260654 9551 260710 9560
rect 259828 6248 259880 6254
rect 259828 6190 259880 6196
rect 259368 4684 259420 4690
rect 259368 4626 259420 4632
rect 259366 4584 259422 4593
rect 259366 4519 259422 4528
rect 259380 4321 259408 4519
rect 259366 4312 259422 4321
rect 259366 4247 259422 4256
rect 259840 480 259868 6190
rect 260760 4758 260788 318106
rect 260852 317898 260880 320076
rect 260840 317892 260892 317898
rect 260840 317834 260892 317840
rect 261312 317830 261340 320076
rect 261694 320062 262076 320090
rect 261852 318164 261904 318170
rect 261852 318106 261904 318112
rect 261300 317824 261352 317830
rect 261300 317766 261352 317772
rect 261864 13258 261892 318106
rect 261944 317892 261996 317898
rect 261944 317834 261996 317840
rect 261956 13326 261984 317834
rect 261944 13320 261996 13326
rect 261944 13262 261996 13268
rect 261852 13252 261904 13258
rect 261852 13194 261904 13200
rect 262048 9314 262076 320062
rect 262140 318170 262168 320076
rect 262128 318164 262180 318170
rect 262128 318106 262180 318112
rect 262128 317824 262180 317830
rect 262128 317766 262180 317772
rect 261024 9308 261076 9314
rect 261024 9250 261076 9256
rect 262036 9308 262088 9314
rect 262036 9250 262088 9256
rect 260748 4752 260800 4758
rect 260748 4694 260800 4700
rect 261036 480 261064 9250
rect 262140 5506 262168 317766
rect 262600 317762 262628 320076
rect 263074 320062 263456 320090
rect 263324 318164 263376 318170
rect 263324 318106 263376 318112
rect 262588 317756 262640 317762
rect 262588 317698 262640 317704
rect 263336 13190 263364 318106
rect 263324 13184 263376 13190
rect 263324 13126 263376 13132
rect 263428 9489 263456 320062
rect 263520 318170 263548 320076
rect 263508 318164 263560 318170
rect 263508 318106 263560 318112
rect 263980 317898 264008 320076
rect 264454 320062 264836 320090
rect 264704 318164 264756 318170
rect 264704 318106 264756 318112
rect 263968 317892 264020 317898
rect 263968 317834 264020 317840
rect 263508 317756 263560 317762
rect 263508 317698 263560 317704
rect 263414 9480 263470 9489
rect 263414 9415 263470 9424
rect 263416 6180 263468 6186
rect 263416 6122 263468 6128
rect 262128 5500 262180 5506
rect 262128 5442 262180 5448
rect 262220 4956 262272 4962
rect 262220 4898 262272 4904
rect 262232 480 262260 4898
rect 263428 480 263456 6122
rect 263520 5438 263548 317698
rect 264716 13122 264744 318106
rect 264704 13116 264756 13122
rect 264704 13058 264756 13064
rect 264808 9246 264836 320062
rect 264900 318170 264928 320076
rect 265268 318170 265296 320076
rect 265742 320062 266124 320090
rect 264888 318164 264940 318170
rect 264888 318106 264940 318112
rect 265256 318164 265308 318170
rect 265256 318106 265308 318112
rect 264888 317892 264940 317898
rect 264888 317834 264940 317840
rect 264612 9240 264664 9246
rect 264612 9182 264664 9188
rect 264796 9240 264848 9246
rect 264796 9182 264848 9188
rect 263508 5432 263560 5438
rect 263508 5374 263560 5380
rect 264624 480 264652 9182
rect 264900 5370 264928 317834
rect 266096 14521 266124 320062
rect 266082 14512 266138 14521
rect 266082 14447 266138 14456
rect 266188 13569 266216 320076
rect 266268 318164 266320 318170
rect 266268 318106 266320 318112
rect 266174 13560 266230 13569
rect 266174 13495 266230 13504
rect 264888 5364 264940 5370
rect 264888 5306 264940 5312
rect 266280 5302 266308 318106
rect 266648 317898 266676 320076
rect 267108 318170 267136 320076
rect 267476 320062 267582 320090
rect 267096 318164 267148 318170
rect 267096 318106 267148 318112
rect 266636 317892 266688 317898
rect 266636 317834 266688 317840
rect 267476 13433 267504 320062
rect 268028 318170 268056 320076
rect 267556 318164 267608 318170
rect 267556 318106 267608 318112
rect 268016 318164 268068 318170
rect 268016 318106 268068 318112
rect 267462 13424 267518 13433
rect 267462 13359 267518 13368
rect 267568 9353 267596 318106
rect 268488 318102 268516 320076
rect 268856 320062 268962 320090
rect 268476 318096 268528 318102
rect 268476 318038 268528 318044
rect 267648 317892 267700 317898
rect 267648 317834 267700 317840
rect 267554 9344 267610 9353
rect 267554 9279 267610 9288
rect 267004 6996 267056 7002
rect 267004 6938 267056 6944
rect 266268 5296 266320 5302
rect 266268 5238 266320 5244
rect 265808 4888 265860 4894
rect 265808 4830 265860 4836
rect 265820 480 265848 4830
rect 267016 480 267044 6938
rect 267660 5234 267688 317834
rect 268856 13297 268884 320062
rect 269316 318170 269344 320076
rect 269028 318164 269080 318170
rect 269028 318106 269080 318112
rect 269304 318164 269356 318170
rect 269304 318106 269356 318112
rect 268936 318096 268988 318102
rect 268936 318038 268988 318044
rect 268842 13288 268898 13297
rect 268842 13223 268898 13232
rect 268948 9178 268976 318038
rect 268108 9172 268160 9178
rect 268108 9114 268160 9120
rect 268936 9172 268988 9178
rect 268936 9114 268988 9120
rect 267648 5228 267700 5234
rect 267648 5170 267700 5176
rect 268120 480 268148 9114
rect 269040 5166 269068 318106
rect 269776 318102 269804 320076
rect 269764 318096 269816 318102
rect 269764 318038 269816 318044
rect 270236 13161 270264 320076
rect 270696 318170 270724 320076
rect 270408 318164 270460 318170
rect 270408 318106 270460 318112
rect 270684 318164 270736 318170
rect 270684 318106 270736 318112
rect 270316 318096 270368 318102
rect 270316 318038 270368 318044
rect 270222 13152 270278 13161
rect 270222 13087 270278 13096
rect 270328 9217 270356 318038
rect 270314 9208 270370 9217
rect 270314 9143 270370 9152
rect 269028 5160 269080 5166
rect 269028 5102 269080 5108
rect 270420 5098 270448 318106
rect 271156 318102 271184 320076
rect 271144 318096 271196 318102
rect 271144 318038 271196 318044
rect 271144 317892 271196 317898
rect 271144 317834 271196 317840
rect 270500 9104 270552 9110
rect 270500 9046 270552 9052
rect 270408 5092 270460 5098
rect 270408 5034 270460 5040
rect 269304 4820 269356 4826
rect 269304 4762 269356 4768
rect 269316 480 269344 4762
rect 270512 480 270540 9046
rect 271156 2854 271184 317834
rect 271236 317688 271288 317694
rect 271236 317630 271288 317636
rect 271248 3126 271276 317630
rect 271616 13025 271644 320076
rect 271788 318164 271840 318170
rect 271788 318106 271840 318112
rect 271696 318096 271748 318102
rect 271696 318038 271748 318044
rect 271602 13016 271658 13025
rect 271602 12951 271658 12960
rect 271708 9110 271736 318038
rect 271696 9104 271748 9110
rect 271696 9046 271748 9052
rect 271800 5030 271828 318106
rect 272076 318102 272104 320076
rect 272536 318170 272564 320076
rect 272904 318510 272932 320076
rect 272892 318504 272944 318510
rect 272892 318446 272944 318452
rect 273364 318170 273392 320076
rect 272524 318164 272576 318170
rect 272524 318106 272576 318112
rect 273076 318164 273128 318170
rect 273076 318106 273128 318112
rect 273352 318164 273404 318170
rect 273352 318106 273404 318112
rect 272064 318096 272116 318102
rect 272064 318038 272116 318044
rect 273088 6254 273116 318106
rect 273824 318102 273852 320076
rect 274298 320062 274404 320090
rect 273168 318096 273220 318102
rect 273168 318038 273220 318044
rect 273812 318096 273864 318102
rect 273812 318038 273864 318044
rect 273076 6248 273128 6254
rect 273076 6190 273128 6196
rect 272890 5128 272946 5137
rect 272890 5063 272946 5072
rect 271788 5024 271840 5030
rect 271788 4966 271840 4972
rect 271696 3392 271748 3398
rect 271696 3334 271748 3340
rect 271236 3120 271288 3126
rect 271236 3062 271288 3068
rect 271144 2848 271196 2854
rect 271144 2790 271196 2796
rect 271708 480 271736 3334
rect 272904 480 272932 5063
rect 273180 4962 273208 318038
rect 274376 16046 274404 320062
rect 274548 318164 274600 318170
rect 274548 318106 274600 318112
rect 274456 318096 274508 318102
rect 274456 318038 274508 318044
rect 274364 16040 274416 16046
rect 274364 15982 274416 15988
rect 274468 9042 274496 318038
rect 274088 9036 274140 9042
rect 274088 8978 274140 8984
rect 274456 9036 274508 9042
rect 274456 8978 274508 8984
rect 273168 4956 273220 4962
rect 273168 4898 273220 4904
rect 273442 4312 273498 4321
rect 273442 4247 273498 4256
rect 273456 2378 273484 4247
rect 273444 2372 273496 2378
rect 273444 2314 273496 2320
rect 274100 480 274128 8978
rect 274560 4894 274588 318106
rect 274744 318102 274772 320076
rect 274732 318096 274784 318102
rect 274732 318038 274784 318044
rect 275204 317830 275232 320076
rect 275664 318170 275692 320076
rect 275652 318164 275704 318170
rect 275652 318106 275704 318112
rect 275928 318096 275980 318102
rect 275928 318038 275980 318044
rect 275284 317892 275336 317898
rect 275284 317834 275336 317840
rect 275192 317824 275244 317830
rect 275192 317766 275244 317772
rect 274548 4888 274600 4894
rect 274548 4830 274600 4836
rect 275296 3398 275324 317834
rect 275836 317824 275888 317830
rect 275836 317766 275888 317772
rect 275848 9081 275876 317766
rect 275834 9072 275890 9081
rect 275834 9007 275890 9016
rect 275940 4826 275968 318038
rect 276124 317898 276152 320076
rect 276492 318102 276520 320076
rect 276966 320062 277164 320090
rect 276480 318096 276532 318102
rect 276480 318038 276532 318044
rect 276112 317892 276164 317898
rect 276112 317834 276164 317840
rect 277136 15978 277164 320062
rect 277216 318096 277268 318102
rect 277216 318038 277268 318044
rect 277124 15972 277176 15978
rect 277124 15914 277176 15920
rect 277228 6186 277256 318038
rect 277308 317892 277360 317898
rect 277308 317834 277360 317840
rect 277216 6180 277268 6186
rect 277216 6122 277268 6128
rect 277320 5137 277348 317834
rect 277412 317830 277440 320076
rect 277872 317898 277900 320076
rect 278346 320062 278544 320090
rect 277860 317892 277912 317898
rect 277860 317834 277912 317840
rect 277400 317824 277452 317830
rect 277400 317766 277452 317772
rect 278516 15910 278544 320062
rect 278792 317898 278820 320076
rect 279266 320062 279648 320090
rect 279424 318436 279476 318442
rect 279424 318378 279476 318384
rect 278596 317892 278648 317898
rect 278596 317834 278648 317840
rect 278780 317892 278832 317898
rect 278780 317834 278832 317840
rect 278504 15904 278556 15910
rect 278504 15846 278556 15852
rect 278608 8974 278636 317834
rect 278688 317824 278740 317830
rect 278688 317766 278740 317772
rect 277676 8968 277728 8974
rect 277676 8910 277728 8916
rect 278596 8968 278648 8974
rect 278596 8910 278648 8916
rect 277306 5128 277362 5137
rect 277306 5063 277362 5072
rect 276478 4992 276534 5001
rect 276478 4927 276534 4936
rect 275928 4820 275980 4826
rect 275928 4762 275980 4768
rect 275284 3392 275336 3398
rect 275284 3334 275336 3340
rect 275284 2916 275336 2922
rect 275284 2858 275336 2864
rect 275296 480 275324 2858
rect 276492 480 276520 4927
rect 277688 480 277716 8910
rect 278700 5001 278728 317766
rect 278686 4992 278742 5001
rect 278686 4927 278742 4936
rect 278872 2984 278924 2990
rect 278872 2926 278924 2932
rect 278884 480 278912 2926
rect 279436 2854 279464 318378
rect 279620 318050 279648 320062
rect 279712 318345 279740 320076
rect 405016 318782 405044 412626
rect 438136 410854 438164 646031
rect 438214 645008 438270 645017
rect 438214 644943 438270 644952
rect 438124 410848 438176 410854
rect 438124 410790 438176 410796
rect 438228 410786 438256 644943
rect 438306 643240 438362 643249
rect 438306 643175 438362 643184
rect 438216 410780 438268 410786
rect 438216 410722 438268 410728
rect 438320 410718 438348 643175
rect 438398 642016 438454 642025
rect 438398 641951 438454 641960
rect 438308 410712 438360 410718
rect 438308 410654 438360 410660
rect 438412 410582 438440 641951
rect 438490 640384 438546 640393
rect 438490 640319 438546 640328
rect 438504 412146 438532 640319
rect 438582 639296 438638 639305
rect 438582 639231 438638 639240
rect 438596 412214 438624 639231
rect 438674 637664 438730 637673
rect 438674 637599 438730 637608
rect 438584 412208 438636 412214
rect 438584 412150 438636 412156
rect 438492 412140 438544 412146
rect 438492 412082 438544 412088
rect 438688 412078 438716 637599
rect 518912 589393 518940 652734
rect 518898 589384 518954 589393
rect 518898 589319 518954 589328
rect 518912 587761 518940 589319
rect 518898 587752 518954 587761
rect 518898 587687 518954 587696
rect 438766 579728 438822 579737
rect 438766 579663 438822 579672
rect 438676 412072 438728 412078
rect 438676 412014 438728 412020
rect 438780 410650 438808 579663
rect 443090 558920 443146 558929
rect 443090 558855 443146 558864
rect 445758 558920 445814 558929
rect 447598 558920 447654 558929
rect 445758 558855 445814 558864
rect 446404 558884 446456 558890
rect 441620 558816 441672 558822
rect 441620 558758 441672 558764
rect 441632 557598 441660 558758
rect 443104 558550 443132 558855
rect 443092 558544 443144 558550
rect 443092 558486 443144 558492
rect 443644 558000 443696 558006
rect 443644 557942 443696 557948
rect 441620 557592 441672 557598
rect 441620 557534 441672 557540
rect 443656 522986 443684 557942
rect 443644 522980 443696 522986
rect 443644 522922 443696 522928
rect 445772 412010 445800 558855
rect 447598 558855 447654 558864
rect 453670 558920 453726 558929
rect 453670 558855 453726 558864
rect 454682 558920 454738 558929
rect 454682 558855 454738 558864
rect 455970 558920 456026 558929
rect 455970 558855 456026 558864
rect 457350 558920 457406 558929
rect 457350 558855 457406 558864
rect 458270 558920 458326 558929
rect 458270 558855 458326 558864
rect 460846 558920 460902 558929
rect 460846 558855 460902 558864
rect 461674 558920 461730 558929
rect 461674 558855 461730 558864
rect 462594 558920 462650 558929
rect 462594 558855 462650 558864
rect 464250 558920 464306 558929
rect 464250 558855 464306 558864
rect 465262 558920 465318 558929
rect 465262 558855 465318 558864
rect 466458 558920 466514 558929
rect 466458 558855 466514 558864
rect 467838 558920 467894 558929
rect 467838 558855 467894 558864
rect 468666 558920 468722 558929
rect 468666 558855 468722 558864
rect 469218 558920 469274 558929
rect 469218 558855 469274 558864
rect 470598 558920 470654 558929
rect 470598 558855 470654 558864
rect 471978 558920 472034 558929
rect 471978 558855 472034 558864
rect 473358 558920 473414 558929
rect 473358 558855 473414 558864
rect 474830 558920 474886 558929
rect 474830 558855 474886 558864
rect 475474 558920 475530 558929
rect 475474 558855 475530 558864
rect 477130 558920 477186 558929
rect 477130 558855 477186 558864
rect 478234 558920 478290 558929
rect 478234 558855 478290 558864
rect 478970 558920 479026 558929
rect 478970 558855 479026 558864
rect 480534 558920 480590 558929
rect 480534 558855 480536 558864
rect 446404 558826 446456 558832
rect 446416 525774 446444 558826
rect 447612 558210 447640 558855
rect 452658 558784 452714 558793
rect 453684 558754 453712 558855
rect 452658 558719 452714 558728
rect 453672 558748 453724 558754
rect 451740 558544 451792 558550
rect 449898 558512 449954 558521
rect 452384 558544 452436 558550
rect 451792 558492 452384 558498
rect 451740 558486 452436 558492
rect 451752 558470 452424 558486
rect 452672 558482 452700 558719
rect 453672 558690 453724 558696
rect 454696 558686 454724 558855
rect 454040 558680 454092 558686
rect 453302 558648 453358 558657
rect 453302 558583 453358 558592
rect 453946 558648 454002 558657
rect 454040 558622 454092 558628
rect 454684 558680 454736 558686
rect 454684 558622 454736 558628
rect 453946 558583 454002 558592
rect 452660 558476 452712 558482
rect 449898 558447 449954 558456
rect 447600 558204 447652 558210
rect 447600 558146 447652 558152
rect 449912 558142 449940 558447
rect 452660 558418 452712 558424
rect 449900 558136 449952 558142
rect 449900 558078 449952 558084
rect 451278 558104 451334 558113
rect 451278 558039 451280 558048
rect 451332 558039 451334 558048
rect 451280 558010 451332 558016
rect 449164 557932 449216 557938
rect 449164 557874 449216 557880
rect 447784 557864 447836 557870
rect 447784 557806 447836 557812
rect 447796 527134 447824 557806
rect 449176 529922 449204 557874
rect 451924 557796 451976 557802
rect 451924 557738 451976 557744
rect 450544 557728 450596 557734
rect 450544 557670 450596 557676
rect 450556 531282 450584 557670
rect 451936 534070 451964 557738
rect 452658 557560 452714 557569
rect 452658 557495 452714 557504
rect 451924 534064 451976 534070
rect 451924 534006 451976 534012
rect 450544 531276 450596 531282
rect 450544 531218 450596 531224
rect 449164 529916 449216 529922
rect 449164 529858 449216 529864
rect 447784 527128 447836 527134
rect 447784 527070 447836 527076
rect 446404 525768 446456 525774
rect 446404 525710 446456 525716
rect 452672 476066 452700 557495
rect 452660 476060 452712 476066
rect 452660 476002 452712 476008
rect 445760 412004 445812 412010
rect 445760 411946 445812 411952
rect 453316 411942 453344 558583
rect 453960 558550 453988 558583
rect 453948 558544 454000 558550
rect 453948 558486 454000 558492
rect 453488 557660 453540 557666
rect 453488 557602 453540 557608
rect 453394 557560 453450 557569
rect 453394 557495 453450 557504
rect 453408 480214 453436 557495
rect 453500 535430 453528 557602
rect 454052 557598 454080 558622
rect 455984 558618 456012 558855
rect 457364 558822 457392 558855
rect 457352 558816 457404 558822
rect 457352 558758 457404 558764
rect 455972 558612 456024 558618
rect 455972 558554 456024 558560
rect 458284 558006 458312 558855
rect 459650 558648 459706 558657
rect 459650 558583 459706 558592
rect 459468 558476 459520 558482
rect 459468 558418 459520 558424
rect 459480 558006 459508 558418
rect 458272 558000 458324 558006
rect 458272 557942 458324 557948
rect 459468 558000 459520 558006
rect 459468 557942 459520 557948
rect 454684 557932 454736 557938
rect 454684 557874 454736 557880
rect 454040 557592 454092 557598
rect 454040 557534 454092 557540
rect 454696 538218 454724 557874
rect 459664 557598 459692 558583
rect 460860 558006 460888 558855
rect 461688 558550 461716 558855
rect 462608 558754 462636 558855
rect 462596 558748 462648 558754
rect 462596 558690 462648 558696
rect 462962 558648 463018 558657
rect 462962 558583 462964 558592
rect 463016 558583 463018 558592
rect 462964 558554 463016 558560
rect 461676 558544 461728 558550
rect 461676 558486 461728 558492
rect 460848 558000 460900 558006
rect 460848 557942 460900 557948
rect 461030 557696 461086 557705
rect 461030 557631 461086 557640
rect 459652 557592 459704 557598
rect 455418 557560 455474 557569
rect 455418 557495 455474 557504
rect 456798 557560 456854 557569
rect 456798 557495 456854 557504
rect 458178 557560 458234 557569
rect 458178 557495 458234 557504
rect 459558 557560 459614 557569
rect 459652 557534 459704 557540
rect 460938 557560 460994 557569
rect 459558 557495 459614 557504
rect 460938 557495 460994 557504
rect 454684 538212 454736 538218
rect 454684 538154 454736 538160
rect 453488 535424 453540 535430
rect 453488 535366 453540 535372
rect 455432 483002 455460 557495
rect 456812 484362 456840 557495
rect 458192 487150 458220 557495
rect 459572 488510 459600 557495
rect 460952 491298 460980 557495
rect 461044 492658 461072 557631
rect 464264 557598 464292 558855
rect 465276 558686 465304 558855
rect 465264 558680 465316 558686
rect 465264 558622 465316 558628
rect 464344 557932 464396 557938
rect 464344 557874 464396 557880
rect 464252 557592 464304 557598
rect 462318 557560 462374 557569
rect 462318 557495 462374 557504
rect 463698 557560 463754 557569
rect 464252 557534 464304 557540
rect 463698 557495 463754 557504
rect 462332 495446 462360 557495
rect 463712 496806 463740 557495
rect 464356 539578 464384 557874
rect 465078 557560 465134 557569
rect 465078 557495 465134 557504
rect 464344 539572 464396 539578
rect 464344 539514 464396 539520
rect 465092 499526 465120 557495
rect 466472 500954 466500 558855
rect 466552 558816 466604 558822
rect 466550 558784 466552 558793
rect 466604 558784 466606 558793
rect 466550 558719 466606 558728
rect 467852 502314 467880 558855
rect 467930 558784 467986 558793
rect 467930 558719 467986 558728
rect 467944 505102 467972 558719
rect 468022 558648 468078 558657
rect 468680 558618 468708 558855
rect 468022 558583 468078 558592
rect 468668 558612 468720 558618
rect 468036 558482 468064 558583
rect 468668 558554 468720 558560
rect 468024 558476 468076 558482
rect 468024 558418 468076 558424
rect 468760 558476 468812 558482
rect 468760 558418 468812 558424
rect 468772 558006 468800 558418
rect 468760 558000 468812 558006
rect 468760 557942 468812 557948
rect 469232 506462 469260 558855
rect 470046 558784 470102 558793
rect 470046 558719 470102 558728
rect 470060 558482 470088 558719
rect 470048 558476 470100 558482
rect 470048 558418 470100 558424
rect 470612 509250 470640 558855
rect 471334 558784 471390 558793
rect 471334 558719 471390 558728
rect 471348 558550 471376 558719
rect 471336 558544 471388 558550
rect 471336 558486 471388 558492
rect 471992 510610 472020 558855
rect 472162 558784 472218 558793
rect 472162 558719 472164 558728
rect 472216 558719 472218 558728
rect 472164 558690 472216 558696
rect 473372 513330 473400 558855
rect 474844 558686 474872 558855
rect 475488 558822 475516 558855
rect 475476 558816 475528 558822
rect 475476 558758 475528 558764
rect 474832 558680 474884 558686
rect 473450 558648 473506 558657
rect 474832 558622 474884 558628
rect 475488 558618 475516 558758
rect 473450 558583 473506 558592
rect 475476 558612 475528 558618
rect 473464 557598 473492 558583
rect 475476 558554 475528 558560
rect 476118 558512 476174 558521
rect 476118 558447 476174 558456
rect 476132 558414 476160 558447
rect 477144 558414 477172 558855
rect 477592 558476 477644 558482
rect 477592 558418 477644 558424
rect 476120 558408 476172 558414
rect 476304 558408 476356 558414
rect 476120 558350 476172 558356
rect 476210 558376 476266 558385
rect 476304 558350 476356 558356
rect 477132 558408 477184 558414
rect 477132 558350 477184 558356
rect 477498 558376 477554 558385
rect 476210 558311 476266 558320
rect 476224 558278 476252 558311
rect 476212 558272 476264 558278
rect 476212 558214 476264 558220
rect 476316 557598 476344 558350
rect 477498 558311 477500 558320
rect 477552 558311 477554 558320
rect 477500 558282 477552 558288
rect 477604 558278 477632 558418
rect 478248 558278 478276 558855
rect 477592 558272 477644 558278
rect 477592 558214 477644 558220
rect 478236 558272 478288 558278
rect 478236 558214 478288 558220
rect 478878 558240 478934 558249
rect 478984 558210 479012 558855
rect 480588 558855 480590 558864
rect 483018 558920 483074 558929
rect 483018 558855 483074 558864
rect 480536 558826 480588 558832
rect 483032 558822 483060 558855
rect 483020 558816 483072 558822
rect 480350 558784 480406 558793
rect 480350 558719 480406 558728
rect 481638 558784 481694 558793
rect 483020 558758 483072 558764
rect 481638 558719 481640 558728
rect 480364 558550 480392 558719
rect 481692 558719 481694 558728
rect 481640 558690 481692 558696
rect 484398 558648 484454 558657
rect 484398 558583 484400 558592
rect 484452 558583 484454 558592
rect 488538 558648 488594 558657
rect 488538 558583 488594 558592
rect 484400 558554 484452 558560
rect 480352 558544 480404 558550
rect 480352 558486 480404 558492
rect 481638 558512 481694 558521
rect 481638 558447 481694 558456
rect 485778 558512 485834 558521
rect 485778 558447 485834 558456
rect 487158 558512 487214 558521
rect 487158 558447 487214 558456
rect 478878 558175 478880 558184
rect 478932 558175 478934 558184
rect 478972 558204 479024 558210
rect 478880 558146 478932 558152
rect 478972 558146 479024 558152
rect 478984 558006 479012 558146
rect 481652 558074 481680 558447
rect 485792 558414 485820 558447
rect 485780 558408 485832 558414
rect 485780 558350 485832 558356
rect 487172 558278 487200 558447
rect 487160 558272 487212 558278
rect 483018 558240 483074 558249
rect 483018 558175 483074 558184
rect 484398 558240 484454 558249
rect 484398 558175 484454 558184
rect 485778 558240 485834 558249
rect 487160 558214 487212 558220
rect 488552 558210 488580 558583
rect 485778 558175 485834 558184
rect 488540 558204 488592 558210
rect 483032 558142 483060 558175
rect 483020 558136 483072 558142
rect 483020 558078 483072 558084
rect 483110 558104 483166 558113
rect 481640 558068 481692 558074
rect 483110 558039 483166 558048
rect 481640 558010 481692 558016
rect 478972 558000 479024 558006
rect 478972 557942 479024 557948
rect 483124 557734 483152 558039
rect 484412 557802 484440 558175
rect 484400 557796 484452 557802
rect 484400 557738 484452 557744
rect 483112 557728 483164 557734
rect 483018 557696 483074 557705
rect 483112 557670 483164 557676
rect 485792 557666 485820 558175
rect 488540 558146 488592 558152
rect 488538 558104 488594 558113
rect 488538 558039 488594 558048
rect 487158 557968 487214 557977
rect 488552 557938 488580 558039
rect 487158 557903 487214 557912
rect 488540 557932 488592 557938
rect 487172 557870 487200 557903
rect 488540 557874 488592 557880
rect 487160 557864 487212 557870
rect 487160 557806 487212 557812
rect 483018 557631 483074 557640
rect 485780 557660 485832 557666
rect 483032 557598 483060 557631
rect 485780 557602 485832 557608
rect 473452 557592 473504 557598
rect 474648 557592 474700 557598
rect 473452 557534 473504 557540
rect 474646 557560 474648 557569
rect 476304 557592 476356 557598
rect 474700 557560 474702 557569
rect 476396 557592 476448 557598
rect 476304 557534 476356 557540
rect 476394 557560 476396 557569
rect 483020 557592 483072 557598
rect 476448 557560 476450 557569
rect 474646 557495 474702 557504
rect 483020 557534 483072 557540
rect 476394 557495 476450 557504
rect 473360 513324 473412 513330
rect 473360 513266 473412 513272
rect 471980 510604 472032 510610
rect 471980 510546 472032 510552
rect 470600 509244 470652 509250
rect 470600 509186 470652 509192
rect 469220 506456 469272 506462
rect 469220 506398 469272 506404
rect 467932 505096 467984 505102
rect 467932 505038 467984 505044
rect 467840 502308 467892 502314
rect 467840 502250 467892 502256
rect 466460 500948 466512 500954
rect 466460 500890 466512 500896
rect 465080 499520 465132 499526
rect 465080 499462 465132 499468
rect 463700 496800 463752 496806
rect 463700 496742 463752 496748
rect 462320 495440 462372 495446
rect 462320 495382 462372 495388
rect 461032 492652 461084 492658
rect 461032 492594 461084 492600
rect 460940 491292 460992 491298
rect 460940 491234 460992 491240
rect 459560 488504 459612 488510
rect 459560 488446 459612 488452
rect 458180 487144 458232 487150
rect 458180 487086 458232 487092
rect 456800 484356 456852 484362
rect 456800 484298 456852 484304
rect 455420 482996 455472 483002
rect 455420 482938 455472 482944
rect 453396 480208 453448 480214
rect 453396 480150 453448 480156
rect 513378 412720 513434 412729
rect 513378 412655 513380 412664
rect 513432 412655 513434 412664
rect 513380 412626 513432 412632
rect 453304 411936 453356 411942
rect 453304 411878 453356 411884
rect 438768 410644 438820 410650
rect 438768 410586 438820 410592
rect 438400 410576 438452 410582
rect 438400 410518 438452 410524
rect 293224 318776 293276 318782
rect 313280 318776 313332 318782
rect 293224 318718 293276 318724
rect 313278 318744 313280 318753
rect 405004 318776 405056 318782
rect 313332 318744 313334 318753
rect 291844 318640 291896 318646
rect 291844 318582 291896 318588
rect 289084 318572 289136 318578
rect 289084 318514 289136 318520
rect 286324 318368 286376 318374
rect 279698 318336 279754 318345
rect 286324 318310 286376 318316
rect 279698 318271 279754 318280
rect 279620 318022 280016 318050
rect 279988 8945 280016 318022
rect 280068 317892 280120 317898
rect 280068 317834 280120 317840
rect 279974 8936 280030 8945
rect 279974 8871 280030 8880
rect 280080 4865 280108 317834
rect 284760 8424 284812 8430
rect 284760 8366 284812 8372
rect 281264 8356 281316 8362
rect 281264 8298 281316 8304
rect 280066 4856 280122 4865
rect 280066 4791 280122 4800
rect 279424 2848 279476 2854
rect 279424 2790 279476 2796
rect 280068 2372 280120 2378
rect 280068 2314 280120 2320
rect 280080 480 280108 2314
rect 281276 480 281304 8298
rect 283654 5536 283710 5545
rect 283654 5471 283710 5480
rect 282460 3324 282512 3330
rect 282460 3266 282512 3272
rect 282472 480 282500 3266
rect 283668 480 283696 5471
rect 284772 480 284800 8366
rect 286336 2922 286364 318310
rect 287060 13864 287112 13870
rect 287060 13806 287112 13812
rect 285956 2916 286008 2922
rect 285956 2858 286008 2864
rect 286324 2916 286376 2922
rect 286324 2858 286376 2864
rect 285968 480 285996 2858
rect 287072 626 287100 13806
rect 288348 8492 288400 8498
rect 288348 8434 288400 8440
rect 287072 598 287192 626
rect 287164 480 287192 598
rect 288360 480 288388 8434
rect 289096 2990 289124 318514
rect 290738 5400 290794 5409
rect 290738 5335 290794 5344
rect 289544 4004 289596 4010
rect 289544 3946 289596 3952
rect 289084 2984 289136 2990
rect 289084 2926 289136 2932
rect 289556 480 289584 3946
rect 290752 480 290780 5335
rect 291856 3126 291884 318582
rect 291936 8560 291988 8566
rect 291936 8502 291988 8508
rect 291844 3120 291896 3126
rect 291844 3062 291896 3068
rect 291948 480 291976 8502
rect 293236 3330 293264 318718
rect 443092 318776 443144 318782
rect 405004 318718 405056 318724
rect 443090 318744 443092 318753
rect 443144 318744 443146 318753
rect 313278 318679 313334 318688
rect 443090 318679 443146 318688
rect 304264 318300 304316 318306
rect 304264 318242 304316 318248
rect 295984 318028 296036 318034
rect 295984 317970 296036 317976
rect 293960 14000 294012 14006
rect 293960 13942 294012 13948
rect 293132 3324 293184 3330
rect 293132 3266 293184 3272
rect 293224 3324 293276 3330
rect 293224 3266 293276 3272
rect 293144 480 293172 3266
rect 293972 626 294000 13942
rect 295340 13932 295392 13938
rect 295340 13874 295392 13880
rect 293972 598 294368 626
rect 295352 610 295380 13874
rect 295996 4010 296024 317970
rect 296076 317960 296128 317966
rect 296076 317902 296128 317908
rect 295984 4004 296036 4010
rect 295984 3946 296036 3952
rect 296088 3233 296116 317902
rect 302240 14136 302292 14142
rect 302240 14078 302292 14084
rect 298100 14068 298152 14074
rect 298100 14010 298152 14016
rect 297916 5568 297968 5574
rect 297916 5510 297968 5516
rect 296074 3224 296130 3233
rect 296074 3159 296130 3168
rect 296720 2848 296772 2854
rect 296720 2790 296772 2796
rect 294340 480 294368 598
rect 295340 604 295392 610
rect 295340 546 295392 552
rect 295524 604 295576 610
rect 295524 546 295576 552
rect 295536 480 295564 546
rect 296732 480 296760 2790
rect 297928 480 297956 5510
rect 298112 610 298140 14010
rect 301412 5636 301464 5642
rect 301412 5578 301464 5584
rect 300308 4140 300360 4146
rect 300308 4082 300360 4088
rect 298100 604 298152 610
rect 298100 546 298152 552
rect 299112 604 299164 610
rect 299112 546 299164 552
rect 299124 480 299152 546
rect 300320 480 300348 4082
rect 301424 480 301452 5578
rect 302252 626 302280 14078
rect 304276 4146 304304 318242
rect 313292 318238 313320 318679
rect 313280 318232 313332 318238
rect 313280 318174 313332 318180
rect 529388 318164 529440 318170
rect 529388 318106 529440 318112
rect 485780 16584 485832 16590
rect 485780 16526 485832 16532
rect 483020 15836 483072 15842
rect 483020 15778 483072 15784
rect 443000 15768 443052 15774
rect 443000 15710 443052 15716
rect 420920 15700 420972 15706
rect 420920 15642 420972 15648
rect 407120 15632 407172 15638
rect 407120 15574 407172 15580
rect 317420 15564 317472 15570
rect 317420 15506 317472 15512
rect 305000 14204 305052 14210
rect 305000 14146 305052 14152
rect 304264 4140 304316 4146
rect 304264 4082 304316 4088
rect 305012 2922 305040 14146
rect 316040 9852 316092 9858
rect 316040 9794 316092 9800
rect 313280 9784 313332 9790
rect 313280 9726 313332 9732
rect 309140 9716 309192 9722
rect 309140 9658 309192 9664
rect 308588 5772 308640 5778
rect 308588 5714 308640 5720
rect 305092 5704 305144 5710
rect 305092 5646 305144 5652
rect 303804 2916 303856 2922
rect 303804 2858 303856 2864
rect 305000 2916 305052 2922
rect 305000 2858 305052 2864
rect 302252 598 302648 626
rect 302620 480 302648 598
rect 303816 480 303844 2858
rect 305104 2802 305132 5646
rect 307392 4140 307444 4146
rect 307392 4082 307444 4088
rect 306196 2916 306248 2922
rect 306196 2858 306248 2864
rect 305012 2774 305132 2802
rect 305012 480 305040 2774
rect 306208 480 306236 2858
rect 307404 480 307432 4082
rect 308600 480 308628 5714
rect 309152 610 309180 9658
rect 312176 5840 312228 5846
rect 312176 5782 312228 5788
rect 310980 4072 311032 4078
rect 310980 4014 311032 4020
rect 309140 604 309192 610
rect 309140 546 309192 552
rect 309784 604 309836 610
rect 309784 546 309836 552
rect 309796 480 309824 546
rect 310992 480 311020 4014
rect 312188 480 312216 5782
rect 313292 626 313320 9726
rect 315764 5908 315816 5914
rect 315764 5850 315816 5856
rect 314566 3360 314622 3369
rect 314566 3295 314622 3304
rect 313292 598 313412 626
rect 313384 480 313412 598
rect 314580 480 314608 3295
rect 315776 480 315804 5850
rect 316052 610 316080 9794
rect 317432 610 317460 15506
rect 405740 14408 405792 14414
rect 405740 14350 405792 14356
rect 401600 14340 401652 14346
rect 401600 14282 401652 14288
rect 390560 14272 390612 14278
rect 390560 14214 390612 14220
rect 385040 12980 385092 12986
rect 385040 12922 385092 12928
rect 378140 12912 378192 12918
rect 378140 12854 378192 12860
rect 374000 12844 374052 12850
rect 374000 12786 374052 12792
rect 371240 12776 371292 12782
rect 371240 12718 371292 12724
rect 364340 12708 364392 12714
rect 364340 12650 364392 12656
rect 356060 12640 356112 12646
rect 356060 12582 356112 12588
rect 349160 12572 349212 12578
rect 349160 12514 349212 12520
rect 342260 12504 342312 12510
rect 342260 12446 342312 12452
rect 340880 11008 340932 11014
rect 340880 10950 340932 10956
rect 338120 10260 338172 10266
rect 338120 10202 338172 10208
rect 333980 10192 334032 10198
rect 333980 10134 334032 10140
rect 331312 10124 331364 10130
rect 331312 10066 331364 10072
rect 327080 10056 327132 10062
rect 327080 9998 327132 10004
rect 322940 9988 322992 9994
rect 322940 9930 322992 9936
rect 320180 9920 320232 9926
rect 320180 9862 320232 9868
rect 319260 5976 319312 5982
rect 319260 5918 319312 5924
rect 316040 604 316092 610
rect 316040 546 316092 552
rect 316960 604 317012 610
rect 316960 546 317012 552
rect 317420 604 317472 610
rect 317420 546 317472 552
rect 318064 604 318116 610
rect 318064 546 318116 552
rect 316972 480 317000 546
rect 318076 480 318104 546
rect 319272 480 319300 5918
rect 320192 626 320220 9862
rect 322848 6044 322900 6050
rect 322848 5986 322900 5992
rect 321650 3360 321706 3369
rect 321650 3295 321706 3304
rect 321834 3360 321890 3369
rect 321834 3295 321890 3304
rect 320192 598 320496 626
rect 320468 480 320496 598
rect 321664 480 321692 3295
rect 321848 3097 321876 3295
rect 321834 3088 321890 3097
rect 321834 3023 321890 3032
rect 322860 480 322888 5986
rect 322952 610 322980 9930
rect 326436 6112 326488 6118
rect 326436 6054 326488 6060
rect 325240 3052 325292 3058
rect 325240 2994 325292 3000
rect 322940 604 322992 610
rect 322940 546 322992 552
rect 324044 604 324096 610
rect 324044 546 324096 552
rect 324056 480 324084 546
rect 325252 480 325280 2994
rect 326448 480 326476 6054
rect 327092 610 327120 9998
rect 330024 6860 330076 6866
rect 330024 6802 330076 6808
rect 328828 3188 328880 3194
rect 328828 3130 328880 3136
rect 327080 604 327132 610
rect 327080 546 327132 552
rect 327632 604 327684 610
rect 327632 546 327684 552
rect 327644 480 327672 546
rect 328840 480 328868 3130
rect 330036 480 330064 6802
rect 331324 626 331352 10066
rect 333612 6792 333664 6798
rect 333612 6734 333664 6740
rect 332416 3936 332468 3942
rect 332416 3878 332468 3884
rect 331232 598 331352 626
rect 331232 480 331260 598
rect 332428 480 332456 3878
rect 333624 480 333652 6734
rect 333992 610 334020 10134
rect 337108 6724 337160 6730
rect 337108 6666 337160 6672
rect 335912 3868 335964 3874
rect 335912 3810 335964 3816
rect 333980 604 334032 610
rect 333980 546 334032 552
rect 334716 604 334768 610
rect 334716 546 334768 552
rect 334728 480 334756 546
rect 335924 480 335952 3810
rect 337120 480 337148 6666
rect 338132 626 338160 10202
rect 340696 6656 340748 6662
rect 340696 6598 340748 6604
rect 339500 3256 339552 3262
rect 339500 3198 339552 3204
rect 338132 598 338344 626
rect 338316 480 338344 598
rect 339512 480 339540 3198
rect 340708 480 340736 6598
rect 340892 610 340920 10950
rect 342272 610 342300 12446
rect 345020 10940 345072 10946
rect 345020 10882 345072 10888
rect 344284 6588 344336 6594
rect 344284 6530 344336 6536
rect 340880 604 340932 610
rect 340880 546 340932 552
rect 341892 604 341944 610
rect 341892 546 341944 552
rect 342260 604 342312 610
rect 342260 546 342312 552
rect 343088 604 343140 610
rect 343088 546 343140 552
rect 341904 480 341932 546
rect 343100 480 343128 546
rect 344296 480 344324 6530
rect 345032 3346 345060 10882
rect 347780 10872 347832 10878
rect 347780 10814 347832 10820
rect 346676 3800 346728 3806
rect 346676 3742 346728 3748
rect 345032 3318 345520 3346
rect 345492 480 345520 3318
rect 346688 480 346716 3742
rect 347792 3262 347820 10814
rect 347870 5264 347926 5273
rect 347870 5199 347926 5208
rect 347780 3256 347832 3262
rect 347780 3198 347832 3204
rect 347884 480 347912 5199
rect 349172 3346 349200 12514
rect 351920 10804 351972 10810
rect 351920 10746 351972 10752
rect 351368 6520 351420 6526
rect 351368 6462 351420 6468
rect 349172 3318 350304 3346
rect 349068 3256 349120 3262
rect 349068 3198 349120 3204
rect 349080 480 349108 3198
rect 350276 480 350304 3318
rect 351380 480 351408 6462
rect 351932 3346 351960 10746
rect 354956 6452 355008 6458
rect 354956 6394 355008 6400
rect 351932 3318 352604 3346
rect 352576 480 352604 3318
rect 353760 2984 353812 2990
rect 353760 2926 353812 2932
rect 353772 480 353800 2926
rect 354968 480 354996 6394
rect 356072 3738 356100 12582
rect 356152 10736 356204 10742
rect 356152 10678 356204 10684
rect 356060 3732 356112 3738
rect 356060 3674 356112 3680
rect 356164 480 356192 10678
rect 358820 10668 358872 10674
rect 358820 10610 358872 10616
rect 358544 6384 358596 6390
rect 358544 6326 358596 6332
rect 357348 3732 357400 3738
rect 357348 3674 357400 3680
rect 357360 480 357388 3674
rect 358556 480 358584 6326
rect 358832 3346 358860 10610
rect 362960 10600 363012 10606
rect 362960 10542 363012 10548
rect 362130 6760 362186 6769
rect 362130 6695 362186 6704
rect 360936 3800 360988 3806
rect 360936 3742 360988 3748
rect 358832 3318 359780 3346
rect 359752 480 359780 3318
rect 360948 480 360976 3742
rect 362144 480 362172 6695
rect 362972 3346 363000 10542
rect 362972 3318 363368 3346
rect 363340 480 363368 3318
rect 364352 610 364380 12650
rect 365720 10532 365772 10538
rect 365720 10474 365772 10480
rect 365732 1426 365760 10474
rect 369860 10464 369912 10470
rect 369860 10406 369912 10412
rect 365810 6624 365866 6633
rect 365810 6559 365866 6568
rect 365720 1420 365772 1426
rect 365720 1362 365772 1368
rect 365824 626 365852 6559
rect 369216 6316 369268 6322
rect 369216 6258 369268 6264
rect 368020 3120 368072 3126
rect 368020 3062 368072 3068
rect 366916 1420 366968 1426
rect 366916 1362 366968 1368
rect 364340 604 364392 610
rect 364340 546 364392 552
rect 364524 604 364576 610
rect 364524 546 364576 552
rect 365732 598 365852 626
rect 364536 480 364564 546
rect 365732 480 365760 598
rect 366928 480 366956 1362
rect 368032 480 368060 3062
rect 369228 480 369256 6258
rect 369872 610 369900 10406
rect 371252 626 371280 12718
rect 372802 6488 372858 6497
rect 372802 6423 372858 6432
rect 369860 604 369912 610
rect 369860 546 369912 552
rect 370412 604 370464 610
rect 371252 598 371648 626
rect 370412 546 370464 552
rect 370424 480 370452 546
rect 371620 480 371648 598
rect 372816 480 372844 6423
rect 374012 3738 374040 12786
rect 374092 10396 374144 10402
rect 374092 10338 374144 10344
rect 374000 3732 374052 3738
rect 374000 3674 374052 3680
rect 374104 1442 374132 10338
rect 376760 10328 376812 10334
rect 376760 10270 376812 10276
rect 376392 4208 376444 4214
rect 376392 4150 376444 4156
rect 375196 3732 375248 3738
rect 375196 3674 375248 3680
rect 374012 1414 374132 1442
rect 374012 480 374040 1414
rect 375208 480 375236 3674
rect 376404 480 376432 4150
rect 376772 610 376800 10270
rect 378152 610 378180 12854
rect 380898 10840 380954 10849
rect 380898 10775 380954 10784
rect 379978 6352 380034 6361
rect 379978 6287 380034 6296
rect 376760 604 376812 610
rect 376760 546 376812 552
rect 377588 604 377640 610
rect 377588 546 377640 552
rect 378140 604 378192 610
rect 378140 546 378192 552
rect 378784 604 378836 610
rect 378784 546 378836 552
rect 377600 480 377628 546
rect 378796 480 378824 546
rect 379992 480 380020 6287
rect 380912 626 380940 10775
rect 383658 10704 383714 10713
rect 383658 10639 383714 10648
rect 383568 4276 383620 4282
rect 383568 4218 383620 4224
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 380912 598 381216 626
rect 381188 480 381216 598
rect 382384 480 382412 3334
rect 383580 480 383608 4218
rect 383672 3346 383700 10639
rect 385052 3346 385080 12922
rect 388260 8628 388312 8634
rect 388260 8570 388312 8576
rect 387062 6216 387118 6225
rect 387062 6151 387118 6160
rect 383672 3318 384712 3346
rect 385052 3318 385908 3346
rect 384684 480 384712 3318
rect 385880 480 385908 3318
rect 387076 480 387104 6151
rect 388272 480 388300 8570
rect 389456 3664 389508 3670
rect 389456 3606 389508 3612
rect 389468 480 389496 3606
rect 390572 1578 390600 14214
rect 391940 13048 391992 13054
rect 391940 12990 391992 12996
rect 390650 10568 390706 10577
rect 390650 10503 390706 10512
rect 390664 3398 390692 10503
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391952 3346 391980 12990
rect 394698 10432 394754 10441
rect 394698 10367 394754 10376
rect 394240 4344 394292 4350
rect 394240 4286 394292 4292
rect 390572 1550 390692 1578
rect 390664 480 390692 1550
rect 391860 480 391888 3334
rect 391952 3318 393084 3346
rect 393056 480 393084 3318
rect 394252 480 394280 4286
rect 394712 3346 394740 10367
rect 398838 10296 398894 10305
rect 398838 10231 398894 10240
rect 397828 7064 397880 7070
rect 397828 7006 397880 7012
rect 396632 3596 396684 3602
rect 396632 3538 396684 3544
rect 394712 3318 395476 3346
rect 395448 480 395476 3318
rect 396644 480 396672 3538
rect 397840 480 397868 7006
rect 398852 3346 398880 10231
rect 401324 7132 401376 7138
rect 401324 7074 401376 7080
rect 398852 3318 399064 3346
rect 399036 480 399064 3318
rect 400220 3324 400272 3330
rect 400220 3266 400272 3272
rect 400232 480 400260 3266
rect 401336 480 401364 7074
rect 401612 3346 401640 14282
rect 402980 13796 403032 13802
rect 402980 13738 403032 13744
rect 402992 3482 403020 13738
rect 404912 7200 404964 7206
rect 404912 7142 404964 7148
rect 402992 3454 403756 3482
rect 401612 3318 402560 3346
rect 402532 480 402560 3318
rect 403728 480 403756 3454
rect 404924 480 404952 7142
rect 405752 3482 405780 14350
rect 407132 3482 407160 15574
rect 408500 15156 408552 15162
rect 408500 15098 408552 15104
rect 408512 3602 408540 15098
rect 414020 13728 414072 13734
rect 414020 13670 414072 13676
rect 412640 11144 412692 11150
rect 412640 11086 412692 11092
rect 412088 7336 412140 7342
rect 412088 7278 412140 7284
rect 408592 7268 408644 7274
rect 408592 7210 408644 7216
rect 408500 3596 408552 3602
rect 408500 3538 408552 3544
rect 408604 3482 408632 7210
rect 409696 3596 409748 3602
rect 409696 3538 409748 3544
rect 405752 3454 406148 3482
rect 407132 3454 407344 3482
rect 406120 480 406148 3454
rect 407316 480 407344 3454
rect 408512 3454 408632 3482
rect 408512 480 408540 3454
rect 409708 480 409736 3538
rect 410892 3528 410944 3534
rect 410892 3470 410944 3476
rect 410904 480 410932 3470
rect 412100 480 412128 7278
rect 412652 610 412680 11086
rect 414032 626 414060 13670
rect 419540 11280 419592 11286
rect 419540 11222 419592 11228
rect 416872 11212 416924 11218
rect 416872 11154 416924 11160
rect 415676 7404 415728 7410
rect 415676 7346 415728 7352
rect 412640 604 412692 610
rect 412640 546 412692 552
rect 413284 604 413336 610
rect 414032 598 414520 626
rect 413284 546 413336 552
rect 413296 480 413324 546
rect 414492 480 414520 598
rect 415688 480 415716 7346
rect 416884 480 416912 11154
rect 419172 7472 419224 7478
rect 419172 7414 419224 7420
rect 417976 4004 418028 4010
rect 417976 3946 418028 3952
rect 417988 480 418016 3946
rect 419184 480 419212 7414
rect 419552 610 419580 11222
rect 420932 610 420960 15642
rect 431960 15088 432012 15094
rect 431960 15030 432012 15036
rect 425060 13660 425112 13666
rect 425060 13602 425112 13608
rect 423680 11348 423732 11354
rect 423680 11290 423732 11296
rect 422760 7540 422812 7546
rect 422760 7482 422812 7488
rect 419540 604 419592 610
rect 419540 546 419592 552
rect 420368 604 420420 610
rect 420368 546 420420 552
rect 420920 604 420972 610
rect 420920 546 420972 552
rect 421564 604 421616 610
rect 421564 546 421616 552
rect 420380 480 420408 546
rect 421576 480 421604 546
rect 422772 480 422800 7482
rect 423692 610 423720 11290
rect 425072 626 425100 13602
rect 430580 11484 430632 11490
rect 430580 11426 430632 11432
rect 426440 11416 426492 11422
rect 426440 11358 426492 11364
rect 426348 8288 426400 8294
rect 426348 8230 426400 8236
rect 423680 604 423732 610
rect 423680 546 423732 552
rect 423956 604 424008 610
rect 425072 598 425192 626
rect 423956 546 424008 552
rect 423968 480 423996 546
rect 425164 480 425192 598
rect 426360 480 426388 8230
rect 426452 610 426480 11358
rect 429936 8220 429988 8226
rect 429936 8162 429988 8168
rect 428740 3460 428792 3466
rect 428740 3402 428792 3408
rect 426440 604 426492 610
rect 426440 546 426492 552
rect 427544 604 427596 610
rect 427544 546 427596 552
rect 427556 480 427584 546
rect 428752 480 428780 3402
rect 429948 480 429976 8162
rect 430592 610 430620 11426
rect 431972 626 432000 15030
rect 438860 15020 438912 15026
rect 438860 14962 438912 14968
rect 437480 11620 437532 11626
rect 437480 11562 437532 11568
rect 433340 11552 433392 11558
rect 433340 11494 433392 11500
rect 433352 3534 433380 11494
rect 433524 8152 433576 8158
rect 433524 8094 433576 8100
rect 433340 3528 433392 3534
rect 433340 3470 433392 3476
rect 430580 604 430632 610
rect 430580 546 430632 552
rect 431132 604 431184 610
rect 431972 598 432276 626
rect 432248 592 432276 598
rect 432248 564 432368 592
rect 431132 546 431184 552
rect 431144 480 431172 546
rect 432340 480 432368 564
rect 433536 480 433564 8094
rect 437020 8084 437072 8090
rect 437020 8026 437072 8032
rect 434628 3528 434680 3534
rect 434628 3470 434680 3476
rect 434640 480 434668 3470
rect 435822 3224 435878 3233
rect 435822 3159 435878 3168
rect 435836 480 435864 3159
rect 437032 480 437060 8026
rect 437492 626 437520 11562
rect 437492 598 438164 626
rect 438872 610 438900 14962
rect 441620 11688 441672 11694
rect 441620 11630 441672 11636
rect 440608 8016 440660 8022
rect 440608 7958 440660 7964
rect 438136 592 438164 598
rect 438860 604 438912 610
rect 438136 564 438256 592
rect 438228 480 438256 564
rect 438860 546 438912 552
rect 439412 604 439464 610
rect 439412 546 439464 552
rect 439424 480 439452 546
rect 440620 480 440648 7958
rect 441632 610 441660 11630
rect 441620 604 441672 610
rect 441620 546 441672 552
rect 441804 604 441856 610
rect 441804 546 441856 552
rect 441816 480 441844 546
rect 443012 480 443040 15710
rect 445760 14952 445812 14958
rect 445760 14894 445812 14900
rect 444380 12436 444432 12442
rect 444380 12378 444432 12384
rect 444196 7948 444248 7954
rect 444196 7890 444248 7896
rect 444208 480 444236 7890
rect 444392 610 444420 12378
rect 445772 610 445800 14894
rect 452660 14884 452712 14890
rect 452660 14826 452712 14832
rect 448520 12368 448572 12374
rect 448520 12310 448572 12316
rect 447784 7880 447836 7886
rect 447784 7822 447836 7828
rect 444380 604 444432 610
rect 444380 546 444432 552
rect 445392 604 445444 610
rect 445392 546 445444 552
rect 445760 604 445812 610
rect 445760 546 445812 552
rect 446588 604 446640 610
rect 446588 546 446640 552
rect 445404 480 445432 546
rect 446600 480 446628 546
rect 447796 480 447824 7822
rect 448532 610 448560 12310
rect 451280 12300 451332 12306
rect 451280 12242 451332 12248
rect 450174 4040 450230 4049
rect 450174 3975 450230 3984
rect 448520 604 448572 610
rect 448520 546 448572 552
rect 448980 604 449032 610
rect 448980 546 449032 552
rect 448992 480 449020 546
rect 450188 480 450216 3975
rect 451292 3534 451320 12242
rect 451372 7812 451424 7818
rect 451372 7754 451424 7760
rect 451280 3528 451332 3534
rect 451280 3470 451332 3476
rect 451384 1442 451412 7754
rect 452476 3528 452528 3534
rect 452476 3470 452528 3476
rect 451292 1414 451412 1442
rect 451292 480 451320 1414
rect 452488 480 452516 3470
rect 452672 610 452700 14826
rect 459560 14816 459612 14822
rect 459560 14758 459612 14764
rect 455420 12232 455472 12238
rect 455420 12174 455472 12180
rect 454868 7744 454920 7750
rect 454868 7686 454920 7692
rect 452660 604 452712 610
rect 452660 546 452712 552
rect 453672 604 453724 610
rect 453672 546 453724 552
rect 453684 480 453712 546
rect 454880 480 454908 7686
rect 455432 610 455460 12174
rect 458456 7676 458508 7682
rect 458456 7618 458508 7624
rect 457258 3904 457314 3913
rect 457258 3839 457314 3848
rect 455420 604 455472 610
rect 455420 546 455472 552
rect 456064 604 456116 610
rect 456064 546 456116 552
rect 456076 480 456104 546
rect 457272 480 457300 3839
rect 458468 480 458496 7618
rect 459572 3534 459600 14758
rect 467840 14748 467892 14754
rect 467840 14690 467892 14696
rect 459652 12164 459704 12170
rect 459652 12106 459704 12112
rect 459560 3528 459612 3534
rect 459560 3470 459612 3476
rect 459664 480 459692 12106
rect 462320 12096 462372 12102
rect 462320 12038 462372 12044
rect 462044 7608 462096 7614
rect 462044 7550 462096 7556
rect 460848 3528 460900 3534
rect 460848 3470 460900 3476
rect 460860 480 460888 3470
rect 462056 480 462084 7550
rect 462332 610 462360 12038
rect 466460 12028 466512 12034
rect 466460 11970 466512 11976
rect 465630 8256 465686 8265
rect 465630 8191 465686 8200
rect 464434 3768 464490 3777
rect 464434 3703 464490 3712
rect 462320 604 462372 610
rect 462320 546 462372 552
rect 463240 604 463292 610
rect 463240 546 463292 552
rect 463252 480 463280 546
rect 464448 480 464476 3703
rect 465644 480 465672 8191
rect 466472 610 466500 11970
rect 467852 626 467880 14690
rect 474740 14680 474792 14686
rect 474740 14622 474792 14628
rect 469220 11960 469272 11966
rect 469220 11902 469272 11908
rect 469126 8120 469182 8129
rect 469126 8055 469182 8064
rect 466460 604 466512 610
rect 466460 546 466512 552
rect 466828 604 466880 610
rect 467852 598 467972 626
rect 466828 546 466880 552
rect 466840 480 466868 546
rect 467944 480 467972 598
rect 469140 480 469168 8055
rect 469232 610 469260 11902
rect 473360 11892 473412 11898
rect 473360 11834 473412 11840
rect 472714 7984 472770 7993
rect 472714 7919 472770 7928
rect 471518 3632 471574 3641
rect 471518 3567 471574 3576
rect 469220 604 469272 610
rect 469220 546 469272 552
rect 470324 604 470376 610
rect 470324 546 470376 552
rect 470336 480 470364 546
rect 471532 480 471560 3567
rect 472728 480 472756 7919
rect 473372 626 473400 11834
rect 474752 626 474780 14622
rect 481640 14612 481692 14618
rect 481640 14554 481692 14560
rect 477500 11824 477552 11830
rect 477500 11766 477552 11772
rect 476302 7848 476358 7857
rect 476302 7783 476358 7792
rect 473372 598 473860 626
rect 474752 598 475056 626
rect 473832 592 473860 598
rect 475028 592 475056 598
rect 473832 564 473952 592
rect 475028 564 475148 592
rect 473924 480 473952 564
rect 475120 480 475148 564
rect 476316 480 476344 7783
rect 477512 480 477540 11766
rect 480260 11756 480312 11762
rect 480260 11698 480312 11704
rect 479890 7712 479946 7721
rect 479890 7647 479946 7656
rect 478694 3496 478750 3505
rect 478694 3431 478750 3440
rect 478708 480 478736 3431
rect 479904 480 479932 7647
rect 480272 3482 480300 11698
rect 481652 3482 481680 14554
rect 483032 3482 483060 15778
rect 484582 7576 484638 7585
rect 484582 7511 484638 7520
rect 480272 3454 481128 3482
rect 481652 3454 482324 3482
rect 483032 3454 483520 3482
rect 481100 480 481128 3454
rect 482296 480 482324 3454
rect 483492 480 483520 3454
rect 484596 480 484624 7511
rect 485792 3602 485820 16526
rect 489920 16516 489972 16522
rect 489920 16458 489972 16464
rect 487160 14544 487212 14550
rect 487160 14486 487212 14492
rect 485870 12200 485926 12209
rect 485870 12135 485926 12144
rect 485780 3596 485832 3602
rect 485780 3538 485832 3544
rect 485884 3482 485912 12135
rect 486976 3596 487028 3602
rect 486976 3538 487028 3544
rect 485792 3454 485912 3482
rect 485792 480 485820 3454
rect 486988 480 487016 3538
rect 487172 3482 487200 14486
rect 488538 12064 488594 12073
rect 488538 11999 488594 12008
rect 488552 3482 488580 11999
rect 487172 3454 488212 3482
rect 488552 3454 489408 3482
rect 488184 480 488212 3454
rect 489380 480 489408 3454
rect 489932 610 489960 16458
rect 494060 16448 494112 16454
rect 494060 16390 494112 16396
rect 491300 14476 491352 14482
rect 491300 14418 491352 14424
rect 491312 626 491340 14418
rect 492678 11928 492734 11937
rect 492678 11863 492734 11872
rect 492692 626 492720 11863
rect 494072 3466 494100 16390
rect 494152 16380 494204 16386
rect 494152 16322 494204 16328
rect 494060 3460 494112 3466
rect 494060 3402 494112 3408
rect 489920 604 489972 610
rect 489920 546 489972 552
rect 490564 604 490616 610
rect 491312 598 491708 626
rect 492692 598 492904 626
rect 491680 592 491708 598
rect 492876 592 492904 598
rect 491680 564 491800 592
rect 492876 564 492996 592
rect 490564 546 490616 552
rect 490576 480 490604 546
rect 491772 480 491800 564
rect 492968 480 492996 564
rect 494164 480 494192 16322
rect 496820 16312 496872 16318
rect 496820 16254 496872 16260
rect 495438 11792 495494 11801
rect 495438 11727 495494 11736
rect 495348 3460 495400 3466
rect 495348 3402 495400 3408
rect 495360 480 495388 3402
rect 495452 610 495480 11727
rect 496832 610 496860 16254
rect 500960 16244 501012 16250
rect 500960 16186 501012 16192
rect 499578 11656 499634 11665
rect 499578 11591 499634 11600
rect 498936 8696 498988 8702
rect 498936 8638 498988 8644
rect 495440 604 495492 610
rect 495440 546 495492 552
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496820 604 496872 610
rect 496820 546 496872 552
rect 497740 604 497792 610
rect 497740 546 497792 552
rect 496556 480 496584 546
rect 497752 480 497780 546
rect 498948 480 498976 8638
rect 499592 610 499620 11591
rect 500972 610 501000 16186
rect 503720 16176 503772 16182
rect 503720 16118 503772 16124
rect 502338 15056 502394 15065
rect 502338 14991 502394 15000
rect 502352 3534 502380 14991
rect 502432 8764 502484 8770
rect 502432 8706 502484 8712
rect 502340 3528 502392 3534
rect 502340 3470 502392 3476
rect 499580 604 499632 610
rect 499580 546 499632 552
rect 500132 604 500184 610
rect 500132 546 500184 552
rect 500960 604 501012 610
rect 500960 546 501012 552
rect 501236 604 501288 610
rect 501236 546 501288 552
rect 500144 480 500172 546
rect 501248 480 501276 546
rect 502444 480 502472 8706
rect 503628 3528 503680 3534
rect 503628 3470 503680 3476
rect 503640 480 503668 3470
rect 503732 610 503760 16118
rect 507860 16108 507912 16114
rect 507860 16050 507912 16056
rect 506478 14920 506534 14929
rect 506478 14855 506534 14864
rect 506020 8832 506072 8838
rect 506020 8774 506072 8780
rect 503720 604 503772 610
rect 503720 546 503772 552
rect 504824 604 504876 610
rect 504824 546 504876 552
rect 504836 480 504864 546
rect 506032 480 506060 8774
rect 506492 610 506520 14855
rect 507872 610 507900 16050
rect 510618 14784 510674 14793
rect 510618 14719 510674 14728
rect 509608 8900 509660 8906
rect 509608 8842 509660 8848
rect 506480 604 506532 610
rect 506480 546 506532 552
rect 507216 604 507268 610
rect 507216 546 507268 552
rect 507860 604 507912 610
rect 507860 546 507912 552
rect 508412 604 508464 610
rect 508412 546 508464 552
rect 507228 480 507256 546
rect 508424 480 508452 546
rect 509620 480 509648 8842
rect 510632 610 510660 14719
rect 513378 14648 513434 14657
rect 513378 14583 513434 14592
rect 513196 9648 513248 9654
rect 513196 9590 513248 9596
rect 512000 4412 512052 4418
rect 512000 4354 512052 4360
rect 510620 604 510672 610
rect 510620 546 510672 552
rect 510804 604 510856 610
rect 510804 546 510856 552
rect 510816 480 510844 546
rect 512012 480 512040 4354
rect 513208 480 513236 9590
rect 513392 610 513420 14583
rect 517520 13592 517572 13598
rect 517520 13534 517572 13540
rect 516784 9580 516836 9586
rect 516784 9522 516836 9528
rect 515588 4480 515640 4486
rect 515588 4422 515640 4428
rect 513380 604 513432 610
rect 513380 546 513432 552
rect 514392 604 514444 610
rect 514392 546 514444 552
rect 514404 480 514432 546
rect 515600 480 515628 4422
rect 516796 480 516824 9522
rect 517532 626 517560 13534
rect 520280 13524 520332 13530
rect 520280 13466 520332 13472
rect 519084 4548 519136 4554
rect 519084 4490 519136 4496
rect 517532 598 517928 626
rect 517900 480 517928 598
rect 519096 480 519124 4490
rect 520292 3534 520320 13466
rect 524420 13456 524472 13462
rect 524420 13398 524472 13404
rect 520372 9512 520424 9518
rect 520372 9454 520424 9460
rect 520280 3528 520332 3534
rect 520280 3470 520332 3476
rect 520384 1442 520412 9454
rect 523868 9444 523920 9450
rect 523868 9386 523920 9392
rect 522672 4616 522724 4622
rect 522672 4558 522724 4564
rect 521476 3528 521528 3534
rect 521476 3470 521528 3476
rect 520292 1414 520412 1442
rect 520292 480 520320 1414
rect 521488 480 521516 3470
rect 522684 480 522712 4558
rect 523880 480 523908 9386
rect 524432 610 524460 13398
rect 528560 13388 528612 13394
rect 528560 13330 528612 13336
rect 527456 9376 527508 9382
rect 527456 9318 527508 9324
rect 526260 4684 526312 4690
rect 526260 4626 526312 4632
rect 524420 604 524472 610
rect 524420 546 524472 552
rect 525064 604 525116 610
rect 525064 546 525116 552
rect 525076 480 525104 546
rect 526272 480 526300 4626
rect 527468 480 527496 9318
rect 528572 3482 528600 13330
rect 528572 3454 528692 3482
rect 529400 3466 529428 318106
rect 529480 318096 529532 318102
rect 529480 318038 529532 318044
rect 529492 3534 529520 318038
rect 567200 16040 567252 16046
rect 567200 15982 567252 15988
rect 545118 14512 545174 14521
rect 545118 14447 545174 14456
rect 531320 13320 531372 13326
rect 531320 13262 531372 13268
rect 531042 9616 531098 9625
rect 531042 9551 531098 9560
rect 529848 4752 529900 4758
rect 529848 4694 529900 4700
rect 529480 3528 529532 3534
rect 529480 3470 529532 3476
rect 528664 480 528692 3454
rect 529388 3460 529440 3466
rect 529388 3402 529440 3408
rect 529860 480 529888 4694
rect 531056 480 531084 9551
rect 531332 3482 531360 13262
rect 535460 13252 535512 13258
rect 535460 13194 535512 13200
rect 534540 9308 534592 9314
rect 534540 9250 534592 9256
rect 533436 5500 533488 5506
rect 533436 5442 533488 5448
rect 531332 3454 532280 3482
rect 532252 480 532280 3454
rect 533448 480 533476 5442
rect 534552 480 534580 9250
rect 535472 3482 535500 13194
rect 538220 13184 538272 13190
rect 538220 13126 538272 13132
rect 538126 9480 538182 9489
rect 538126 9415 538182 9424
rect 536932 5432 536984 5438
rect 536932 5374 536984 5380
rect 535472 3454 535776 3482
rect 535748 480 535776 3454
rect 536944 480 536972 5374
rect 538140 480 538168 9415
rect 538232 610 538260 13126
rect 542360 13116 542412 13122
rect 542360 13058 542412 13064
rect 541716 9240 541768 9246
rect 541716 9182 541768 9188
rect 540520 5364 540572 5370
rect 540520 5306 540572 5312
rect 538220 604 538272 610
rect 538220 546 538272 552
rect 539324 604 539376 610
rect 539324 546 539376 552
rect 539336 480 539364 546
rect 540532 480 540560 5306
rect 541728 480 541756 9182
rect 542372 610 542400 13058
rect 544108 5296 544160 5302
rect 544108 5238 544160 5244
rect 542360 604 542412 610
rect 542360 546 542412 552
rect 542912 604 542964 610
rect 542912 546 542964 552
rect 542924 480 542952 546
rect 544120 480 544148 5238
rect 545132 626 545160 14447
rect 546498 13560 546554 13569
rect 546498 13495 546554 13504
rect 545132 598 545344 626
rect 545316 480 545344 598
rect 546512 480 546540 13495
rect 549258 13424 549314 13433
rect 549258 13359 549314 13368
rect 548890 9344 548946 9353
rect 548890 9279 548946 9288
rect 547696 5228 547748 5234
rect 547696 5170 547748 5176
rect 547708 480 547736 5170
rect 548904 480 548932 9279
rect 549272 610 549300 13359
rect 553398 13288 553454 13297
rect 553398 13223 553454 13232
rect 552388 9172 552440 9178
rect 552388 9114 552440 9120
rect 551192 5160 551244 5166
rect 551192 5102 551244 5108
rect 549260 604 549312 610
rect 549260 546 549312 552
rect 550088 604 550140 610
rect 550088 546 550140 552
rect 550100 480 550128 546
rect 551204 480 551232 5102
rect 552400 480 552428 9114
rect 553412 626 553440 13223
rect 556158 13152 556214 13161
rect 556158 13087 556214 13096
rect 555974 9208 556030 9217
rect 555974 9143 556030 9152
rect 554780 5092 554832 5098
rect 554780 5034 554832 5040
rect 553412 598 553624 626
rect 553596 480 553624 598
rect 554792 480 554820 5034
rect 555988 480 556016 9143
rect 556172 610 556200 13087
rect 560298 13016 560354 13025
rect 560298 12951 560354 12960
rect 559564 9104 559616 9110
rect 559564 9046 559616 9052
rect 558368 5024 558420 5030
rect 558368 4966 558420 4972
rect 556160 604 556212 610
rect 556160 546 556212 552
rect 557172 604 557224 610
rect 557172 546 557224 552
rect 557184 480 557212 546
rect 558380 480 558408 4966
rect 559576 480 559604 9046
rect 560312 3482 560340 12951
rect 566740 9036 566792 9042
rect 566740 8978 566792 8984
rect 563152 6248 563204 6254
rect 563152 6190 563204 6196
rect 561956 4956 562008 4962
rect 561956 4898 562008 4904
rect 560312 3454 560800 3482
rect 560772 480 560800 3454
rect 561968 480 561996 4898
rect 563164 480 563192 6190
rect 565544 4888 565596 4894
rect 565544 4830 565596 4836
rect 564348 3528 564400 3534
rect 564348 3470 564400 3476
rect 564360 480 564388 3470
rect 565556 480 565584 4830
rect 566752 480 566780 8978
rect 567212 3482 567240 15982
rect 574100 15972 574152 15978
rect 574100 15914 574152 15920
rect 570234 9072 570290 9081
rect 570234 9007 570290 9016
rect 569040 4820 569092 4826
rect 569040 4762 569092 4768
rect 567212 3454 567884 3482
rect 567856 480 567884 3454
rect 569052 480 569080 4762
rect 570248 480 570276 9007
rect 573824 6180 573876 6186
rect 573824 6122 573876 6128
rect 572626 5128 572682 5137
rect 572626 5063 572682 5072
rect 571432 3460 571484 3466
rect 571432 3402 571484 3408
rect 571444 480 571472 3402
rect 572640 480 572668 5063
rect 573836 480 573864 6122
rect 574112 3482 574140 15914
rect 578240 15904 578292 15910
rect 578240 15846 578292 15852
rect 577412 8968 577464 8974
rect 577412 8910 577464 8916
rect 576214 4992 576270 5001
rect 576214 4927 576270 4936
rect 574112 3454 575060 3482
rect 575032 480 575060 3454
rect 576228 480 576256 4927
rect 577424 480 577452 8910
rect 578252 626 578280 15846
rect 580998 8936 581054 8945
rect 580998 8871 581054 8880
rect 579802 4856 579858 4865
rect 579802 4791 579858 4800
rect 578252 598 578648 626
rect 578620 480 578648 598
rect 579816 480 579844 4791
rect 581012 480 581040 8871
rect 582194 3360 582250 3369
rect 582194 3295 582250 3304
rect 582208 480 582236 3295
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 129278 652840 129334 652896
rect 133694 652840 133750 652896
rect 259182 652876 259184 652896
rect 259184 652876 259236 652896
rect 259236 652876 259238 652896
rect 259182 652840 259238 652876
rect 263598 652876 263600 652896
rect 263600 652876 263652 652896
rect 263652 652876 263654 652896
rect 263598 652840 263654 652876
rect 378138 652876 378140 652896
rect 378140 652876 378192 652896
rect 378192 652876 378194 652896
rect 378138 652840 378194 652876
rect 383566 652876 383568 652896
rect 383568 652876 383620 652896
rect 383620 652876 383622 652896
rect 383566 652840 383622 652876
rect 508410 652860 508466 652896
rect 508410 652840 508412 652860
rect 508412 652840 508464 652860
rect 508464 652840 508466 652860
rect 513378 652860 513434 652896
rect 513378 652840 513380 652860
rect 513380 652840 513432 652860
rect 513432 652840 513434 652860
rect 266450 649848 266506 649904
rect 137650 649655 137706 649711
rect 57886 646040 57942 646096
rect 57794 644952 57850 645008
rect 57702 643184 57758 643240
rect 57610 641960 57666 642016
rect 57518 640328 57574 640384
rect 57426 639240 57482 639296
rect 57334 637608 57390 637664
rect 57242 579672 57298 579728
rect 387154 649848 387210 649904
rect 516414 649848 516470 649904
rect 282274 648624 282330 648680
rect 188342 646040 188398 646096
rect 307390 646040 307446 646096
rect 438122 646040 438178 646096
rect 139398 589600 139454 589656
rect 139398 580352 139454 580408
rect 187698 578992 187754 579048
rect 67546 558864 67602 558920
rect 68926 558864 68982 558920
rect 70214 558864 70270 558920
rect 71686 558864 71742 558920
rect 72514 558864 72570 558920
rect 73066 558864 73122 558920
rect 73710 558864 73766 558920
rect 74262 558864 74318 558920
rect 74998 558864 75054 558920
rect 75826 558864 75882 558920
rect 76838 558864 76894 558920
rect 77390 558864 77446 558920
rect 78586 558864 78642 558920
rect 79322 558864 79378 558920
rect 79966 558864 80022 558920
rect 80794 558864 80850 558920
rect 81254 558864 81310 558920
rect 81990 558864 82046 558920
rect 82726 558864 82782 558920
rect 83830 558864 83886 558920
rect 84198 558864 84254 558920
rect 85486 558864 85542 558920
rect 86774 558864 86830 558920
rect 87878 558864 87934 558920
rect 88246 558864 88302 558920
rect 88890 558864 88946 558920
rect 89350 558864 89406 558920
rect 89810 558864 89866 558920
rect 91006 558864 91062 558920
rect 92294 558864 92350 558920
rect 92478 558864 92534 558920
rect 93674 558864 93730 558920
rect 94870 558864 94926 558920
rect 95054 558864 95110 558920
rect 95698 558864 95754 558920
rect 96526 558864 96582 558920
rect 97078 558864 97134 558920
rect 97630 558864 97686 558920
rect 98550 558864 98606 558920
rect 99286 558864 99342 558920
rect 100574 558864 100630 558920
rect 102046 558864 102102 558920
rect 104806 558864 104862 558920
rect 107474 558864 107530 558920
rect 108486 558864 108542 558920
rect 62026 558320 62082 558376
rect 63406 558184 63462 558240
rect 70306 558728 70362 558784
rect 75918 558728 75974 558784
rect 78494 558728 78550 558784
rect 79506 558748 79562 558784
rect 79506 558728 79508 558748
rect 79508 558728 79560 558748
rect 79560 558728 79562 558748
rect 77574 542952 77630 543008
rect 82910 558728 82966 558784
rect 85394 558728 85450 558784
rect 86682 558612 86738 558648
rect 86682 558592 86684 558612
rect 86684 558592 86736 558612
rect 86736 558592 86738 558612
rect 86866 558728 86922 558784
rect 91098 558728 91154 558784
rect 93582 558592 93638 558648
rect 93766 558728 93822 558784
rect 96250 543224 96306 543280
rect 99378 558476 99434 558512
rect 104898 558748 104954 558784
rect 104898 558728 104900 558748
rect 104900 558728 104952 558748
rect 104952 558728 104954 558748
rect 99378 558456 99380 558476
rect 99380 558456 99432 558476
rect 99432 558456 99434 558476
rect 100022 557776 100078 557832
rect 100850 557660 100906 557696
rect 100850 557640 100852 557660
rect 100852 557640 100904 557660
rect 100904 557640 100906 557660
rect 101402 557640 101458 557696
rect 106278 557640 106334 557696
rect 106922 557640 106978 557696
rect 102046 557504 102102 557560
rect 102782 557504 102838 557560
rect 103426 557504 103482 557560
rect 104162 557504 104218 557560
rect 105542 557504 105598 557560
rect 106186 557504 106242 557560
rect 103426 543088 103482 543144
rect 108302 558456 108358 558512
rect 107658 557504 107714 557560
rect 108486 557504 108542 557560
rect 110326 557504 110382 557560
rect 140042 543632 140098 543688
rect 141422 543360 141478 543416
rect 148322 543496 148378 543552
rect 188434 644952 188490 645008
rect 188526 643184 188582 643240
rect 188618 641960 188674 642016
rect 188710 640328 188766 640384
rect 188802 639240 188858 639296
rect 188894 637608 188950 637664
rect 282182 587152 282238 587208
rect 282182 586472 282238 586528
rect 188986 579672 189042 579728
rect 188342 543224 188398 543280
rect 229374 559952 229430 560008
rect 225970 559816 226026 559872
rect 194414 558864 194470 558920
rect 195978 558864 196034 558920
rect 200210 558884 200266 558920
rect 200210 558864 200212 558884
rect 200212 558864 200264 558884
rect 200264 558864 200266 558884
rect 194414 558048 194470 558104
rect 188986 542952 189042 543008
rect 201498 558864 201554 558920
rect 202786 558864 202842 558920
rect 203798 558864 203854 558920
rect 204166 558864 204222 558920
rect 205546 558864 205602 558920
rect 206374 558864 206430 558920
rect 208490 558864 208546 558920
rect 211894 558864 211950 558920
rect 213090 558864 213146 558920
rect 213918 558864 213974 558920
rect 215298 558864 215354 558920
rect 218794 558864 218850 558920
rect 220082 558864 220138 558920
rect 221094 558864 221150 558920
rect 222290 558864 222346 558920
rect 223578 558864 223634 558920
rect 223946 558864 224002 558920
rect 202142 558728 202198 558784
rect 200026 543632 200082 543688
rect 202050 543088 202106 543144
rect 204902 558592 204958 558648
rect 210514 558592 210570 558648
rect 211158 558592 211214 558648
rect 207662 557640 207718 557696
rect 209042 557640 209098 557696
rect 217966 558748 218022 558784
rect 217966 558728 217968 558748
rect 217968 558728 218020 558748
rect 218020 558728 218022 558748
rect 206926 557504 206982 557560
rect 210974 557640 211030 557696
rect 217874 557640 217930 557696
rect 208306 557504 208362 557560
rect 209686 557504 209742 557560
rect 210422 543496 210478 543552
rect 208306 543360 208362 543416
rect 211066 557504 211122 557560
rect 212446 557504 212502 557560
rect 213826 557504 213882 557560
rect 215206 557504 215262 557560
rect 216586 557504 216642 557560
rect 220726 558628 220728 558648
rect 220728 558628 220780 558648
rect 220780 558628 220782 558648
rect 220726 558592 220782 558628
rect 227258 559272 227314 559328
rect 228086 558864 228142 558920
rect 235906 558864 235962 558920
rect 237286 558864 237342 558920
rect 240046 558864 240102 558920
rect 231950 558728 232006 558784
rect 233238 558728 233294 558784
rect 234618 558748 234674 558784
rect 234618 558728 234620 558748
rect 234620 558728 234672 558748
rect 234672 558728 234674 558748
rect 231858 558612 231914 558648
rect 231858 558592 231860 558612
rect 231860 558592 231912 558612
rect 231912 558592 231914 558612
rect 230478 558456 230534 558512
rect 226246 557640 226302 557696
rect 233146 557640 233202 557696
rect 217966 557504 218022 557560
rect 219346 557504 219402 557560
rect 220726 557504 220782 557560
rect 222106 557504 222162 557560
rect 223486 557504 223542 557560
rect 224866 557504 224922 557560
rect 226154 557504 226210 557560
rect 227626 557504 227682 557560
rect 229006 557504 229062 557560
rect 230386 557504 230442 557560
rect 231766 557504 231822 557560
rect 233054 557504 233110 557560
rect 234526 557504 234582 557560
rect 235998 558728 236054 558784
rect 237378 558592 237434 558648
rect 238758 558340 238814 558376
rect 238758 558320 238760 558340
rect 238760 558320 238812 558340
rect 238812 558320 238814 558340
rect 238666 558048 238722 558104
rect 281722 539008 281778 539064
rect 281722 536968 281778 537024
rect 281722 534928 281778 534984
rect 281722 532888 281778 532944
rect 281722 530848 281778 530904
rect 281722 528808 281778 528864
rect 281722 526768 281778 526824
rect 281722 524728 281778 524784
rect 281722 522688 281778 522744
rect 281722 520648 281778 520704
rect 281722 518608 281778 518664
rect 281722 516568 281778 516624
rect 281722 514528 281778 514584
rect 281722 512488 281778 512544
rect 281722 510448 281778 510504
rect 281722 508408 281778 508464
rect 281722 506404 281724 506424
rect 281724 506404 281776 506424
rect 281776 506404 281778 506424
rect 281722 506368 281778 506404
rect 281722 504328 281778 504384
rect 281722 502308 281778 502344
rect 281722 502288 281724 502308
rect 281724 502288 281776 502308
rect 281776 502288 281778 502308
rect 281722 500248 281778 500304
rect 281722 498208 281778 498264
rect 281722 496168 281778 496224
rect 281722 494128 281778 494184
rect 281722 492088 281778 492144
rect 281722 490048 281778 490104
rect 281722 488008 281778 488064
rect 281722 485968 281778 486024
rect 281722 483928 281778 483984
rect 281722 481888 281778 481944
rect 281722 479848 281778 479904
rect 281722 477808 281778 477864
rect 281722 475768 281778 475824
rect 281722 473728 281778 473784
rect 281722 471688 281778 471744
rect 281722 469648 281778 469704
rect 281722 467608 281778 467664
rect 281722 465568 281778 465624
rect 281722 463528 281778 463584
rect 281722 461488 281778 461544
rect 281722 459484 281724 459504
rect 281724 459484 281776 459504
rect 281776 459484 281778 459504
rect 281722 459448 281778 459484
rect 281722 457408 281778 457464
rect 281722 455388 281778 455424
rect 281722 455368 281724 455388
rect 281724 455368 281776 455388
rect 281776 455368 281778 455388
rect 281722 453328 281778 453384
rect 281722 451288 281778 451344
rect 281722 449248 281778 449304
rect 281722 447208 281778 447264
rect 281722 445168 281778 445224
rect 281722 443128 281778 443184
rect 281722 441088 281778 441144
rect 281722 439048 281778 439104
rect 281722 437008 281778 437064
rect 281722 434968 281778 435024
rect 281722 432928 281778 432984
rect 281722 431024 281778 431080
rect 281722 428984 281778 429040
rect 281722 426944 281778 427000
rect 281722 424904 281778 424960
rect 281722 422864 281778 422920
rect 281722 420860 281724 420880
rect 281724 420860 281776 420880
rect 281776 420860 281778 420880
rect 281722 420824 281778 420860
rect 281722 418784 281778 418840
rect 281722 416744 281778 416800
rect 281722 414704 281778 414760
rect 281722 412664 281778 412720
rect 281814 408584 281870 408640
rect 281998 410624 282054 410680
rect 281906 406544 281962 406600
rect 281722 404504 281778 404560
rect 281538 402464 281594 402520
rect 281630 400424 281686 400480
rect 281722 398384 281778 398440
rect 281538 396344 281594 396400
rect 282090 394304 282146 394360
rect 281906 378020 281908 378040
rect 281908 378020 281960 378040
rect 281960 378020 281962 378040
rect 281906 377984 281962 378020
rect 281722 365780 281724 365800
rect 281724 365780 281776 365800
rect 281776 365780 281778 365800
rect 281722 365744 281778 365780
rect 281906 361664 281962 361720
rect 281906 359624 281962 359680
rect 281722 357620 281724 357640
rect 281724 357620 281776 357640
rect 281776 357620 281778 357640
rect 281722 357584 281778 357620
rect 282090 355544 282146 355600
rect 281538 345344 281594 345400
rect 281538 341300 281540 341320
rect 281540 341300 281592 341320
rect 281592 341300 281594 341320
rect 281538 341264 281594 341300
rect 281722 339260 281724 339280
rect 281724 339260 281776 339280
rect 281776 339260 281778 339280
rect 281722 339224 281778 339260
rect 281538 337184 281594 337240
rect 281630 335180 281632 335200
rect 281632 335180 281684 335200
rect 281684 335180 281686 335200
rect 281630 335144 281686 335180
rect 281538 333104 281594 333160
rect 281538 331100 281540 331120
rect 281540 331100 281592 331120
rect 281592 331100 281594 331120
rect 281538 331064 281594 331100
rect 281538 329060 281540 329080
rect 281540 329060 281592 329080
rect 281592 329060 281594 329080
rect 281538 329024 281594 329060
rect 281538 327020 281540 327040
rect 281540 327020 281592 327040
rect 281592 327020 281594 327040
rect 281538 326984 281594 327020
rect 281538 324944 281594 325000
rect 283654 558184 283710 558240
rect 282826 392264 282882 392320
rect 282734 390224 282790 390280
rect 282642 388184 282698 388240
rect 282550 386144 282606 386200
rect 282458 384104 282514 384160
rect 282366 382064 282422 382120
rect 282274 380024 282330 380080
rect 282826 375944 282882 376000
rect 282826 373940 282828 373960
rect 282828 373940 282880 373960
rect 282880 373940 282882 373960
rect 282826 373904 282882 373940
rect 282826 371864 282882 371920
rect 282366 369824 282422 369880
rect 282274 367784 282330 367840
rect 282826 363704 282882 363760
rect 282826 353504 282882 353560
rect 282826 351464 282882 351520
rect 282826 349424 282882 349480
rect 282826 347656 282882 347712
rect 282826 343304 282882 343360
rect 292578 558612 292634 558648
rect 292578 558592 292580 558612
rect 292580 558592 292632 558612
rect 292632 558592 292634 558612
rect 307114 644952 307170 645008
rect 307114 643456 307170 643512
rect 307666 642096 307722 642152
rect 307666 640464 307722 640520
rect 306654 639376 306710 639432
rect 306838 637880 306894 637936
rect 389178 580896 389234 580952
rect 306930 579944 306986 580000
rect 302146 558592 302202 558648
rect 437846 579128 437902 579184
rect 307666 578892 307668 578912
rect 307668 578892 307720 578912
rect 307720 578892 307722 578912
rect 307666 578856 307722 578892
rect 348422 559272 348478 559328
rect 357714 559272 357770 559328
rect 313738 558864 313794 558920
rect 316038 558864 316094 558920
rect 317418 558884 317474 558920
rect 317418 558864 317420 558884
rect 317420 558864 317472 558884
rect 317472 558864 317474 558884
rect 320270 558864 320326 558920
rect 322846 558864 322902 558920
rect 323490 558864 323546 558920
rect 320178 558748 320234 558784
rect 320178 558728 320180 558748
rect 320180 558728 320232 558748
rect 320232 558728 320234 558748
rect 318798 558592 318854 558648
rect 328550 558864 328606 558920
rect 329562 558864 329618 558920
rect 330482 558864 330538 558920
rect 332506 558864 332562 558920
rect 333150 558864 333206 558920
rect 334254 558884 334310 558920
rect 334254 558864 334256 558884
rect 334256 558864 334308 558884
rect 334308 558864 334310 558884
rect 335910 558864 335966 558920
rect 336278 558864 336334 558920
rect 337750 558864 337806 558920
rect 339038 558864 339094 558920
rect 339866 558864 339922 558920
rect 341246 558864 341302 558920
rect 342534 558864 342590 558920
rect 343638 558884 343694 558920
rect 343638 558864 343640 558884
rect 343640 558864 343692 558884
rect 343692 558864 343694 558884
rect 344834 558884 344890 558920
rect 344834 558864 344836 558884
rect 344836 558864 344888 558884
rect 344888 558864 344890 558884
rect 345754 558864 345810 558920
rect 346490 558864 346546 558920
rect 348238 558864 348294 558920
rect 349342 558864 349398 558920
rect 350538 558864 350594 558920
rect 352010 558864 352066 558920
rect 353298 558884 353354 558920
rect 353298 558864 353300 558884
rect 353300 558864 353352 558884
rect 353352 558864 353354 558884
rect 354678 558728 354734 558784
rect 356058 558728 356114 558784
rect 357438 558476 357494 558512
rect 357438 558456 357440 558476
rect 357440 558456 357492 558476
rect 357492 558456 357494 558476
rect 356702 558320 356758 558376
rect 324962 557640 325018 557696
rect 326342 557640 326398 557696
rect 327722 557640 327778 557696
rect 329930 557640 329986 557696
rect 336830 557640 336886 557696
rect 343730 557640 343786 557696
rect 352010 557640 352066 557696
rect 321558 557504 321614 557560
rect 322938 557504 322994 557560
rect 324318 557504 324374 557560
rect 325698 557504 325754 557560
rect 327078 557504 327134 557560
rect 328458 557504 328514 557560
rect 329838 557504 329894 557560
rect 331218 557504 331274 557560
rect 332598 557504 332654 557560
rect 333978 557504 334034 557560
rect 335358 557504 335414 557560
rect 336738 557504 336794 557560
rect 338118 557504 338174 557560
rect 339498 557504 339554 557560
rect 340878 557504 340934 557560
rect 342258 557504 342314 557560
rect 343638 557504 343694 557560
rect 345018 557504 345074 557560
rect 346398 557504 346454 557560
rect 347778 557504 347834 557560
rect 349158 557504 349214 557560
rect 350538 557504 350594 557560
rect 353298 557504 353354 557560
rect 354678 557504 354734 557560
rect 356058 557504 356114 557560
rect 352194 555464 352250 555520
rect 357530 557504 357586 557560
rect 358910 555464 358966 555520
rect 383566 413244 383568 413264
rect 383568 413244 383620 413264
rect 383620 413244 383622 413264
rect 383566 413208 383622 413244
rect 282182 321000 282238 321056
rect 12346 318416 12402 318472
rect 9586 318144 9642 318200
rect 5446 318008 5502 318064
rect 4066 3440 4122 3496
rect 2870 3304 2926 3360
rect 13634 318280 13690 318336
rect 24306 3576 24362 3632
rect 34978 3712 35034 3768
rect 40958 3984 41014 4040
rect 39762 3848 39818 3904
rect 60738 3440 60794 3496
rect 61934 318008 61990 318064
rect 63314 318144 63370 318200
rect 64142 318416 64198 318472
rect 65062 318280 65118 318336
rect 66350 241440 66406 241496
rect 66534 241440 66590 241496
rect 66350 222128 66406 222184
rect 66534 222128 66590 222184
rect 66350 202816 66406 202872
rect 66534 202816 66590 202872
rect 66350 183504 66406 183560
rect 66534 183504 66590 183560
rect 66350 154536 66406 154592
rect 66626 154536 66682 154592
rect 66350 135224 66406 135280
rect 66626 135224 66682 135280
rect 66350 115912 66406 115968
rect 66626 115912 66682 115968
rect 66350 96600 66406 96656
rect 66626 96600 66682 96656
rect 60830 3304 60886 3360
rect 72054 241440 72110 241496
rect 72238 241440 72294 241496
rect 72054 222128 72110 222184
rect 72238 222128 72294 222184
rect 72054 202816 72110 202872
rect 72238 202816 72294 202872
rect 72054 183504 72110 183560
rect 72238 183504 72294 183560
rect 72238 145016 72294 145072
rect 72238 144880 72294 144936
rect 72238 125704 72294 125760
rect 72238 125568 72294 125624
rect 69294 3576 69350 3632
rect 74262 278704 74318 278760
rect 74446 278704 74502 278760
rect 74262 259392 74318 259448
rect 74446 259392 74502 259448
rect 74262 240080 74318 240136
rect 74446 240080 74502 240136
rect 74262 220768 74318 220824
rect 74446 220768 74502 220824
rect 74262 211112 74318 211168
rect 74446 211112 74502 211168
rect 74262 191800 74318 191856
rect 74446 191800 74502 191856
rect 74262 172488 74318 172544
rect 74446 172488 74502 172544
rect 74446 145016 74502 145072
rect 74446 144880 74502 144936
rect 74446 125704 74502 125760
rect 74446 125568 74502 125624
rect 73250 3712 73306 3768
rect 74814 241440 74870 241496
rect 74998 241440 75054 241496
rect 74814 222128 74870 222184
rect 74998 222128 75054 222184
rect 74814 202816 74870 202872
rect 74998 202816 75054 202872
rect 74814 183504 74870 183560
rect 74998 183504 75054 183560
rect 74998 145016 75054 145072
rect 74998 144880 75054 144936
rect 74998 125704 75054 125760
rect 74998 125568 75054 125624
rect 74722 3984 74778 4040
rect 74630 3848 74686 3904
rect 77574 222128 77630 222184
rect 77758 222128 77814 222184
rect 77482 124208 77538 124264
rect 77850 124208 77906 124264
rect 78862 125704 78918 125760
rect 78770 125588 78826 125624
rect 78770 125568 78772 125588
rect 78772 125568 78824 125588
rect 78824 125568 78826 125588
rect 78862 106392 78918 106448
rect 78770 106256 78826 106312
rect 81714 278740 81716 278760
rect 81716 278740 81768 278760
rect 81768 278740 81770 278760
rect 81714 278704 81770 278740
rect 81898 270408 81954 270464
rect 85854 212472 85910 212528
rect 86130 212472 86186 212528
rect 85854 193160 85910 193216
rect 86130 193160 86186 193216
rect 85946 144900 86002 144936
rect 85946 144880 85948 144900
rect 85948 144880 86000 144900
rect 86000 144880 86002 144900
rect 86130 144880 86186 144936
rect 85854 135224 85910 135280
rect 86038 135224 86094 135280
rect 85946 125588 86002 125624
rect 85946 125568 85948 125588
rect 85948 125568 86000 125588
rect 86000 125568 86002 125588
rect 86130 125568 86186 125624
rect 85854 115912 85910 115968
rect 86038 115912 86094 115968
rect 95422 241440 95478 241496
rect 95606 241440 95662 241496
rect 95422 222128 95478 222184
rect 95606 222128 95662 222184
rect 95422 202816 95478 202872
rect 95606 202816 95662 202872
rect 95422 183504 95478 183560
rect 95606 183504 95662 183560
rect 95422 154536 95478 154592
rect 95698 154536 95754 154592
rect 95422 135224 95478 135280
rect 95698 135224 95754 135280
rect 95422 115912 95478 115968
rect 95698 115912 95754 115968
rect 95422 96600 95478 96656
rect 95698 96600 95754 96656
rect 114466 3304 114522 3360
rect 115754 2896 115810 2952
rect 119986 3440 120042 3496
rect 118606 3032 118662 3088
rect 121366 3576 121422 3632
rect 124310 144880 124366 144936
rect 124586 144880 124642 144936
rect 124310 125568 124366 125624
rect 124586 125568 124642 125624
rect 124310 106256 124366 106312
rect 124586 106256 124642 106312
rect 124310 86944 124366 87000
rect 124586 86944 124642 87000
rect 124494 42064 124550 42120
rect 124402 32408 124458 32464
rect 124034 3168 124090 3224
rect 129554 2796 129556 2816
rect 129556 2796 129608 2816
rect 129608 2796 129610 2816
rect 129554 2760 129610 2796
rect 134614 317908 134616 317928
rect 134616 317908 134668 317928
rect 134668 317908 134670 317928
rect 134614 317872 134670 317908
rect 136454 318144 136510 318200
rect 134982 280064 135038 280120
rect 134982 270544 135038 270600
rect 134982 260752 135038 260808
rect 134982 251232 135038 251288
rect 134798 193160 134854 193216
rect 134982 193160 135038 193216
rect 134798 173848 134854 173904
rect 134982 173848 135038 173904
rect 134706 77288 134762 77344
rect 134890 77288 134946 77344
rect 134890 67768 134946 67824
rect 134890 67632 134946 67688
rect 135074 61376 135130 61432
rect 134982 48320 135038 48376
rect 135074 42064 135130 42120
rect 134982 29008 135038 29064
rect 137926 317872 137982 317928
rect 133970 2796 133972 2816
rect 133972 2796 134024 2816
rect 134024 2796 134026 2816
rect 133970 2760 134026 2796
rect 140870 183504 140926 183560
rect 141146 183504 141202 183560
rect 140686 3984 140742 4040
rect 142066 3848 142122 3904
rect 143446 3712 143502 3768
rect 144458 3304 144514 3360
rect 144826 3304 144882 3360
rect 146850 2896 146906 2952
rect 149702 318416 149758 318472
rect 149702 318144 149758 318200
rect 150070 183504 150126 183560
rect 150254 183504 150310 183560
rect 150162 77152 150218 77208
rect 150346 77152 150402 77208
rect 153934 3032 153990 3088
rect 157890 318144 157946 318200
rect 158718 3440 158774 3496
rect 160558 202816 160614 202872
rect 160742 202816 160798 202872
rect 159362 3032 159418 3088
rect 162306 3576 162362 3632
rect 162122 3440 162178 3496
rect 162766 3440 162822 3496
rect 162766 3032 162822 3088
rect 164146 5072 164202 5128
rect 165526 4936 165582 4992
rect 166906 4800 166962 4856
rect 168286 5480 168342 5536
rect 169666 5344 169722 5400
rect 169390 3168 169446 3224
rect 172334 4800 172390 4856
rect 172518 4800 172574 4856
rect 171782 3032 171838 3088
rect 176566 4256 176622 4312
rect 176750 4256 176806 4312
rect 176474 4120 176530 4176
rect 176842 4120 176898 4176
rect 176750 3032 176806 3088
rect 178682 318144 178738 318200
rect 178682 4120 178738 4176
rect 181350 318008 181406 318064
rect 180706 4800 180762 4856
rect 180706 4528 180762 4584
rect 182086 4800 182142 4856
rect 182086 4528 182142 4584
rect 181534 4120 181590 4176
rect 186134 3168 186190 3224
rect 186410 3168 186466 3224
rect 191654 5208 191710 5264
rect 197174 6704 197230 6760
rect 198646 6568 198702 6624
rect 204074 10784 204130 10840
rect 201406 6432 201462 6488
rect 205454 10648 205510 10704
rect 204166 6296 204222 6352
rect 205454 4800 205510 4856
rect 205454 4528 205510 4584
rect 206834 6160 206890 6216
rect 208306 10512 208362 10568
rect 209502 10376 209558 10432
rect 210974 10240 211030 10296
rect 212446 4800 212502 4856
rect 212446 4528 212502 4584
rect 211066 3984 211122 4040
rect 214654 3848 214710 3904
rect 218150 3712 218206 3768
rect 221738 3304 221794 3360
rect 230386 3984 230442 4040
rect 231766 4528 231822 4584
rect 231766 4120 231822 4176
rect 235814 8200 235870 8256
rect 233146 3848 233202 3904
rect 234526 4528 234582 4584
rect 234710 4392 234766 4448
rect 237286 8064 237342 8120
rect 238574 7928 238630 7984
rect 235906 3712 235962 3768
rect 234802 3440 234858 3496
rect 240046 7792 240102 7848
rect 241334 7656 241390 7712
rect 238390 3576 238446 3632
rect 238666 3576 238722 3632
rect 241426 3440 241482 3496
rect 244186 12144 244242 12200
rect 245566 12008 245622 12064
rect 242806 7520 242862 7576
rect 244094 4392 244150 4448
rect 244278 4392 244334 4448
rect 246946 11872 247002 11928
rect 248234 11736 248290 11792
rect 249614 11600 249670 11656
rect 250994 15000 251050 15056
rect 252374 14864 252430 14920
rect 253662 14728 253718 14784
rect 255042 14592 255098 14648
rect 260654 9560 260710 9616
rect 259366 4528 259422 4584
rect 259366 4256 259422 4312
rect 263414 9424 263470 9480
rect 266082 14456 266138 14512
rect 266174 13504 266230 13560
rect 267462 13368 267518 13424
rect 267554 9288 267610 9344
rect 268842 13232 268898 13288
rect 270222 13096 270278 13152
rect 270314 9152 270370 9208
rect 271602 12960 271658 13016
rect 272890 5072 272946 5128
rect 273442 4256 273498 4312
rect 275834 9016 275890 9072
rect 277306 5072 277362 5128
rect 276478 4936 276534 4992
rect 278686 4936 278742 4992
rect 438214 644952 438270 645008
rect 438306 643184 438362 643240
rect 438398 641960 438454 642016
rect 438490 640328 438546 640384
rect 438582 639240 438638 639296
rect 438674 637608 438730 637664
rect 518898 589328 518954 589384
rect 518898 587696 518954 587752
rect 438766 579672 438822 579728
rect 443090 558864 443146 558920
rect 445758 558864 445814 558920
rect 447598 558864 447654 558920
rect 453670 558864 453726 558920
rect 454682 558864 454738 558920
rect 455970 558864 456026 558920
rect 457350 558864 457406 558920
rect 458270 558864 458326 558920
rect 460846 558864 460902 558920
rect 461674 558864 461730 558920
rect 462594 558864 462650 558920
rect 464250 558864 464306 558920
rect 465262 558864 465318 558920
rect 466458 558864 466514 558920
rect 467838 558864 467894 558920
rect 468666 558864 468722 558920
rect 469218 558864 469274 558920
rect 470598 558864 470654 558920
rect 471978 558864 472034 558920
rect 473358 558864 473414 558920
rect 474830 558864 474886 558920
rect 475474 558864 475530 558920
rect 477130 558864 477186 558920
rect 478234 558864 478290 558920
rect 478970 558864 479026 558920
rect 480534 558884 480590 558920
rect 480534 558864 480536 558884
rect 480536 558864 480588 558884
rect 480588 558864 480590 558884
rect 452658 558728 452714 558784
rect 449898 558456 449954 558512
rect 453302 558592 453358 558648
rect 453946 558592 454002 558648
rect 451278 558068 451334 558104
rect 451278 558048 451280 558068
rect 451280 558048 451332 558068
rect 451332 558048 451334 558068
rect 452658 557504 452714 557560
rect 453394 557504 453450 557560
rect 459650 558592 459706 558648
rect 462962 558612 463018 558648
rect 462962 558592 462964 558612
rect 462964 558592 463016 558612
rect 463016 558592 463018 558612
rect 461030 557640 461086 557696
rect 455418 557504 455474 557560
rect 456798 557504 456854 557560
rect 458178 557504 458234 557560
rect 459558 557504 459614 557560
rect 460938 557504 460994 557560
rect 462318 557504 462374 557560
rect 463698 557504 463754 557560
rect 465078 557504 465134 557560
rect 466550 558764 466552 558784
rect 466552 558764 466604 558784
rect 466604 558764 466606 558784
rect 466550 558728 466606 558764
rect 467930 558728 467986 558784
rect 468022 558592 468078 558648
rect 470046 558728 470102 558784
rect 471334 558728 471390 558784
rect 472162 558748 472218 558784
rect 472162 558728 472164 558748
rect 472164 558728 472216 558748
rect 472216 558728 472218 558748
rect 473450 558592 473506 558648
rect 476118 558456 476174 558512
rect 476210 558320 476266 558376
rect 477498 558340 477554 558376
rect 477498 558320 477500 558340
rect 477500 558320 477552 558340
rect 477552 558320 477554 558340
rect 478878 558204 478934 558240
rect 483018 558864 483074 558920
rect 480350 558728 480406 558784
rect 481638 558748 481694 558784
rect 481638 558728 481640 558748
rect 481640 558728 481692 558748
rect 481692 558728 481694 558748
rect 484398 558612 484454 558648
rect 484398 558592 484400 558612
rect 484400 558592 484452 558612
rect 484452 558592 484454 558612
rect 488538 558592 488594 558648
rect 481638 558456 481694 558512
rect 485778 558456 485834 558512
rect 487158 558456 487214 558512
rect 478878 558184 478880 558204
rect 478880 558184 478932 558204
rect 478932 558184 478934 558204
rect 483018 558184 483074 558240
rect 484398 558184 484454 558240
rect 485778 558184 485834 558240
rect 483110 558048 483166 558104
rect 483018 557640 483074 557696
rect 488538 558048 488594 558104
rect 487158 557912 487214 557968
rect 474646 557540 474648 557560
rect 474648 557540 474700 557560
rect 474700 557540 474702 557560
rect 474646 557504 474702 557540
rect 476394 557540 476396 557560
rect 476396 557540 476448 557560
rect 476448 557540 476450 557560
rect 476394 557504 476450 557540
rect 513378 412684 513434 412720
rect 513378 412664 513380 412684
rect 513380 412664 513432 412684
rect 513432 412664 513434 412684
rect 313278 318724 313280 318744
rect 313280 318724 313332 318744
rect 313332 318724 313334 318744
rect 279698 318280 279754 318336
rect 279974 8880 280030 8936
rect 280066 4800 280122 4856
rect 283654 5480 283710 5536
rect 290738 5344 290794 5400
rect 313278 318688 313334 318724
rect 443090 318724 443092 318744
rect 443092 318724 443144 318744
rect 443144 318724 443146 318744
rect 443090 318688 443146 318724
rect 296074 3168 296130 3224
rect 314566 3304 314622 3360
rect 321650 3304 321706 3360
rect 321834 3304 321890 3360
rect 321834 3032 321890 3088
rect 347870 5208 347926 5264
rect 362130 6704 362186 6760
rect 365810 6568 365866 6624
rect 372802 6432 372858 6488
rect 380898 10784 380954 10840
rect 379978 6296 380034 6352
rect 383658 10648 383714 10704
rect 387062 6160 387118 6216
rect 390650 10512 390706 10568
rect 394698 10376 394754 10432
rect 398838 10240 398894 10296
rect 435822 3168 435878 3224
rect 450174 3984 450230 4040
rect 457258 3848 457314 3904
rect 465630 8200 465686 8256
rect 464434 3712 464490 3768
rect 469126 8064 469182 8120
rect 472714 7928 472770 7984
rect 471518 3576 471574 3632
rect 476302 7792 476358 7848
rect 479890 7656 479946 7712
rect 478694 3440 478750 3496
rect 484582 7520 484638 7576
rect 485870 12144 485926 12200
rect 488538 12008 488594 12064
rect 492678 11872 492734 11928
rect 495438 11736 495494 11792
rect 499578 11600 499634 11656
rect 502338 15000 502394 15056
rect 506478 14864 506534 14920
rect 510618 14728 510674 14784
rect 513378 14592 513434 14648
rect 545118 14456 545174 14512
rect 531042 9560 531098 9616
rect 538126 9424 538182 9480
rect 546498 13504 546554 13560
rect 549258 13368 549314 13424
rect 548890 9288 548946 9344
rect 553398 13232 553454 13288
rect 556158 13096 556214 13152
rect 555974 9152 556030 9208
rect 560298 12960 560354 13016
rect 570234 9016 570290 9072
rect 572626 5072 572682 5128
rect 576214 4936 576270 4992
rect 580998 8880 581054 8936
rect 579802 4800 579858 4856
rect 582194 3304 582250 3360
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 583520 686204 584960 686444
rect -960 682124 480 682364
rect 583520 674508 584960 674748
rect -960 667844 480 668084
rect 583520 662676 584960 662916
rect -960 653428 480 653668
rect 129273 652900 129339 652901
rect 133689 652900 133755 652901
rect 259177 652900 259243 652901
rect 263593 652900 263659 652901
rect 129222 652898 129228 652900
rect 129182 652838 129228 652898
rect 129292 652896 129339 652900
rect 133638 652898 133644 652900
rect 129334 652840 129339 652896
rect 129222 652836 129228 652838
rect 129292 652836 129339 652840
rect 133598 652838 133644 652898
rect 133708 652896 133755 652900
rect 259126 652898 259132 652900
rect 133750 652840 133755 652896
rect 133638 652836 133644 652838
rect 133708 652836 133755 652840
rect 259086 652838 259132 652898
rect 259196 652896 259243 652900
rect 259238 652840 259243 652896
rect 259126 652836 259132 652838
rect 259196 652836 259243 652840
rect 263542 652836 263548 652900
rect 263612 652898 263659 652900
rect 378133 652900 378199 652901
rect 383561 652900 383627 652901
rect 263612 652896 263704 652898
rect 263654 652840 263704 652896
rect 263612 652838 263704 652840
rect 378133 652896 378180 652900
rect 378244 652898 378250 652900
rect 383510 652898 383516 652900
rect 378133 652840 378138 652896
rect 263612 652836 263659 652838
rect 129273 652835 129339 652836
rect 133689 652835 133755 652836
rect 259177 652835 259243 652836
rect 263593 652835 263659 652836
rect 378133 652836 378180 652840
rect 378244 652838 378290 652898
rect 383470 652838 383516 652898
rect 383580 652896 383627 652900
rect 383622 652840 383627 652896
rect 378244 652836 378250 652838
rect 383510 652836 383516 652838
rect 383580 652836 383627 652840
rect 378133 652835 378199 652836
rect 383561 652835 383627 652836
rect 508405 652900 508471 652901
rect 513373 652900 513439 652901
rect 508405 652896 508452 652900
rect 508516 652898 508522 652900
rect 508405 652840 508410 652896
rect 508405 652836 508452 652840
rect 508516 652838 508562 652898
rect 513373 652896 513420 652900
rect 513484 652898 513490 652900
rect 513373 652840 513378 652896
rect 508516 652836 508522 652838
rect 513373 652836 513420 652840
rect 513484 652838 513530 652898
rect 513484 652836 513490 652838
rect 508405 652835 508471 652836
rect 513373 652835 513439 652836
rect 583520 650980 584960 651220
rect 266445 649906 266511 649909
rect 387149 649906 387215 649909
rect 516409 649906 516475 649909
rect 266445 649904 266554 649906
rect 266445 649848 266450 649904
rect 266506 649848 266554 649904
rect 266445 649843 266554 649848
rect 387149 649904 387258 649906
rect 387149 649848 387154 649904
rect 387210 649848 387258 649904
rect 387149 649843 387258 649848
rect 516409 649904 516610 649906
rect 516409 649848 516414 649904
rect 516470 649848 516610 649904
rect 516409 649846 516610 649848
rect 516409 649843 516475 649846
rect 137645 649713 137711 649716
rect 137172 649711 137711 649713
rect 137172 649655 137650 649711
rect 137706 649655 137711 649711
rect 266494 649683 266554 649843
rect 387198 649683 387258 649843
rect 516550 649683 516610 649846
rect 137172 649653 137711 649655
rect 137645 649650 137711 649653
rect 282269 648684 282335 648685
rect 282269 648680 282316 648684
rect 282380 648682 282386 648684
rect 282269 648624 282274 648680
rect 282269 648620 282316 648624
rect 282380 648622 282426 648682
rect 282380 648620 282386 648622
rect 282269 648619 282335 648620
rect 57881 646098 57947 646101
rect 60046 646098 60106 646587
rect 57881 646096 60106 646098
rect 57881 646040 57886 646096
rect 57942 646040 60106 646096
rect 57881 646038 60106 646040
rect 188337 646098 188403 646101
rect 190134 646098 190194 646587
rect 188337 646096 190194 646098
rect 188337 646040 188342 646096
rect 188398 646040 190194 646096
rect 188337 646038 190194 646040
rect 307385 646098 307451 646101
rect 310102 646098 310162 646587
rect 307385 646096 310162 646098
rect 307385 646040 307390 646096
rect 307446 646040 310162 646096
rect 307385 646038 310162 646040
rect 438117 646098 438183 646101
rect 440006 646098 440066 646587
rect 438117 646096 440066 646098
rect 438117 646040 438122 646096
rect 438178 646040 440066 646096
rect 438117 646038 440066 646040
rect 57881 646035 57947 646038
rect 188337 646035 188403 646038
rect 307385 646035 307451 646038
rect 438117 646035 438183 646038
rect 57789 645010 57855 645013
rect 60046 645010 60106 645459
rect 57789 645008 60106 645010
rect 57789 644952 57794 645008
rect 57850 644952 60106 645008
rect 57789 644950 60106 644952
rect 188429 645010 188495 645013
rect 190134 645010 190194 645459
rect 188429 645008 190194 645010
rect 188429 644952 188434 645008
rect 188490 644952 190194 645008
rect 188429 644950 190194 644952
rect 307109 645010 307175 645013
rect 310102 645010 310162 645459
rect 307109 645008 310162 645010
rect 307109 644952 307114 645008
rect 307170 644952 310162 645008
rect 307109 644950 310162 644952
rect 438209 645010 438275 645013
rect 440006 645010 440066 645459
rect 438209 645008 440066 645010
rect 438209 644952 438214 645008
rect 438270 644952 440066 645008
rect 438209 644950 440066 644952
rect 57789 644947 57855 644950
rect 188429 644947 188495 644950
rect 307109 644947 307175 644950
rect 438209 644947 438275 644950
rect 57697 643242 57763 643245
rect 60046 643242 60106 643759
rect 57697 643240 60106 643242
rect 57697 643184 57702 643240
rect 57758 643184 60106 643240
rect 57697 643182 60106 643184
rect 188521 643242 188587 643245
rect 190134 643242 190194 643759
rect 307109 643514 307175 643517
rect 310102 643514 310162 643759
rect 307109 643512 310162 643514
rect 307109 643456 307114 643512
rect 307170 643456 310162 643512
rect 307109 643454 310162 643456
rect 307109 643451 307175 643454
rect 188521 643240 190194 643242
rect 188521 643184 188526 643240
rect 188582 643184 190194 643240
rect 188521 643182 190194 643184
rect 438301 643242 438367 643245
rect 440006 643242 440066 643759
rect 438301 643240 440066 643242
rect 438301 643184 438306 643240
rect 438362 643184 440066 643240
rect 438301 643182 440066 643184
rect 57697 643179 57763 643182
rect 188521 643179 188587 643182
rect 438301 643179 438367 643182
rect 57605 642018 57671 642021
rect 60046 642018 60106 642631
rect 57605 642016 60106 642018
rect 57605 641960 57610 642016
rect 57666 641960 60106 642016
rect 57605 641958 60106 641960
rect 188613 642018 188679 642021
rect 190134 642018 190194 642631
rect 307661 642154 307727 642157
rect 310102 642154 310162 642631
rect 307661 642152 310162 642154
rect 307661 642096 307666 642152
rect 307722 642096 310162 642152
rect 307661 642094 310162 642096
rect 307661 642091 307727 642094
rect 188613 642016 190194 642018
rect 188613 641960 188618 642016
rect 188674 641960 190194 642016
rect 188613 641958 190194 641960
rect 438393 642018 438459 642021
rect 440006 642018 440066 642631
rect 438393 642016 440066 642018
rect 438393 641960 438398 642016
rect 438454 641960 440066 642016
rect 438393 641958 440066 641960
rect 57605 641955 57671 641958
rect 188613 641955 188679 641958
rect 438393 641955 438459 641958
rect 57513 640386 57579 640389
rect 60046 640386 60106 640931
rect 57513 640384 60106 640386
rect 57513 640328 57518 640384
rect 57574 640328 60106 640384
rect 57513 640326 60106 640328
rect 188705 640386 188771 640389
rect 190134 640386 190194 640931
rect 307661 640522 307727 640525
rect 310102 640522 310162 640931
rect 307661 640520 310162 640522
rect 307661 640464 307666 640520
rect 307722 640464 310162 640520
rect 307661 640462 310162 640464
rect 307661 640459 307727 640462
rect 188705 640384 190194 640386
rect 188705 640328 188710 640384
rect 188766 640328 190194 640384
rect 188705 640326 190194 640328
rect 438485 640386 438551 640389
rect 440006 640386 440066 640931
rect 438485 640384 440066 640386
rect 438485 640328 438490 640384
rect 438546 640328 440066 640384
rect 438485 640326 440066 640328
rect 57513 640323 57579 640326
rect 188705 640323 188771 640326
rect 438485 640323 438551 640326
rect 57421 639298 57487 639301
rect 60046 639298 60106 639803
rect 57421 639296 60106 639298
rect -960 639012 480 639252
rect 57421 639240 57426 639296
rect 57482 639240 60106 639296
rect 57421 639238 60106 639240
rect 188797 639298 188863 639301
rect 190134 639298 190194 639803
rect 306649 639434 306715 639437
rect 310102 639434 310162 639803
rect 306649 639432 310162 639434
rect 306649 639376 306654 639432
rect 306710 639376 310162 639432
rect 306649 639374 310162 639376
rect 306649 639371 306715 639374
rect 188797 639296 190194 639298
rect 188797 639240 188802 639296
rect 188858 639240 190194 639296
rect 188797 639238 190194 639240
rect 438577 639298 438643 639301
rect 440006 639298 440066 639803
rect 438577 639296 440066 639298
rect 438577 639240 438582 639296
rect 438638 639240 440066 639296
rect 583520 639284 584960 639524
rect 438577 639238 440066 639240
rect 57421 639235 57487 639238
rect 188797 639235 188863 639238
rect 438577 639235 438643 639238
rect 57329 637666 57395 637669
rect 60046 637666 60106 638103
rect 57329 637664 60106 637666
rect 57329 637608 57334 637664
rect 57390 637608 60106 637664
rect 57329 637606 60106 637608
rect 188889 637666 188955 637669
rect 190134 637666 190194 638103
rect 306833 637938 306899 637941
rect 310102 637938 310162 638103
rect 306833 637936 310162 637938
rect 306833 637880 306838 637936
rect 306894 637880 310162 637936
rect 306833 637878 310162 637880
rect 306833 637875 306899 637878
rect 188889 637664 190194 637666
rect 188889 637608 188894 637664
rect 188950 637608 190194 637664
rect 188889 637606 190194 637608
rect 438669 637666 438735 637669
rect 440006 637666 440066 638103
rect 438669 637664 440066 637666
rect 438669 637608 438674 637664
rect 438730 637608 440066 637664
rect 438669 637606 440066 637608
rect 57329 637603 57395 637606
rect 188889 637603 188955 637606
rect 438669 637603 438735 637606
rect 583520 627588 584960 627828
rect -960 624732 480 624972
rect 583520 615756 584960 615996
rect -960 610316 480 610556
rect 583520 604060 584960 604300
rect -960 595900 480 596140
rect 583520 592364 584960 592604
rect 139393 589658 139459 589661
rect 136958 589656 139459 589658
rect 136958 589600 139398 589656
rect 139454 589600 139459 589656
rect 136958 589598 139459 589600
rect 136958 586614 137018 589598
rect 139393 589595 139459 589598
rect 267046 586666 267106 589412
rect 282177 587210 282243 587213
rect 282678 587210 282684 587212
rect 282177 587208 282684 587210
rect 282177 587152 282182 587208
rect 282238 587152 282684 587208
rect 282177 587150 282684 587152
rect 282177 587147 282243 587150
rect 282678 587148 282684 587150
rect 282748 587148 282754 587212
rect 387198 587210 387258 589412
rect 517102 589386 517162 589412
rect 518893 589386 518959 589389
rect 517102 589384 518959 589386
rect 517102 589328 518898 589384
rect 518954 589328 518959 589384
rect 517102 589326 518959 589328
rect 518893 589323 518959 589326
rect 518893 587754 518959 587757
rect 517102 587752 518959 587754
rect 517102 587696 518898 587752
rect 518954 587696 518959 587752
rect 517102 587694 518959 587696
rect 387558 587210 387564 587212
rect 387198 587150 387564 587210
rect 267046 586614 267290 586666
rect 136958 586584 137172 586614
rect 267046 586606 267658 586614
rect 136988 586554 137202 586584
rect -960 581620 480 581860
rect 137142 580410 137202 586554
rect 267046 583786 267106 586606
rect 267230 586584 267658 586606
rect 267260 586554 267658 586584
rect 267598 586530 267658 586554
rect 282177 586530 282243 586533
rect 267598 586528 282243 586530
rect 267598 586472 282182 586528
rect 282238 586472 282243 586528
rect 267598 586470 282243 586472
rect 282177 586467 282243 586470
rect 267046 583756 267260 583786
rect 267076 583726 267290 583756
rect 267230 580954 267290 583726
rect 269062 580954 269068 580956
rect 267230 580894 269068 580954
rect 269062 580892 269068 580894
rect 269132 580892 269138 580956
rect 387198 580954 387258 587150
rect 387558 587148 387564 587150
rect 387628 587148 387634 587212
rect 389173 580954 389239 580957
rect 387198 580952 389239 580954
rect 387198 580896 389178 580952
rect 389234 580896 389239 580952
rect 387198 580894 389239 580896
rect 517102 580954 517162 587694
rect 518893 587691 518959 587694
rect 518934 580954 518940 580956
rect 517102 580894 518940 580954
rect 389173 580891 389239 580894
rect 518934 580892 518940 580894
rect 519004 580892 519010 580956
rect 583520 580668 584960 580908
rect 137502 580410 137508 580412
rect 137142 580350 137508 580410
rect 137502 580348 137508 580350
rect 137572 580410 137578 580412
rect 139393 580410 139459 580413
rect 137572 580408 139459 580410
rect 137572 580352 139398 580408
rect 139454 580352 139459 580408
rect 137572 580350 139459 580352
rect 137572 580348 137578 580350
rect 139393 580347 139459 580350
rect 57237 579730 57303 579733
rect 60046 579730 60106 580255
rect 57237 579728 60106 579730
rect 57237 579672 57242 579728
rect 57298 579672 60106 579728
rect 57237 579670 60106 579672
rect 188981 579730 189047 579733
rect 190134 579730 190194 580255
rect 306925 580002 306991 580005
rect 310102 580002 310162 580255
rect 306925 580000 310162 580002
rect 306925 579944 306930 580000
rect 306986 579944 310162 580000
rect 306925 579942 310162 579944
rect 306925 579939 306991 579942
rect 188981 579728 190194 579730
rect 188981 579672 188986 579728
rect 189042 579672 190194 579728
rect 188981 579670 190194 579672
rect 438761 579730 438827 579733
rect 440006 579730 440066 580255
rect 438761 579728 440066 579730
rect 438761 579672 438766 579728
rect 438822 579672 440066 579728
rect 438761 579670 440066 579672
rect 57237 579667 57303 579670
rect 188981 579667 189047 579670
rect 438761 579667 438827 579670
rect 437841 579186 437907 579189
rect 439998 579186 440004 579188
rect 437841 579184 440004 579186
rect 437841 579128 437846 579184
rect 437902 579128 440004 579184
rect 437841 579126 440004 579128
rect 437841 579123 437907 579126
rect 439998 579124 440004 579126
rect 440068 579124 440074 579188
rect 60590 578988 60596 579052
rect 60660 578988 60666 579052
rect 187693 579050 187759 579053
rect 190126 579050 190132 579052
rect 187693 579048 190132 579050
rect 187693 578992 187698 579048
rect 187754 578992 190132 579048
rect 187693 578990 190132 578992
rect 60598 578555 60658 578988
rect 187693 578987 187759 578990
rect 190126 578988 190132 578990
rect 190196 578988 190202 579052
rect 190134 578555 190194 578988
rect 307661 578914 307727 578917
rect 307661 578912 310162 578914
rect 307661 578856 307666 578912
rect 307722 578856 310162 578912
rect 307661 578854 310162 578856
rect 307661 578851 307727 578854
rect 310102 578555 310162 578854
rect 440006 578555 440066 579124
rect 583520 568836 584960 569076
rect -960 567204 480 567444
rect 229369 560012 229435 560013
rect 229318 560010 229324 560012
rect 229278 559950 229324 560010
rect 229388 560008 229435 560012
rect 229430 559952 229435 560008
rect 229318 559948 229324 559950
rect 229388 559948 229435 559952
rect 229369 559947 229435 559948
rect 225822 559812 225828 559876
rect 225892 559874 225898 559876
rect 225965 559874 226031 559877
rect 225892 559872 226031 559874
rect 225892 559816 225970 559872
rect 226026 559816 226031 559872
rect 225892 559814 226031 559816
rect 225892 559812 225898 559814
rect 225965 559811 226031 559814
rect 227110 559268 227116 559332
rect 227180 559330 227186 559332
rect 227253 559330 227319 559333
rect 227180 559328 227319 559330
rect 227180 559272 227258 559328
rect 227314 559272 227319 559328
rect 227180 559270 227319 559272
rect 227180 559268 227186 559270
rect 227253 559267 227319 559270
rect 348417 559330 348483 559333
rect 351862 559330 351868 559332
rect 348417 559328 351868 559330
rect 348417 559272 348422 559328
rect 348478 559272 351868 559328
rect 348417 559270 351868 559272
rect 348417 559267 348483 559270
rect 351862 559268 351868 559270
rect 351932 559268 351938 559332
rect 357709 559330 357775 559333
rect 358854 559330 358860 559332
rect 357709 559328 358860 559330
rect 357709 559272 357714 559328
rect 357770 559272 358860 559328
rect 357709 559270 358860 559272
rect 357709 559267 357775 559270
rect 358854 559268 358860 559270
rect 358924 559268 358930 559332
rect 67398 558860 67404 558924
rect 67468 558922 67474 558924
rect 67541 558922 67607 558925
rect 67468 558920 67607 558922
rect 67468 558864 67546 558920
rect 67602 558864 67607 558920
rect 67468 558862 67607 558864
rect 67468 558860 67474 558862
rect 67541 558859 67607 558862
rect 68502 558860 68508 558924
rect 68572 558922 68578 558924
rect 68921 558922 68987 558925
rect 70209 558924 70275 558925
rect 71681 558924 71747 558925
rect 68572 558920 68987 558922
rect 68572 558864 68926 558920
rect 68982 558864 68987 558920
rect 68572 558862 68987 558864
rect 68572 558860 68578 558862
rect 68921 558859 68987 558862
rect 70158 558860 70164 558924
rect 70228 558922 70275 558924
rect 70228 558920 70320 558922
rect 70270 558864 70320 558920
rect 70228 558862 70320 558864
rect 70228 558860 70275 558862
rect 71630 558860 71636 558924
rect 71700 558922 71747 558924
rect 71700 558920 71792 558922
rect 71742 558864 71792 558920
rect 71700 558862 71792 558864
rect 71700 558860 71747 558862
rect 72366 558860 72372 558924
rect 72436 558922 72442 558924
rect 72509 558922 72575 558925
rect 72436 558920 72575 558922
rect 72436 558864 72514 558920
rect 72570 558864 72575 558920
rect 72436 558862 72575 558864
rect 72436 558860 72442 558862
rect 70209 558859 70275 558860
rect 71681 558859 71747 558860
rect 72509 558859 72575 558862
rect 72918 558860 72924 558924
rect 72988 558922 72994 558924
rect 73061 558922 73127 558925
rect 73705 558924 73771 558925
rect 74257 558924 74323 558925
rect 74993 558924 75059 558925
rect 73654 558922 73660 558924
rect 72988 558920 73127 558922
rect 72988 558864 73066 558920
rect 73122 558864 73127 558920
rect 72988 558862 73127 558864
rect 73614 558862 73660 558922
rect 73724 558920 73771 558924
rect 74206 558922 74212 558924
rect 73766 558864 73771 558920
rect 72988 558860 72994 558862
rect 73061 558859 73127 558862
rect 73654 558860 73660 558862
rect 73724 558860 73771 558864
rect 74166 558862 74212 558922
rect 74276 558920 74323 558924
rect 74942 558922 74948 558924
rect 74318 558864 74323 558920
rect 74206 558860 74212 558862
rect 74276 558860 74323 558864
rect 74902 558862 74948 558922
rect 75012 558920 75059 558924
rect 75054 558864 75059 558920
rect 74942 558860 74948 558862
rect 75012 558860 75059 558864
rect 75678 558860 75684 558924
rect 75748 558922 75754 558924
rect 75821 558922 75887 558925
rect 76833 558924 76899 558925
rect 77385 558924 77451 558925
rect 76782 558922 76788 558924
rect 75748 558920 75887 558922
rect 75748 558864 75826 558920
rect 75882 558864 75887 558920
rect 75748 558862 75887 558864
rect 76742 558862 76788 558922
rect 76852 558920 76899 558924
rect 77334 558922 77340 558924
rect 76894 558864 76899 558920
rect 75748 558860 75754 558862
rect 73705 558859 73771 558860
rect 74257 558859 74323 558860
rect 74993 558859 75059 558860
rect 75821 558859 75887 558862
rect 76782 558860 76788 558862
rect 76852 558860 76899 558864
rect 77294 558862 77340 558922
rect 77404 558920 77451 558924
rect 77446 558864 77451 558920
rect 77334 558860 77340 558862
rect 77404 558860 77451 558864
rect 78070 558860 78076 558924
rect 78140 558922 78146 558924
rect 78581 558922 78647 558925
rect 78140 558920 78647 558922
rect 78140 558864 78586 558920
rect 78642 558864 78647 558920
rect 78140 558862 78647 558864
rect 78140 558860 78146 558862
rect 76833 558859 76899 558860
rect 77385 558859 77451 558860
rect 78581 558859 78647 558862
rect 79174 558860 79180 558924
rect 79244 558922 79250 558924
rect 79317 558922 79383 558925
rect 79961 558924 80027 558925
rect 79244 558920 79383 558922
rect 79244 558864 79322 558920
rect 79378 558864 79383 558920
rect 79244 558862 79383 558864
rect 79244 558860 79250 558862
rect 79317 558859 79383 558862
rect 79910 558860 79916 558924
rect 79980 558922 80027 558924
rect 79980 558920 80072 558922
rect 80022 558864 80072 558920
rect 79980 558862 80072 558864
rect 79980 558860 80027 558862
rect 80646 558860 80652 558924
rect 80716 558922 80722 558924
rect 80789 558922 80855 558925
rect 81249 558924 81315 558925
rect 81985 558924 82051 558925
rect 82721 558924 82787 558925
rect 83825 558924 83891 558925
rect 84193 558924 84259 558925
rect 81198 558922 81204 558924
rect 80716 558920 80855 558922
rect 80716 558864 80794 558920
rect 80850 558864 80855 558920
rect 80716 558862 80855 558864
rect 81158 558862 81204 558922
rect 81268 558920 81315 558924
rect 81934 558922 81940 558924
rect 81310 558864 81315 558920
rect 80716 558860 80722 558862
rect 79961 558859 80027 558860
rect 80789 558859 80855 558862
rect 81198 558860 81204 558862
rect 81268 558860 81315 558864
rect 81894 558862 81940 558922
rect 82004 558920 82051 558924
rect 82046 558864 82051 558920
rect 81934 558860 81940 558862
rect 82004 558860 82051 558864
rect 82670 558860 82676 558924
rect 82740 558922 82787 558924
rect 83774 558922 83780 558924
rect 82740 558920 82832 558922
rect 82782 558864 82832 558920
rect 82740 558862 82832 558864
rect 83734 558862 83780 558922
rect 83844 558920 83891 558924
rect 83886 558864 83891 558920
rect 82740 558860 82787 558862
rect 83774 558860 83780 558862
rect 83844 558860 83891 558864
rect 84142 558860 84148 558924
rect 84212 558922 84259 558924
rect 84212 558920 84304 558922
rect 84254 558864 84304 558920
rect 84212 558862 84304 558864
rect 84212 558860 84259 558862
rect 85062 558860 85068 558924
rect 85132 558922 85138 558924
rect 85481 558922 85547 558925
rect 86769 558924 86835 558925
rect 87873 558924 87939 558925
rect 88241 558924 88307 558925
rect 85132 558920 85547 558922
rect 85132 558864 85486 558920
rect 85542 558864 85547 558920
rect 85132 558862 85547 558864
rect 85132 558860 85138 558862
rect 81249 558859 81315 558860
rect 81985 558859 82051 558860
rect 82721 558859 82787 558860
rect 83825 558859 83891 558860
rect 84193 558859 84259 558860
rect 85481 558859 85547 558862
rect 86718 558860 86724 558924
rect 86788 558922 86835 558924
rect 87822 558922 87828 558924
rect 86788 558920 86880 558922
rect 86830 558864 86880 558920
rect 86788 558862 86880 558864
rect 87782 558862 87828 558922
rect 87892 558920 87939 558924
rect 87934 558864 87939 558920
rect 86788 558860 86835 558862
rect 87822 558860 87828 558862
rect 87892 558860 87939 558864
rect 88190 558860 88196 558924
rect 88260 558922 88307 558924
rect 88885 558924 88951 558925
rect 88260 558920 88352 558922
rect 88302 558864 88352 558920
rect 88260 558862 88352 558864
rect 88885 558920 88932 558924
rect 88996 558922 89002 558924
rect 88885 558864 88890 558920
rect 88260 558860 88307 558862
rect 86769 558859 86835 558860
rect 87873 558859 87939 558860
rect 88241 558859 88307 558860
rect 88885 558860 88932 558864
rect 88996 558862 89042 558922
rect 88996 558860 89002 558862
rect 89110 558860 89116 558924
rect 89180 558922 89186 558924
rect 89345 558922 89411 558925
rect 89180 558920 89411 558922
rect 89180 558864 89350 558920
rect 89406 558864 89411 558920
rect 89180 558862 89411 558864
rect 89180 558860 89186 558862
rect 88885 558859 88951 558860
rect 89345 558859 89411 558862
rect 89805 558924 89871 558925
rect 91001 558924 91067 558925
rect 89805 558920 89852 558924
rect 89916 558922 89922 558924
rect 89805 558864 89810 558920
rect 89805 558860 89852 558864
rect 89916 558862 89962 558922
rect 89916 558860 89922 558862
rect 90950 558860 90956 558924
rect 91020 558922 91067 558924
rect 91020 558920 91112 558922
rect 91062 558864 91112 558920
rect 91020 558862 91112 558864
rect 91020 558860 91067 558862
rect 92054 558860 92060 558924
rect 92124 558922 92130 558924
rect 92289 558922 92355 558925
rect 92473 558924 92539 558925
rect 92124 558920 92355 558922
rect 92124 558864 92294 558920
rect 92350 558864 92355 558920
rect 92124 558862 92355 558864
rect 92124 558860 92130 558862
rect 89805 558859 89871 558860
rect 91001 558859 91067 558860
rect 92289 558859 92355 558862
rect 92422 558860 92428 558924
rect 92492 558922 92539 558924
rect 92492 558920 92584 558922
rect 92534 558864 92584 558920
rect 92492 558862 92584 558864
rect 92492 558860 92539 558862
rect 93158 558860 93164 558924
rect 93228 558922 93234 558924
rect 93669 558922 93735 558925
rect 94865 558924 94931 558925
rect 95049 558924 95115 558925
rect 94814 558922 94820 558924
rect 93228 558920 93735 558922
rect 93228 558864 93674 558920
rect 93730 558864 93735 558920
rect 93228 558862 93735 558864
rect 94774 558862 94820 558922
rect 94884 558920 94931 558924
rect 94926 558864 94931 558920
rect 93228 558860 93234 558862
rect 92473 558859 92539 558860
rect 93669 558859 93735 558862
rect 94814 558860 94820 558862
rect 94884 558860 94931 558864
rect 94998 558860 95004 558924
rect 95068 558922 95115 558924
rect 95693 558924 95759 558925
rect 96521 558924 96587 558925
rect 97073 558924 97139 558925
rect 97625 558924 97691 558925
rect 95068 558920 95160 558922
rect 95110 558864 95160 558920
rect 95068 558862 95160 558864
rect 95693 558920 95740 558924
rect 95804 558922 95810 558924
rect 95693 558864 95698 558920
rect 95068 558860 95115 558862
rect 94865 558859 94931 558860
rect 95049 558859 95115 558860
rect 95693 558860 95740 558864
rect 95804 558862 95850 558922
rect 95804 558860 95810 558862
rect 96470 558860 96476 558924
rect 96540 558922 96587 558924
rect 97022 558922 97028 558924
rect 96540 558920 96632 558922
rect 96582 558864 96632 558920
rect 96540 558862 96632 558864
rect 96982 558862 97028 558922
rect 97092 558920 97139 558924
rect 97574 558922 97580 558924
rect 97134 558864 97139 558920
rect 96540 558860 96587 558862
rect 97022 558860 97028 558862
rect 97092 558860 97139 558864
rect 97534 558862 97580 558922
rect 97644 558920 97691 558924
rect 97686 558864 97691 558920
rect 97574 558860 97580 558862
rect 97644 558860 97691 558864
rect 98310 558860 98316 558924
rect 98380 558922 98386 558924
rect 98545 558922 98611 558925
rect 98380 558920 98611 558922
rect 98380 558864 98550 558920
rect 98606 558864 98611 558920
rect 98380 558862 98611 558864
rect 98380 558860 98386 558862
rect 95693 558859 95759 558860
rect 96521 558859 96587 558860
rect 97073 558859 97139 558860
rect 97625 558859 97691 558860
rect 98545 558859 98611 558862
rect 99046 558860 99052 558924
rect 99116 558922 99122 558924
rect 99281 558922 99347 558925
rect 99116 558920 99347 558922
rect 99116 558864 99286 558920
rect 99342 558864 99347 558920
rect 99116 558862 99347 558864
rect 99116 558860 99122 558862
rect 99281 558859 99347 558862
rect 100150 558860 100156 558924
rect 100220 558922 100226 558924
rect 100569 558922 100635 558925
rect 102041 558924 102107 558925
rect 104801 558924 104867 558925
rect 101990 558922 101996 558924
rect 100220 558920 100635 558922
rect 100220 558864 100574 558920
rect 100630 558864 100635 558920
rect 100220 558862 100635 558864
rect 101950 558862 101996 558922
rect 102060 558920 102107 558924
rect 104750 558922 104756 558924
rect 102102 558864 102107 558920
rect 100220 558860 100226 558862
rect 100569 558859 100635 558862
rect 101990 558860 101996 558862
rect 102060 558860 102107 558864
rect 104710 558862 104756 558922
rect 104820 558920 104867 558924
rect 104862 558864 104867 558920
rect 104750 558860 104756 558862
rect 104820 558860 104867 558864
rect 107142 558860 107148 558924
rect 107212 558922 107218 558924
rect 107469 558922 107535 558925
rect 108481 558924 108547 558925
rect 194409 558924 194475 558925
rect 108430 558922 108436 558924
rect 107212 558920 107535 558922
rect 107212 558864 107474 558920
rect 107530 558864 107535 558920
rect 107212 558862 107535 558864
rect 108390 558862 108436 558922
rect 108500 558920 108547 558924
rect 194358 558922 194364 558924
rect 108542 558864 108547 558920
rect 107212 558860 107218 558862
rect 102041 558859 102107 558860
rect 104801 558859 104867 558860
rect 107469 558859 107535 558862
rect 108430 558860 108436 558862
rect 108500 558860 108547 558864
rect 194318 558862 194364 558922
rect 194428 558920 194475 558924
rect 194470 558864 194475 558920
rect 194358 558860 194364 558862
rect 194428 558860 194475 558864
rect 108481 558859 108547 558860
rect 194409 558859 194475 558860
rect 195973 558922 196039 558925
rect 200205 558924 200271 558925
rect 201493 558924 201559 558925
rect 196198 558922 196204 558924
rect 195973 558920 196204 558922
rect 195973 558864 195978 558920
rect 196034 558864 196204 558920
rect 195973 558862 196204 558864
rect 195973 558859 196039 558862
rect 196198 558860 196204 558862
rect 196268 558860 196274 558924
rect 200205 558922 200252 558924
rect 200160 558920 200252 558922
rect 200160 558864 200210 558920
rect 200160 558862 200252 558864
rect 200205 558860 200252 558862
rect 200316 558860 200322 558924
rect 201493 558922 201540 558924
rect 201448 558920 201540 558922
rect 201448 558864 201498 558920
rect 201448 558862 201540 558864
rect 201493 558860 201540 558862
rect 201604 558860 201610 558924
rect 202638 558860 202644 558924
rect 202708 558922 202714 558924
rect 202781 558922 202847 558925
rect 203793 558924 203859 558925
rect 203742 558922 203748 558924
rect 202708 558920 202847 558922
rect 202708 558864 202786 558920
rect 202842 558864 202847 558920
rect 202708 558862 202847 558864
rect 203702 558862 203748 558922
rect 203812 558920 203859 558924
rect 203854 558864 203859 558920
rect 202708 558860 202714 558862
rect 200205 558859 200271 558860
rect 201493 558859 201559 558860
rect 202781 558859 202847 558862
rect 203742 558860 203748 558862
rect 203812 558860 203859 558864
rect 203926 558860 203932 558924
rect 203996 558922 204002 558924
rect 204161 558922 204227 558925
rect 203996 558920 204227 558922
rect 203996 558864 204166 558920
rect 204222 558864 204227 558920
rect 203996 558862 204227 558864
rect 203996 558860 204002 558862
rect 203793 558859 203859 558860
rect 204161 558859 204227 558862
rect 205398 558860 205404 558924
rect 205468 558922 205474 558924
rect 205541 558922 205607 558925
rect 205468 558920 205607 558922
rect 205468 558864 205546 558920
rect 205602 558864 205607 558920
rect 205468 558862 205607 558864
rect 205468 558860 205474 558862
rect 205541 558859 205607 558862
rect 206134 558860 206140 558924
rect 206204 558922 206210 558924
rect 206369 558922 206435 558925
rect 206204 558920 206435 558922
rect 206204 558864 206374 558920
rect 206430 558864 206435 558920
rect 206204 558862 206435 558864
rect 206204 558860 206210 558862
rect 206369 558859 206435 558862
rect 208342 558860 208348 558924
rect 208412 558922 208418 558924
rect 208485 558922 208551 558925
rect 211889 558924 211955 558925
rect 211838 558922 211844 558924
rect 208412 558920 208551 558922
rect 208412 558864 208490 558920
rect 208546 558864 208551 558920
rect 208412 558862 208551 558864
rect 211798 558862 211844 558922
rect 211908 558920 211955 558924
rect 211950 558864 211955 558920
rect 208412 558860 208418 558862
rect 208485 558859 208551 558862
rect 211838 558860 211844 558862
rect 211908 558860 211955 558864
rect 211889 558859 211955 558860
rect 213085 558924 213151 558925
rect 213085 558920 213132 558924
rect 213196 558922 213202 558924
rect 213913 558922 213979 558925
rect 215293 558924 215359 558925
rect 218789 558924 218855 558925
rect 220077 558924 220143 558925
rect 221089 558924 221155 558925
rect 214046 558922 214052 558924
rect 213085 558864 213090 558920
rect 213085 558860 213132 558864
rect 213196 558862 213242 558922
rect 213913 558920 214052 558922
rect 213913 558864 213918 558920
rect 213974 558864 214052 558920
rect 213913 558862 214052 558864
rect 213196 558860 213202 558862
rect 213085 558859 213151 558860
rect 213913 558859 213979 558862
rect 214046 558860 214052 558862
rect 214116 558860 214122 558924
rect 215293 558920 215340 558924
rect 215404 558922 215410 558924
rect 215293 558864 215298 558920
rect 215293 558860 215340 558864
rect 215404 558862 215450 558922
rect 218789 558920 218836 558924
rect 218900 558922 218906 558924
rect 218789 558864 218794 558920
rect 215404 558860 215410 558862
rect 218789 558860 218836 558864
rect 218900 558862 218946 558922
rect 220077 558920 220124 558924
rect 220188 558922 220194 558924
rect 221038 558922 221044 558924
rect 220077 558864 220082 558920
rect 218900 558860 218906 558862
rect 220077 558860 220124 558864
rect 220188 558862 220234 558922
rect 220998 558862 221044 558922
rect 221108 558920 221155 558924
rect 221150 558864 221155 558920
rect 220188 558860 220194 558862
rect 221038 558860 221044 558862
rect 221108 558860 221155 558864
rect 215293 558859 215359 558860
rect 218789 558859 218855 558860
rect 220077 558859 220143 558860
rect 221089 558859 221155 558860
rect 222285 558924 222351 558925
rect 223573 558924 223639 558925
rect 222285 558920 222332 558924
rect 222396 558922 222402 558924
rect 222285 558864 222290 558920
rect 222285 558860 222332 558864
rect 222396 558862 222442 558922
rect 223573 558920 223620 558924
rect 223684 558922 223690 558924
rect 223941 558922 224007 558925
rect 228081 558924 228147 558925
rect 224534 558922 224540 558924
rect 223573 558864 223578 558920
rect 222396 558860 222402 558862
rect 223573 558860 223620 558864
rect 223684 558862 223730 558922
rect 223941 558920 224540 558922
rect 223941 558864 223946 558920
rect 224002 558864 224540 558920
rect 223941 558862 224540 558864
rect 223684 558860 223690 558862
rect 222285 558859 222351 558860
rect 223573 558859 223639 558860
rect 223941 558859 224007 558862
rect 224534 558860 224540 558862
rect 224604 558860 224610 558924
rect 228030 558922 228036 558924
rect 227990 558862 228036 558922
rect 228100 558920 228147 558924
rect 228142 558864 228147 558920
rect 228030 558860 228036 558862
rect 228100 558860 228147 558864
rect 235758 558860 235764 558924
rect 235828 558922 235834 558924
rect 235901 558922 235967 558925
rect 237281 558924 237347 558925
rect 235828 558920 235967 558922
rect 235828 558864 235906 558920
rect 235962 558864 235967 558920
rect 235828 558862 235967 558864
rect 235828 558860 235834 558862
rect 228081 558859 228147 558860
rect 235901 558859 235967 558862
rect 237230 558860 237236 558924
rect 237300 558922 237347 558924
rect 237300 558920 237392 558922
rect 237342 558864 237392 558920
rect 237300 558862 237392 558864
rect 237300 558860 237347 558862
rect 239622 558860 239628 558924
rect 239692 558922 239698 558924
rect 240041 558922 240107 558925
rect 239692 558920 240107 558922
rect 239692 558864 240046 558920
rect 240102 558864 240107 558920
rect 239692 558862 240107 558864
rect 239692 558860 239698 558862
rect 237281 558859 237347 558860
rect 240041 558859 240107 558862
rect 313733 558924 313799 558925
rect 313733 558920 313780 558924
rect 313844 558922 313850 558924
rect 316033 558922 316099 558925
rect 317413 558924 317479 558925
rect 316166 558922 316172 558924
rect 313733 558864 313738 558920
rect 313733 558860 313780 558864
rect 313844 558862 313890 558922
rect 316033 558920 316172 558922
rect 316033 558864 316038 558920
rect 316094 558864 316172 558920
rect 316033 558862 316172 558864
rect 313844 558860 313850 558862
rect 313733 558859 313799 558860
rect 316033 558859 316099 558862
rect 316166 558860 316172 558862
rect 316236 558860 316242 558924
rect 317413 558922 317460 558924
rect 317368 558920 317460 558922
rect 317368 558864 317418 558920
rect 317368 558862 317460 558864
rect 317413 558860 317460 558862
rect 317524 558860 317530 558924
rect 320265 558922 320331 558925
rect 320950 558922 320956 558924
rect 320265 558920 320956 558922
rect 320265 558864 320270 558920
rect 320326 558864 320956 558920
rect 320265 558862 320956 558864
rect 317413 558859 317479 558860
rect 320265 558859 320331 558862
rect 320950 558860 320956 558862
rect 321020 558860 321026 558924
rect 322606 558860 322612 558924
rect 322676 558922 322682 558924
rect 322841 558922 322907 558925
rect 322676 558920 322907 558922
rect 322676 558864 322846 558920
rect 322902 558864 322907 558920
rect 322676 558862 322907 558864
rect 322676 558860 322682 558862
rect 322841 558859 322907 558862
rect 323485 558924 323551 558925
rect 328545 558924 328611 558925
rect 323485 558920 323532 558924
rect 323596 558922 323602 558924
rect 328494 558922 328500 558924
rect 323485 558864 323490 558920
rect 323485 558860 323532 558864
rect 323596 558862 323642 558922
rect 328454 558862 328500 558922
rect 328564 558920 328611 558924
rect 328606 558864 328611 558920
rect 323596 558860 323602 558862
rect 328494 558860 328500 558862
rect 328564 558860 328611 558864
rect 323485 558859 323551 558860
rect 328545 558859 328611 558860
rect 329557 558924 329623 558925
rect 330477 558924 330543 558925
rect 329557 558920 329604 558924
rect 329668 558922 329674 558924
rect 329557 558864 329562 558920
rect 329557 558860 329604 558864
rect 329668 558862 329714 558922
rect 330477 558920 330524 558924
rect 330588 558922 330594 558924
rect 330477 558864 330482 558920
rect 329668 558860 329674 558862
rect 330477 558860 330524 558864
rect 330588 558862 330634 558922
rect 330588 558860 330594 558862
rect 331806 558860 331812 558924
rect 331876 558922 331882 558924
rect 332501 558922 332567 558925
rect 333145 558924 333211 558925
rect 333094 558922 333100 558924
rect 331876 558920 332567 558922
rect 331876 558864 332506 558920
rect 332562 558864 332567 558920
rect 331876 558862 332567 558864
rect 333054 558862 333100 558922
rect 333164 558920 333211 558924
rect 333206 558864 333211 558920
rect 331876 558860 331882 558862
rect 329557 558859 329623 558860
rect 330477 558859 330543 558860
rect 332501 558859 332567 558862
rect 333094 558860 333100 558862
rect 333164 558860 333211 558864
rect 334014 558860 334020 558924
rect 334084 558922 334090 558924
rect 334249 558922 334315 558925
rect 334084 558920 334315 558922
rect 334084 558864 334254 558920
rect 334310 558864 334315 558920
rect 334084 558862 334315 558864
rect 334084 558860 334090 558862
rect 333145 558859 333211 558860
rect 334249 558859 334315 558862
rect 335486 558860 335492 558924
rect 335556 558922 335562 558924
rect 335905 558922 335971 558925
rect 335556 558920 335971 558922
rect 335556 558864 335910 558920
rect 335966 558864 335971 558920
rect 335556 558862 335971 558864
rect 335556 558860 335562 558862
rect 335905 558859 335971 558862
rect 336273 558922 336339 558925
rect 337745 558924 337811 558925
rect 339033 558924 339099 558925
rect 336406 558922 336412 558924
rect 336273 558920 336412 558922
rect 336273 558864 336278 558920
rect 336334 558864 336412 558920
rect 336273 558862 336412 558864
rect 336273 558859 336339 558862
rect 336406 558860 336412 558862
rect 336476 558860 336482 558924
rect 337694 558922 337700 558924
rect 337654 558862 337700 558922
rect 337764 558920 337811 558924
rect 338982 558922 338988 558924
rect 337806 558864 337811 558920
rect 337694 558860 337700 558862
rect 337764 558860 337811 558864
rect 338942 558862 338988 558922
rect 339052 558920 339099 558924
rect 339094 558864 339099 558920
rect 338982 558860 338988 558862
rect 339052 558860 339099 558864
rect 337745 558859 337811 558860
rect 339033 558859 339099 558860
rect 339861 558924 339927 558925
rect 341241 558924 341307 558925
rect 342529 558924 342595 558925
rect 343633 558924 343699 558925
rect 339861 558920 339908 558924
rect 339972 558922 339978 558924
rect 341190 558922 341196 558924
rect 339861 558864 339866 558920
rect 339861 558860 339908 558864
rect 339972 558862 340018 558922
rect 341150 558862 341196 558922
rect 341260 558920 341307 558924
rect 342478 558922 342484 558924
rect 341302 558864 341307 558920
rect 339972 558860 339978 558862
rect 341190 558860 341196 558862
rect 341260 558860 341307 558864
rect 342438 558862 342484 558922
rect 342548 558920 342595 558924
rect 343582 558922 343588 558924
rect 342590 558864 342595 558920
rect 342478 558860 342484 558862
rect 342548 558860 342595 558864
rect 343542 558862 343588 558922
rect 343652 558920 343699 558924
rect 343694 558864 343699 558920
rect 343582 558860 343588 558862
rect 343652 558860 343699 558864
rect 344686 558860 344692 558924
rect 344756 558922 344762 558924
rect 344829 558922 344895 558925
rect 344756 558920 344895 558922
rect 344756 558864 344834 558920
rect 344890 558864 344895 558920
rect 344756 558862 344895 558864
rect 344756 558860 344762 558862
rect 339861 558859 339927 558860
rect 341241 558859 341307 558860
rect 342529 558859 342595 558860
rect 343633 558859 343699 558860
rect 344829 558859 344895 558862
rect 345749 558924 345815 558925
rect 346485 558924 346551 558925
rect 348233 558924 348299 558925
rect 345749 558920 345796 558924
rect 345860 558922 345866 558924
rect 345749 558864 345754 558920
rect 345749 558860 345796 558864
rect 345860 558862 345906 558922
rect 346485 558920 346532 558924
rect 346596 558922 346602 558924
rect 348182 558922 348188 558924
rect 346485 558864 346490 558920
rect 345860 558860 345866 558862
rect 346485 558860 346532 558864
rect 346596 558862 346642 558922
rect 348142 558862 348188 558922
rect 348252 558920 348299 558924
rect 348294 558864 348299 558920
rect 346596 558860 346602 558862
rect 348182 558860 348188 558862
rect 348252 558860 348299 558864
rect 345749 558859 345815 558860
rect 346485 558859 346551 558860
rect 348233 558859 348299 558860
rect 349337 558922 349403 558925
rect 350533 558924 350599 558925
rect 349470 558922 349476 558924
rect 349337 558920 349476 558922
rect 349337 558864 349342 558920
rect 349398 558864 349476 558920
rect 349337 558862 349476 558864
rect 349337 558859 349403 558862
rect 349470 558860 349476 558862
rect 349540 558860 349546 558924
rect 350533 558920 350580 558924
rect 350644 558922 350650 558924
rect 352005 558922 352071 558925
rect 352414 558922 352420 558924
rect 350533 558864 350538 558920
rect 350533 558860 350580 558864
rect 350644 558862 350690 558922
rect 352005 558920 352420 558922
rect 352005 558864 352010 558920
rect 352066 558864 352420 558920
rect 352005 558862 352420 558864
rect 350644 558860 350650 558862
rect 350533 558859 350599 558860
rect 352005 558859 352071 558862
rect 352414 558860 352420 558862
rect 352484 558860 352490 558924
rect 353293 558922 353359 558925
rect 443085 558924 443151 558925
rect 353518 558922 353524 558924
rect 353293 558920 353524 558922
rect 353293 558864 353298 558920
rect 353354 558864 353524 558920
rect 353293 558862 353524 558864
rect 353293 558859 353359 558862
rect 353518 558860 353524 558862
rect 353588 558860 353594 558924
rect 443085 558920 443132 558924
rect 443196 558922 443202 558924
rect 445753 558922 445819 558925
rect 446254 558922 446260 558924
rect 443085 558864 443090 558920
rect 443085 558860 443132 558864
rect 443196 558862 443242 558922
rect 445753 558920 446260 558922
rect 445753 558864 445758 558920
rect 445814 558864 446260 558920
rect 445753 558862 446260 558864
rect 443196 558860 443202 558862
rect 443085 558859 443151 558860
rect 445753 558859 445819 558862
rect 446254 558860 446260 558862
rect 446324 558860 446330 558924
rect 447593 558922 447659 558925
rect 453665 558924 453731 558925
rect 447726 558922 447732 558924
rect 447593 558920 447732 558922
rect 447593 558864 447598 558920
rect 447654 558864 447732 558920
rect 447593 558862 447732 558864
rect 447593 558859 447659 558862
rect 447726 558860 447732 558862
rect 447796 558860 447802 558924
rect 453614 558922 453620 558924
rect 453574 558862 453620 558922
rect 453684 558920 453731 558924
rect 453726 558864 453731 558920
rect 453614 558860 453620 558862
rect 453684 558860 453731 558864
rect 453665 558859 453731 558860
rect 454677 558924 454743 558925
rect 455965 558924 456031 558925
rect 457345 558924 457411 558925
rect 458265 558924 458331 558925
rect 460841 558924 460907 558925
rect 454677 558920 454724 558924
rect 454788 558922 454794 558924
rect 454677 558864 454682 558920
rect 454677 558860 454724 558864
rect 454788 558862 454834 558922
rect 455965 558920 456012 558924
rect 456076 558922 456082 558924
rect 457294 558922 457300 558924
rect 455965 558864 455970 558920
rect 454788 558860 454794 558862
rect 455965 558860 456012 558864
rect 456076 558862 456122 558922
rect 457254 558862 457300 558922
rect 457364 558920 457411 558924
rect 458214 558922 458220 558924
rect 457406 558864 457411 558920
rect 456076 558860 456082 558862
rect 457294 558860 457300 558862
rect 457364 558860 457411 558864
rect 458174 558862 458220 558922
rect 458284 558920 458331 558924
rect 460790 558922 460796 558924
rect 458326 558864 458331 558920
rect 458214 558860 458220 558862
rect 458284 558860 458331 558864
rect 460750 558862 460796 558922
rect 460860 558920 460907 558924
rect 460902 558864 460907 558920
rect 460790 558860 460796 558862
rect 460860 558860 460907 558864
rect 454677 558859 454743 558860
rect 455965 558859 456031 558860
rect 457345 558859 457411 558860
rect 458265 558859 458331 558860
rect 460841 558859 460907 558860
rect 461669 558924 461735 558925
rect 462589 558924 462655 558925
rect 464245 558924 464311 558925
rect 465257 558924 465323 558925
rect 461669 558920 461716 558924
rect 461780 558922 461786 558924
rect 461669 558864 461674 558920
rect 461669 558860 461716 558864
rect 461780 558862 461826 558922
rect 462589 558920 462636 558924
rect 462700 558922 462706 558924
rect 462589 558864 462594 558920
rect 461780 558860 461786 558862
rect 462589 558860 462636 558864
rect 462700 558862 462746 558922
rect 464245 558920 464292 558924
rect 464356 558922 464362 558924
rect 465206 558922 465212 558924
rect 464245 558864 464250 558920
rect 462700 558860 462706 558862
rect 464245 558860 464292 558864
rect 464356 558862 464402 558922
rect 465166 558862 465212 558922
rect 465276 558920 465323 558924
rect 465318 558864 465323 558920
rect 464356 558860 464362 558862
rect 465206 558860 465212 558862
rect 465276 558860 465323 558864
rect 461669 558859 461735 558860
rect 462589 558859 462655 558860
rect 464245 558859 464311 558860
rect 465257 558859 465323 558860
rect 466453 558922 466519 558925
rect 466862 558922 466868 558924
rect 466453 558920 466868 558922
rect 466453 558864 466458 558920
rect 466514 558864 466868 558920
rect 466453 558862 466868 558864
rect 466453 558859 466519 558862
rect 466862 558860 466868 558862
rect 466932 558860 466938 558924
rect 467833 558922 467899 558925
rect 468661 558924 468727 558925
rect 467966 558922 467972 558924
rect 467833 558920 467972 558922
rect 467833 558864 467838 558920
rect 467894 558864 467972 558920
rect 467833 558862 467972 558864
rect 467833 558859 467899 558862
rect 467966 558860 467972 558862
rect 468036 558860 468042 558924
rect 468661 558920 468708 558924
rect 468772 558922 468778 558924
rect 469213 558922 469279 558925
rect 470358 558922 470364 558924
rect 468661 558864 468666 558920
rect 468661 558860 468708 558864
rect 468772 558862 468818 558922
rect 469213 558920 470364 558922
rect 469213 558864 469218 558920
rect 469274 558864 470364 558920
rect 469213 558862 470364 558864
rect 468772 558860 468778 558862
rect 468661 558859 468727 558860
rect 469213 558859 469279 558862
rect 470358 558860 470364 558862
rect 470428 558860 470434 558924
rect 470593 558922 470659 558925
rect 471462 558922 471468 558924
rect 470593 558920 471468 558922
rect 470593 558864 470598 558920
rect 470654 558864 471468 558920
rect 470593 558862 471468 558864
rect 470593 558859 470659 558862
rect 471462 558860 471468 558862
rect 471532 558860 471538 558924
rect 471973 558922 472039 558925
rect 472750 558922 472756 558924
rect 471973 558920 472756 558922
rect 471973 558864 471978 558920
rect 472034 558864 472756 558920
rect 471973 558862 472756 558864
rect 471973 558859 472039 558862
rect 472750 558860 472756 558862
rect 472820 558860 472826 558924
rect 473353 558922 473419 558925
rect 474825 558924 474891 558925
rect 474038 558922 474044 558924
rect 473353 558920 474044 558922
rect 473353 558864 473358 558920
rect 473414 558864 474044 558920
rect 473353 558862 474044 558864
rect 473353 558859 473419 558862
rect 474038 558860 474044 558862
rect 474108 558860 474114 558924
rect 474774 558922 474780 558924
rect 474734 558862 474780 558922
rect 474844 558920 474891 558924
rect 474886 558864 474891 558920
rect 474774 558860 474780 558862
rect 474844 558860 474891 558864
rect 474825 558859 474891 558860
rect 475469 558924 475535 558925
rect 477125 558924 477191 558925
rect 478229 558924 478295 558925
rect 478965 558924 479031 558925
rect 475469 558920 475516 558924
rect 475580 558922 475586 558924
rect 475469 558864 475474 558920
rect 475469 558860 475516 558864
rect 475580 558862 475626 558922
rect 477125 558920 477172 558924
rect 477236 558922 477242 558924
rect 477125 558864 477130 558920
rect 475580 558860 475586 558862
rect 477125 558860 477172 558864
rect 477236 558862 477282 558922
rect 478229 558920 478276 558924
rect 478340 558922 478346 558924
rect 478229 558864 478234 558920
rect 477236 558860 477242 558862
rect 478229 558860 478276 558864
rect 478340 558862 478386 558922
rect 478965 558920 479012 558924
rect 479076 558922 479082 558924
rect 480529 558922 480595 558925
rect 480846 558922 480852 558924
rect 478965 558864 478970 558920
rect 478340 558860 478346 558862
rect 478965 558860 479012 558864
rect 479076 558862 479122 558922
rect 480529 558920 480852 558922
rect 480529 558864 480534 558920
rect 480590 558864 480852 558920
rect 480529 558862 480852 558864
rect 479076 558860 479082 558862
rect 475469 558859 475535 558860
rect 477125 558859 477191 558860
rect 478229 558859 478295 558860
rect 478965 558859 479031 558860
rect 480529 558859 480595 558862
rect 480846 558860 480852 558862
rect 480916 558860 480922 558924
rect 483013 558922 483079 558925
rect 483606 558922 483612 558924
rect 483013 558920 483612 558922
rect 483013 558864 483018 558920
rect 483074 558864 483612 558920
rect 483013 558862 483612 558864
rect 483013 558859 483079 558862
rect 483606 558860 483612 558862
rect 483676 558860 483682 558924
rect 69790 558724 69796 558788
rect 69860 558786 69866 558788
rect 70301 558786 70367 558789
rect 75913 558788 75979 558789
rect 78489 558788 78555 558789
rect 75862 558786 75868 558788
rect 69860 558784 70367 558786
rect 69860 558728 70306 558784
rect 70362 558728 70367 558784
rect 69860 558726 70367 558728
rect 75822 558726 75868 558786
rect 75932 558784 75979 558788
rect 78438 558786 78444 558788
rect 75974 558728 75979 558784
rect 69860 558724 69866 558726
rect 70301 558723 70367 558726
rect 75862 558724 75868 558726
rect 75932 558724 75979 558728
rect 78398 558726 78444 558786
rect 78508 558784 78555 558788
rect 78550 558728 78555 558784
rect 78438 558724 78444 558726
rect 78508 558724 78555 558728
rect 79358 558724 79364 558788
rect 79428 558786 79434 558788
rect 79501 558786 79567 558789
rect 82905 558788 82971 558789
rect 82854 558786 82860 558788
rect 79428 558784 79567 558786
rect 79428 558728 79506 558784
rect 79562 558728 79567 558784
rect 79428 558726 79567 558728
rect 82814 558726 82860 558786
rect 82924 558784 82971 558788
rect 82966 558728 82971 558784
rect 79428 558724 79434 558726
rect 75913 558723 75979 558724
rect 78489 558723 78555 558724
rect 79501 558723 79567 558726
rect 82854 558724 82860 558726
rect 82924 558724 82971 558728
rect 82905 558723 82971 558724
rect 85389 558788 85455 558789
rect 85389 558784 85436 558788
rect 85500 558786 85506 558788
rect 85389 558728 85394 558784
rect 85389 558724 85436 558728
rect 85500 558726 85546 558786
rect 85500 558724 85506 558726
rect 86166 558724 86172 558788
rect 86236 558786 86242 558788
rect 86861 558786 86927 558789
rect 86236 558784 86927 558786
rect 86236 558728 86866 558784
rect 86922 558728 86927 558784
rect 86236 558726 86927 558728
rect 86236 558724 86242 558726
rect 85389 558723 85455 558724
rect 86861 558723 86927 558726
rect 91093 558788 91159 558789
rect 93761 558788 93827 558789
rect 91093 558784 91140 558788
rect 91204 558786 91210 558788
rect 93710 558786 93716 558788
rect 91093 558728 91098 558784
rect 91093 558724 91140 558728
rect 91204 558726 91250 558786
rect 93670 558726 93716 558786
rect 93780 558784 93827 558788
rect 93822 558728 93827 558784
rect 91204 558724 91210 558726
rect 93710 558724 93716 558726
rect 93780 558724 93827 558728
rect 91093 558723 91159 558724
rect 93761 558723 93827 558724
rect 104893 558786 104959 558789
rect 105302 558786 105308 558788
rect 104893 558784 105308 558786
rect 104893 558728 104898 558784
rect 104954 558728 105308 558784
rect 104893 558726 105308 558728
rect 104893 558723 104959 558726
rect 105302 558724 105308 558726
rect 105372 558724 105378 558788
rect 202137 558786 202203 558789
rect 202454 558786 202460 558788
rect 202137 558784 202460 558786
rect 202137 558728 202142 558784
rect 202198 558728 202460 558784
rect 202137 558726 202460 558728
rect 202137 558723 202203 558726
rect 202454 558724 202460 558726
rect 202524 558724 202530 558788
rect 216622 558724 216628 558788
rect 216692 558786 216698 558788
rect 217961 558786 218027 558789
rect 216692 558784 218027 558786
rect 216692 558728 217966 558784
rect 218022 558728 218027 558784
rect 216692 558726 218027 558728
rect 216692 558724 216698 558726
rect 217961 558723 218027 558726
rect 231945 558786 232011 558789
rect 232814 558786 232820 558788
rect 231945 558784 232820 558786
rect 231945 558728 231950 558784
rect 232006 558728 232820 558784
rect 231945 558726 232820 558728
rect 231945 558723 232011 558726
rect 232814 558724 232820 558726
rect 232884 558724 232890 558788
rect 233233 558786 233299 558789
rect 234613 558788 234679 558789
rect 233550 558786 233556 558788
rect 233233 558784 233556 558786
rect 233233 558728 233238 558784
rect 233294 558728 233556 558784
rect 233233 558726 233556 558728
rect 233233 558723 233299 558726
rect 233550 558724 233556 558726
rect 233620 558724 233626 558788
rect 234613 558786 234660 558788
rect 234568 558784 234660 558786
rect 234568 558728 234618 558784
rect 234568 558726 234660 558728
rect 234613 558724 234660 558726
rect 234724 558724 234730 558788
rect 235993 558786 236059 558789
rect 320173 558788 320239 558789
rect 236126 558786 236132 558788
rect 235993 558784 236132 558786
rect 235993 558728 235998 558784
rect 236054 558728 236132 558784
rect 235993 558726 236132 558728
rect 234613 558723 234679 558724
rect 235993 558723 236059 558726
rect 236126 558724 236132 558726
rect 236196 558724 236202 558788
rect 320173 558786 320220 558788
rect 320128 558784 320220 558786
rect 320128 558728 320178 558784
rect 320128 558726 320220 558728
rect 320173 558724 320220 558726
rect 320284 558724 320290 558788
rect 354673 558786 354739 558789
rect 356053 558788 356119 558789
rect 354806 558786 354812 558788
rect 354673 558784 354812 558786
rect 354673 558728 354678 558784
rect 354734 558728 354812 558784
rect 354673 558726 354812 558728
rect 320173 558723 320239 558724
rect 354673 558723 354739 558726
rect 354806 558724 354812 558726
rect 354876 558724 354882 558788
rect 356053 558786 356100 558788
rect 356008 558784 356100 558786
rect 356008 558728 356058 558784
rect 356008 558726 356100 558728
rect 356053 558724 356100 558726
rect 356164 558724 356170 558788
rect 452653 558786 452719 558789
rect 466545 558788 466611 558789
rect 453798 558786 453804 558788
rect 452653 558784 453804 558786
rect 452653 558728 452658 558784
rect 452714 558728 453804 558784
rect 452653 558726 453804 558728
rect 356053 558723 356119 558724
rect 452653 558723 452719 558726
rect 453798 558724 453804 558726
rect 453868 558724 453874 558788
rect 466494 558786 466500 558788
rect 466454 558726 466500 558786
rect 466564 558784 466611 558788
rect 466606 558728 466611 558784
rect 466494 558724 466500 558726
rect 466564 558724 466611 558728
rect 466545 558723 466611 558724
rect 467925 558786 467991 558789
rect 470041 558788 470107 558789
rect 471329 558788 471395 558789
rect 469070 558786 469076 558788
rect 467925 558784 469076 558786
rect 467925 558728 467930 558784
rect 467986 558728 469076 558784
rect 467925 558726 469076 558728
rect 467925 558723 467991 558726
rect 469070 558724 469076 558726
rect 469140 558724 469146 558788
rect 469990 558786 469996 558788
rect 469950 558726 469996 558786
rect 470060 558784 470107 558788
rect 471278 558786 471284 558788
rect 470102 558728 470107 558784
rect 469990 558724 469996 558726
rect 470060 558724 470107 558728
rect 471238 558726 471284 558786
rect 471348 558784 471395 558788
rect 471390 558728 471395 558784
rect 471278 558724 471284 558726
rect 471348 558724 471395 558728
rect 470041 558723 470107 558724
rect 471329 558723 471395 558724
rect 472157 558788 472223 558789
rect 472157 558784 472204 558788
rect 472268 558786 472274 558788
rect 480345 558786 480411 558789
rect 481633 558788 481699 558789
rect 480478 558786 480484 558788
rect 472157 558728 472162 558784
rect 472157 558724 472204 558728
rect 472268 558726 472314 558786
rect 480345 558784 480484 558786
rect 480345 558728 480350 558784
rect 480406 558728 480484 558784
rect 480345 558726 480484 558728
rect 472268 558724 472274 558726
rect 472157 558723 472223 558724
rect 480345 558723 480411 558726
rect 480478 558724 480484 558726
rect 480548 558724 480554 558788
rect 481582 558724 481588 558788
rect 481652 558786 481699 558788
rect 481652 558784 481744 558786
rect 481694 558728 481744 558784
rect 481652 558726 481744 558728
rect 481652 558724 481699 558726
rect 481633 558723 481699 558724
rect 86350 558588 86356 558652
rect 86420 558650 86426 558652
rect 86677 558650 86743 558653
rect 93577 558652 93643 558653
rect 204897 558652 204963 558653
rect 93526 558650 93532 558652
rect 86420 558648 86743 558650
rect 86420 558592 86682 558648
rect 86738 558592 86743 558648
rect 86420 558590 86743 558592
rect 93486 558590 93532 558650
rect 93596 558648 93643 558652
rect 204846 558650 204852 558652
rect 93638 558592 93643 558648
rect 86420 558588 86426 558590
rect 86677 558587 86743 558590
rect 93526 558588 93532 558590
rect 93596 558588 93643 558592
rect 204806 558590 204852 558650
rect 204916 558648 204963 558652
rect 204958 558592 204963 558648
rect 204846 558588 204852 558590
rect 204916 558588 204963 558592
rect 93577 558587 93643 558588
rect 204897 558587 204963 558588
rect 210509 558652 210575 558653
rect 210509 558648 210556 558652
rect 210620 558650 210626 558652
rect 211153 558650 211219 558653
rect 217542 558650 217548 558652
rect 210509 558592 210514 558648
rect 210509 558588 210556 558592
rect 210620 558590 210666 558650
rect 211153 558648 217548 558650
rect 211153 558592 211158 558648
rect 211214 558592 217548 558648
rect 211153 558590 217548 558592
rect 210620 558588 210626 558590
rect 210509 558587 210575 558588
rect 211153 558587 211219 558590
rect 217542 558588 217548 558590
rect 217612 558650 217618 558652
rect 220721 558650 220787 558653
rect 231853 558652 231919 558653
rect 237373 558652 237439 558653
rect 231853 558650 231900 558652
rect 217612 558648 220787 558650
rect 217612 558592 220726 558648
rect 220782 558592 220787 558648
rect 217612 558590 220787 558592
rect 231808 558648 231900 558650
rect 231808 558592 231858 558648
rect 231808 558590 231900 558592
rect 217612 558588 217618 558590
rect 220721 558587 220787 558590
rect 231853 558588 231900 558590
rect 231964 558588 231970 558652
rect 237373 558650 237420 558652
rect 237328 558648 237420 558650
rect 237328 558592 237378 558648
rect 237328 558590 237420 558592
rect 237373 558588 237420 558590
rect 237484 558588 237490 558652
rect 292573 558650 292639 558653
rect 302141 558650 302207 558653
rect 292573 558648 302207 558650
rect 292573 558592 292578 558648
rect 292634 558592 302146 558648
rect 302202 558592 302207 558648
rect 292573 558590 302207 558592
rect 231853 558587 231919 558588
rect 237373 558587 237439 558588
rect 292573 558587 292639 558590
rect 302141 558587 302207 558590
rect 318793 558650 318859 558653
rect 318926 558650 318932 558652
rect 318793 558648 318932 558650
rect 318793 558592 318798 558648
rect 318854 558592 318932 558648
rect 318793 558590 318932 558592
rect 318793 558587 318859 558590
rect 318926 558588 318932 558590
rect 318996 558588 319002 558652
rect 452694 558588 452700 558652
rect 452764 558650 452770 558652
rect 453297 558650 453363 558653
rect 453941 558650 454007 558653
rect 452764 558648 454007 558650
rect 452764 558592 453302 558648
rect 453358 558592 453946 558648
rect 454002 558592 454007 558648
rect 452764 558590 454007 558592
rect 452764 558588 452770 558590
rect 453297 558587 453363 558590
rect 453941 558587 454007 558590
rect 459502 558588 459508 558652
rect 459572 558650 459578 558652
rect 459645 558650 459711 558653
rect 462957 558650 463023 558653
rect 459572 558648 463023 558650
rect 459572 558592 459650 558648
rect 459706 558592 462962 558648
rect 463018 558592 463023 558648
rect 459572 558590 463023 558592
rect 459572 558588 459578 558590
rect 459645 558587 459711 558590
rect 462957 558587 463023 558590
rect 467782 558588 467788 558652
rect 467852 558650 467858 558652
rect 468017 558650 468083 558653
rect 467852 558648 468083 558650
rect 467852 558592 468022 558648
rect 468078 558592 468083 558648
rect 467852 558590 468083 558592
rect 467852 558588 467858 558590
rect 468017 558587 468083 558590
rect 473445 558652 473511 558653
rect 473445 558648 473492 558652
rect 473556 558650 473562 558652
rect 484393 558650 484459 558653
rect 488533 558652 488599 558653
rect 484710 558650 484716 558652
rect 473445 558592 473450 558648
rect 473445 558588 473492 558592
rect 473556 558590 473602 558650
rect 484393 558648 484716 558650
rect 484393 558592 484398 558648
rect 484454 558592 484716 558648
rect 484393 558590 484716 558592
rect 473556 558588 473562 558590
rect 473445 558587 473511 558588
rect 484393 558587 484459 558590
rect 484710 558588 484716 558590
rect 484780 558588 484786 558652
rect 488533 558650 488580 558652
rect 488488 558648 488580 558650
rect 488488 558592 488538 558648
rect 488488 558590 488580 558592
rect 488533 558588 488580 558590
rect 488644 558588 488650 558652
rect 488533 558587 488599 558588
rect 99373 558516 99439 558517
rect 99373 558512 99420 558516
rect 99484 558514 99490 558516
rect 108297 558514 108363 558517
rect 108614 558514 108620 558516
rect 99373 558456 99378 558512
rect 99373 558452 99420 558456
rect 99484 558454 99530 558514
rect 108297 558512 108620 558514
rect 108297 558456 108302 558512
rect 108358 558456 108620 558512
rect 108297 558454 108620 558456
rect 99484 558452 99490 558454
rect 99373 558451 99439 558452
rect 108297 558451 108363 558454
rect 108614 558452 108620 558454
rect 108684 558452 108690 558516
rect 230473 558514 230539 558517
rect 230606 558514 230612 558516
rect 230473 558512 230612 558514
rect 230473 558456 230478 558512
rect 230534 558456 230612 558512
rect 230473 558454 230612 558456
rect 230473 558451 230539 558454
rect 230606 558452 230612 558454
rect 230676 558452 230682 558516
rect 357433 558514 357499 558517
rect 449893 558516 449959 558517
rect 357566 558514 357572 558516
rect 357433 558512 357572 558514
rect 357433 558456 357438 558512
rect 357494 558456 357572 558512
rect 357433 558454 357572 558456
rect 357433 558451 357499 558454
rect 357566 558452 357572 558454
rect 357636 558452 357642 558516
rect 449893 558514 449940 558516
rect 449848 558512 449940 558514
rect 449848 558456 449898 558512
rect 449848 558454 449940 558456
rect 449893 558452 449940 558454
rect 450004 558452 450010 558516
rect 476113 558514 476179 558517
rect 477350 558514 477356 558516
rect 476113 558512 477356 558514
rect 476113 558456 476118 558512
rect 476174 558456 477356 558512
rect 476113 558454 477356 558456
rect 449893 558451 449959 558452
rect 476113 558451 476179 558454
rect 477350 558452 477356 558454
rect 477420 558452 477426 558516
rect 481633 558514 481699 558517
rect 482134 558514 482140 558516
rect 481633 558512 482140 558514
rect 481633 558456 481638 558512
rect 481694 558456 482140 558512
rect 481633 558454 482140 558456
rect 481633 558451 481699 558454
rect 482134 558452 482140 558454
rect 482204 558452 482210 558516
rect 485773 558514 485839 558517
rect 485998 558514 486004 558516
rect 485773 558512 486004 558514
rect 485773 558456 485778 558512
rect 485834 558456 486004 558512
rect 485773 558454 486004 558456
rect 485773 558451 485839 558454
rect 485998 558452 486004 558454
rect 486068 558452 486074 558516
rect 487153 558514 487219 558517
rect 487286 558514 487292 558516
rect 487153 558512 487292 558514
rect 487153 558456 487158 558512
rect 487214 558456 487292 558512
rect 487153 558454 487292 558456
rect 487153 558451 487219 558454
rect 487286 558452 487292 558454
rect 487356 558452 487362 558516
rect 62021 558378 62087 558381
rect 238753 558380 238819 558381
rect 197302 558378 197308 558380
rect 62021 558376 197308 558378
rect 62021 558320 62026 558376
rect 62082 558320 197308 558376
rect 62021 558318 197308 558320
rect 62021 558315 62087 558318
rect 197302 558316 197308 558318
rect 197372 558316 197378 558380
rect 238702 558316 238708 558380
rect 238772 558378 238819 558380
rect 356697 558378 356763 558381
rect 476205 558380 476271 558381
rect 474958 558378 474964 558380
rect 238772 558376 238864 558378
rect 238814 558320 238864 558376
rect 238772 558318 238864 558320
rect 356697 558376 474964 558378
rect 356697 558320 356702 558376
rect 356758 558320 474964 558376
rect 356697 558318 474964 558320
rect 238772 558316 238819 558318
rect 238753 558315 238819 558316
rect 356697 558315 356763 558318
rect 474958 558316 474964 558318
rect 475028 558316 475034 558380
rect 476205 558378 476252 558380
rect 476160 558376 476252 558378
rect 476160 558320 476210 558376
rect 476160 558318 476252 558320
rect 476205 558316 476252 558318
rect 476316 558316 476322 558380
rect 477493 558378 477559 558381
rect 478454 558378 478460 558380
rect 477493 558376 478460 558378
rect 477493 558320 477498 558376
rect 477554 558320 478460 558376
rect 477493 558318 478460 558320
rect 476205 558315 476271 558316
rect 477493 558315 477559 558318
rect 478454 558316 478460 558318
rect 478524 558316 478530 558380
rect 63401 558242 63467 558245
rect 198774 558242 198780 558244
rect 63401 558240 198780 558242
rect 63401 558184 63406 558240
rect 63462 558184 198780 558240
rect 63401 558182 198780 558184
rect 63401 558179 63467 558182
rect 198774 558180 198780 558182
rect 198844 558180 198850 558244
rect 283649 558242 283715 558245
rect 448462 558242 448468 558244
rect 283649 558240 448468 558242
rect 283649 558184 283654 558240
rect 283710 558184 448468 558240
rect 283649 558182 448468 558184
rect 283649 558179 283715 558182
rect 448462 558180 448468 558182
rect 448532 558180 448538 558244
rect 478873 558242 478939 558245
rect 479742 558242 479748 558244
rect 478873 558240 479748 558242
rect 478873 558184 478878 558240
rect 478934 558184 479748 558240
rect 478873 558182 479748 558184
rect 478873 558179 478939 558182
rect 479742 558180 479748 558182
rect 479812 558180 479818 558244
rect 483013 558242 483079 558245
rect 483422 558242 483428 558244
rect 483013 558240 483428 558242
rect 483013 558184 483018 558240
rect 483074 558184 483428 558240
rect 483013 558182 483428 558184
rect 483013 558179 483079 558182
rect 483422 558180 483428 558182
rect 483492 558180 483498 558244
rect 484393 558242 484459 558245
rect 485630 558242 485636 558244
rect 484393 558240 485636 558242
rect 484393 558184 484398 558240
rect 484454 558184 485636 558240
rect 484393 558182 485636 558184
rect 484393 558179 484459 558182
rect 485630 558180 485636 558182
rect 485700 558180 485706 558244
rect 485773 558242 485839 558245
rect 486918 558242 486924 558244
rect 485773 558240 486924 558242
rect 485773 558184 485778 558240
rect 485834 558184 486924 558240
rect 485773 558182 486924 558184
rect 485773 558179 485839 558182
rect 486918 558180 486924 558182
rect 486988 558180 486994 558244
rect 64270 558044 64276 558108
rect 64340 558106 64346 558108
rect 194409 558106 194475 558109
rect 64340 558104 194475 558106
rect 64340 558048 194414 558104
rect 194470 558048 194475 558104
rect 64340 558046 194475 558048
rect 64340 558044 64346 558046
rect 194409 558043 194475 558046
rect 238334 558044 238340 558108
rect 238404 558106 238410 558108
rect 238661 558106 238727 558109
rect 238404 558104 238727 558106
rect 238404 558048 238666 558104
rect 238722 558048 238727 558104
rect 238404 558046 238727 558048
rect 238404 558044 238410 558046
rect 238661 558043 238727 558046
rect 451273 558106 451339 558109
rect 451406 558106 451412 558108
rect 451273 558104 451412 558106
rect 451273 558048 451278 558104
rect 451334 558048 451412 558104
rect 451273 558046 451412 558048
rect 451273 558043 451339 558046
rect 451406 558044 451412 558046
rect 451476 558044 451482 558108
rect 483105 558106 483171 558109
rect 484158 558106 484164 558108
rect 483105 558104 484164 558106
rect 483105 558048 483110 558104
rect 483166 558048 484164 558104
rect 483105 558046 484164 558048
rect 483105 558043 483171 558046
rect 484158 558044 484164 558046
rect 484228 558044 484234 558108
rect 488533 558106 488599 558109
rect 489126 558106 489132 558108
rect 488533 558104 489132 558106
rect 488533 558048 488538 558104
rect 488594 558048 489132 558104
rect 488533 558046 489132 558048
rect 488533 558043 488599 558046
rect 489126 558044 489132 558046
rect 489196 558044 489202 558108
rect 487153 557970 487219 557973
rect 487838 557970 487844 557972
rect 487153 557968 487844 557970
rect 487153 557912 487158 557968
rect 487214 557912 487844 557968
rect 487153 557910 487844 557912
rect 487153 557907 487219 557910
rect 487838 557908 487844 557910
rect 487908 557908 487914 557972
rect 100017 557834 100083 557837
rect 100334 557834 100340 557836
rect 100017 557832 100340 557834
rect 100017 557776 100022 557832
rect 100078 557776 100340 557832
rect 100017 557774 100340 557776
rect 100017 557771 100083 557774
rect 100334 557772 100340 557774
rect 100404 557772 100410 557836
rect 100845 557698 100911 557701
rect 101397 557698 101463 557701
rect 106273 557700 106339 557701
rect 101622 557698 101628 557700
rect 100845 557696 101628 557698
rect 100845 557640 100850 557696
rect 100906 557640 101402 557696
rect 101458 557640 101628 557696
rect 100845 557638 101628 557640
rect 100845 557635 100911 557638
rect 101397 557635 101463 557638
rect 101622 557636 101628 557638
rect 101692 557636 101698 557700
rect 106222 557698 106228 557700
rect 106146 557638 106228 557698
rect 106292 557698 106339 557700
rect 106917 557698 106983 557701
rect 106292 557696 106983 557698
rect 106334 557640 106922 557696
rect 106978 557640 106983 557696
rect 106222 557636 106228 557638
rect 106292 557638 106983 557640
rect 106292 557636 106339 557638
rect 106273 557635 106339 557636
rect 106917 557635 106983 557638
rect 207054 557636 207060 557700
rect 207124 557698 207130 557700
rect 207657 557698 207723 557701
rect 207124 557696 207723 557698
rect 207124 557640 207662 557696
rect 207718 557640 207723 557696
rect 207124 557638 207723 557640
rect 207124 557636 207130 557638
rect 207657 557635 207723 557638
rect 209037 557698 209103 557701
rect 209630 557698 209636 557700
rect 209037 557696 209636 557698
rect 209037 557640 209042 557696
rect 209098 557640 209636 557696
rect 209037 557638 209636 557640
rect 209037 557635 209103 557638
rect 209630 557636 209636 557638
rect 209700 557636 209706 557700
rect 210366 557636 210372 557700
rect 210436 557698 210442 557700
rect 210969 557698 211035 557701
rect 210436 557696 211035 557698
rect 210436 557640 210974 557696
rect 211030 557640 211035 557696
rect 210436 557638 211035 557640
rect 210436 557636 210442 557638
rect 210969 557635 211035 557638
rect 217358 557636 217364 557700
rect 217428 557698 217434 557700
rect 217869 557698 217935 557701
rect 217428 557696 217935 557698
rect 217428 557640 217874 557696
rect 217930 557640 217935 557696
rect 217428 557638 217935 557640
rect 217428 557636 217434 557638
rect 217869 557635 217935 557638
rect 225638 557636 225644 557700
rect 225708 557698 225714 557700
rect 226241 557698 226307 557701
rect 225708 557696 226307 557698
rect 225708 557640 226246 557696
rect 226302 557640 226307 557696
rect 225708 557638 226307 557640
rect 225708 557636 225714 557638
rect 226241 557635 226307 557638
rect 232630 557636 232636 557700
rect 232700 557698 232706 557700
rect 233141 557698 233207 557701
rect 232700 557696 233207 557698
rect 232700 557640 233146 557696
rect 233202 557640 233207 557696
rect 232700 557638 233207 557640
rect 232700 557636 232706 557638
rect 233141 557635 233207 557638
rect 324814 557636 324820 557700
rect 324884 557698 324890 557700
rect 324957 557698 325023 557701
rect 324884 557696 325023 557698
rect 324884 557640 324962 557696
rect 325018 557640 325023 557696
rect 324884 557638 325023 557640
rect 324884 557636 324890 557638
rect 324957 557635 325023 557638
rect 326102 557636 326108 557700
rect 326172 557698 326178 557700
rect 326337 557698 326403 557701
rect 326172 557696 326403 557698
rect 326172 557640 326342 557696
rect 326398 557640 326403 557696
rect 326172 557638 326403 557640
rect 326172 557636 326178 557638
rect 326337 557635 326403 557638
rect 327022 557636 327028 557700
rect 327092 557698 327098 557700
rect 327717 557698 327783 557701
rect 327092 557696 327783 557698
rect 327092 557640 327722 557696
rect 327778 557640 327783 557696
rect 327092 557638 327783 557640
rect 327092 557636 327098 557638
rect 327717 557635 327783 557638
rect 329925 557698 329991 557701
rect 331070 557698 331076 557700
rect 329925 557696 331076 557698
rect 329925 557640 329930 557696
rect 329986 557640 331076 557696
rect 329925 557638 331076 557640
rect 329925 557635 329991 557638
rect 331070 557636 331076 557638
rect 331140 557636 331146 557700
rect 336825 557698 336891 557701
rect 337878 557698 337884 557700
rect 336825 557696 337884 557698
rect 336825 557640 336830 557696
rect 336886 557640 337884 557696
rect 336825 557638 337884 557640
rect 336825 557635 336891 557638
rect 337878 557636 337884 557638
rect 337948 557636 337954 557700
rect 343725 557698 343791 557701
rect 344870 557698 344876 557700
rect 343725 557696 344876 557698
rect 343725 557640 343730 557696
rect 343786 557640 344876 557696
rect 343725 557638 344876 557640
rect 343725 557635 343791 557638
rect 344870 557636 344876 557638
rect 344940 557636 344946 557700
rect 352005 557698 352071 557701
rect 353150 557698 353156 557700
rect 352005 557696 353156 557698
rect 352005 557640 352010 557696
rect 352066 557640 353156 557696
rect 352005 557638 353156 557640
rect 352005 557635 352071 557638
rect 353150 557636 353156 557638
rect 353220 557636 353226 557700
rect 461025 557698 461091 557701
rect 483013 557700 483079 557701
rect 462078 557698 462084 557700
rect 461025 557696 462084 557698
rect 461025 557640 461030 557696
rect 461086 557640 462084 557696
rect 461025 557638 462084 557640
rect 461025 557635 461091 557638
rect 462078 557636 462084 557638
rect 462148 557636 462154 557700
rect 483013 557698 483060 557700
rect 482968 557696 483060 557698
rect 482968 557640 483018 557696
rect 482968 557638 483060 557640
rect 483013 557636 483060 557638
rect 483124 557636 483130 557700
rect 483013 557635 483079 557636
rect 101438 557500 101444 557564
rect 101508 557562 101514 557564
rect 102041 557562 102107 557565
rect 102777 557564 102843 557565
rect 102726 557562 102732 557564
rect 101508 557560 102107 557562
rect 101508 557504 102046 557560
rect 102102 557504 102107 557560
rect 101508 557502 102107 557504
rect 102686 557502 102732 557562
rect 102796 557560 102843 557564
rect 102838 557504 102843 557560
rect 101508 557500 101514 557502
rect 102041 557499 102107 557502
rect 102726 557500 102732 557502
rect 102796 557500 102843 557504
rect 103278 557500 103284 557564
rect 103348 557562 103354 557564
rect 103421 557562 103487 557565
rect 103348 557560 103487 557562
rect 103348 557504 103426 557560
rect 103482 557504 103487 557560
rect 103348 557502 103487 557504
rect 103348 557500 103354 557502
rect 102777 557499 102843 557500
rect 103421 557499 103487 557502
rect 104014 557500 104020 557564
rect 104084 557562 104090 557564
rect 104157 557562 104223 557565
rect 104084 557560 104223 557562
rect 104084 557504 104162 557560
rect 104218 557504 104223 557560
rect 104084 557502 104223 557504
rect 104084 557500 104090 557502
rect 104157 557499 104223 557502
rect 105302 557500 105308 557564
rect 105372 557562 105378 557564
rect 105537 557562 105603 557565
rect 105372 557560 105603 557562
rect 105372 557504 105542 557560
rect 105598 557504 105603 557560
rect 105372 557502 105603 557504
rect 105372 557500 105378 557502
rect 105537 557499 105603 557502
rect 106038 557500 106044 557564
rect 106108 557562 106114 557564
rect 106181 557562 106247 557565
rect 107653 557564 107719 557565
rect 107653 557562 107700 557564
rect 106108 557560 106247 557562
rect 106108 557504 106186 557560
rect 106242 557504 106247 557560
rect 106108 557502 106247 557504
rect 107572 557560 107700 557562
rect 107764 557562 107770 557564
rect 108481 557562 108547 557565
rect 107764 557560 108547 557562
rect 107572 557504 107658 557560
rect 107764 557504 108486 557560
rect 108542 557504 108547 557560
rect 107572 557502 107700 557504
rect 106108 557500 106114 557502
rect 106181 557499 106247 557502
rect 107653 557500 107700 557502
rect 107764 557502 108547 557504
rect 107764 557500 107770 557502
rect 107653 557499 107719 557500
rect 108481 557499 108547 557502
rect 108982 557500 108988 557564
rect 109052 557562 109058 557564
rect 110321 557562 110387 557565
rect 206921 557564 206987 557565
rect 109052 557560 110387 557562
rect 109052 557504 110326 557560
rect 110382 557504 110387 557560
rect 109052 557502 110387 557504
rect 109052 557500 109058 557502
rect 110321 557499 110387 557502
rect 206870 557500 206876 557564
rect 206940 557562 206987 557564
rect 206940 557560 207032 557562
rect 206982 557504 207032 557560
rect 206940 557502 207032 557504
rect 206940 557500 206987 557502
rect 207974 557500 207980 557564
rect 208044 557562 208050 557564
rect 208301 557562 208367 557565
rect 208044 557560 208367 557562
rect 208044 557504 208306 557560
rect 208362 557504 208367 557560
rect 208044 557502 208367 557504
rect 208044 557500 208050 557502
rect 206921 557499 206987 557500
rect 208301 557499 208367 557502
rect 209262 557500 209268 557564
rect 209332 557562 209338 557564
rect 209681 557562 209747 557565
rect 209332 557560 209747 557562
rect 209332 557504 209686 557560
rect 209742 557504 209747 557560
rect 209332 557502 209747 557504
rect 209332 557500 209338 557502
rect 209681 557499 209747 557502
rect 210918 557500 210924 557564
rect 210988 557562 210994 557564
rect 211061 557562 211127 557565
rect 212441 557564 212507 557565
rect 210988 557560 211127 557562
rect 210988 557504 211066 557560
rect 211122 557504 211127 557560
rect 210988 557502 211127 557504
rect 210988 557500 210994 557502
rect 211061 557499 211127 557502
rect 212390 557500 212396 557564
rect 212460 557562 212507 557564
rect 212460 557560 212552 557562
rect 212502 557504 212552 557560
rect 212460 557502 212552 557504
rect 212460 557500 212507 557502
rect 213494 557500 213500 557564
rect 213564 557562 213570 557564
rect 213821 557562 213887 557565
rect 213564 557560 213887 557562
rect 213564 557504 213826 557560
rect 213882 557504 213887 557560
rect 213564 557502 213887 557504
rect 213564 557500 213570 557502
rect 212441 557499 212507 557500
rect 213821 557499 213887 557502
rect 214782 557500 214788 557564
rect 214852 557562 214858 557564
rect 215201 557562 215267 557565
rect 214852 557560 215267 557562
rect 214852 557504 215206 557560
rect 215262 557504 215267 557560
rect 214852 557502 215267 557504
rect 214852 557500 214858 557502
rect 215201 557499 215267 557502
rect 216254 557500 216260 557564
rect 216324 557562 216330 557564
rect 216581 557562 216647 557565
rect 217961 557564 218027 557565
rect 216324 557560 216647 557562
rect 216324 557504 216586 557560
rect 216642 557504 216647 557560
rect 216324 557502 216647 557504
rect 216324 557500 216330 557502
rect 216581 557499 216647 557502
rect 217910 557500 217916 557564
rect 217980 557562 218027 557564
rect 217980 557560 218072 557562
rect 218022 557504 218072 557560
rect 217980 557502 218072 557504
rect 217980 557500 218027 557502
rect 219198 557500 219204 557564
rect 219268 557562 219274 557564
rect 219341 557562 219407 557565
rect 220721 557564 220787 557565
rect 219268 557560 219407 557562
rect 219268 557504 219346 557560
rect 219402 557504 219407 557560
rect 219268 557502 219407 557504
rect 219268 557500 219274 557502
rect 217961 557499 218027 557500
rect 219341 557499 219407 557502
rect 220670 557500 220676 557564
rect 220740 557562 220787 557564
rect 220740 557560 220832 557562
rect 220782 557504 220832 557560
rect 220740 557502 220832 557504
rect 220740 557500 220787 557502
rect 221958 557500 221964 557564
rect 222028 557562 222034 557564
rect 222101 557562 222167 557565
rect 222028 557560 222167 557562
rect 222028 557504 222106 557560
rect 222162 557504 222167 557560
rect 222028 557502 222167 557504
rect 222028 557500 222034 557502
rect 220721 557499 220787 557500
rect 222101 557499 222167 557502
rect 223246 557500 223252 557564
rect 223316 557562 223322 557564
rect 223481 557562 223547 557565
rect 223316 557560 223547 557562
rect 223316 557504 223486 557560
rect 223542 557504 223547 557560
rect 223316 557502 223547 557504
rect 223316 557500 223322 557502
rect 223481 557499 223547 557502
rect 224350 557500 224356 557564
rect 224420 557562 224426 557564
rect 224861 557562 224927 557565
rect 226149 557564 226215 557565
rect 226149 557562 226196 557564
rect 224420 557560 224927 557562
rect 224420 557504 224866 557560
rect 224922 557504 224927 557560
rect 224420 557502 224927 557504
rect 226104 557560 226196 557562
rect 226104 557504 226154 557560
rect 226104 557502 226196 557504
rect 224420 557500 224426 557502
rect 224861 557499 224927 557502
rect 226149 557500 226196 557502
rect 226260 557500 226266 557564
rect 227478 557500 227484 557564
rect 227548 557562 227554 557564
rect 227621 557562 227687 557565
rect 227548 557560 227687 557562
rect 227548 557504 227626 557560
rect 227682 557504 227687 557560
rect 227548 557502 227687 557504
rect 227548 557500 227554 557502
rect 226149 557499 226215 557500
rect 227621 557499 227687 557502
rect 228766 557500 228772 557564
rect 228836 557562 228842 557564
rect 229001 557562 229067 557565
rect 228836 557560 229067 557562
rect 228836 557504 229006 557560
rect 229062 557504 229067 557560
rect 228836 557502 229067 557504
rect 228836 557500 228842 557502
rect 229001 557499 229067 557502
rect 230238 557500 230244 557564
rect 230308 557562 230314 557564
rect 230381 557562 230447 557565
rect 230308 557560 230447 557562
rect 230308 557504 230386 557560
rect 230442 557504 230447 557560
rect 230308 557502 230447 557504
rect 230308 557500 230314 557502
rect 230381 557499 230447 557502
rect 230790 557500 230796 557564
rect 230860 557562 230866 557564
rect 231761 557562 231827 557565
rect 233049 557564 233115 557565
rect 234521 557564 234587 557565
rect 230860 557560 231827 557562
rect 230860 557504 231766 557560
rect 231822 557504 231827 557560
rect 230860 557502 231827 557504
rect 230860 557500 230866 557502
rect 231761 557499 231827 557502
rect 232998 557500 233004 557564
rect 233068 557562 233115 557564
rect 234470 557562 234476 557564
rect 233068 557560 233160 557562
rect 233110 557504 233160 557560
rect 233068 557502 233160 557504
rect 234430 557502 234476 557562
rect 234540 557560 234587 557564
rect 234582 557504 234587 557560
rect 233068 557500 233115 557502
rect 234470 557500 234476 557502
rect 234540 557500 234587 557504
rect 233049 557499 233115 557500
rect 234521 557499 234587 557500
rect 321553 557562 321619 557565
rect 322790 557562 322796 557564
rect 321553 557560 322796 557562
rect 321553 557504 321558 557560
rect 321614 557504 322796 557560
rect 321553 557502 322796 557504
rect 321553 557499 321619 557502
rect 322790 557500 322796 557502
rect 322860 557500 322866 557564
rect 322933 557562 322999 557565
rect 324078 557562 324084 557564
rect 322933 557560 324084 557562
rect 322933 557504 322938 557560
rect 322994 557504 324084 557560
rect 322933 557502 324084 557504
rect 322933 557499 322999 557502
rect 324078 557500 324084 557502
rect 324148 557500 324154 557564
rect 324313 557562 324379 557565
rect 325366 557562 325372 557564
rect 324313 557560 325372 557562
rect 324313 557504 324318 557560
rect 324374 557504 325372 557560
rect 324313 557502 325372 557504
rect 324313 557499 324379 557502
rect 325366 557500 325372 557502
rect 325436 557500 325442 557564
rect 325693 557562 325759 557565
rect 326286 557562 326292 557564
rect 325693 557560 326292 557562
rect 325693 557504 325698 557560
rect 325754 557504 326292 557560
rect 325693 557502 326292 557504
rect 325693 557499 325759 557502
rect 326286 557500 326292 557502
rect 326356 557500 326362 557564
rect 327073 557562 327139 557565
rect 327574 557562 327580 557564
rect 327073 557560 327580 557562
rect 327073 557504 327078 557560
rect 327134 557504 327580 557560
rect 327073 557502 327580 557504
rect 327073 557499 327139 557502
rect 327574 557500 327580 557502
rect 327644 557500 327650 557564
rect 328453 557562 328519 557565
rect 329833 557564 329899 557565
rect 328862 557562 328868 557564
rect 328453 557560 328868 557562
rect 328453 557504 328458 557560
rect 328514 557504 328868 557560
rect 328453 557502 328868 557504
rect 328453 557499 328519 557502
rect 328862 557500 328868 557502
rect 328932 557500 328938 557564
rect 329782 557500 329788 557564
rect 329852 557562 329899 557564
rect 331213 557562 331279 557565
rect 332358 557562 332364 557564
rect 329852 557560 329944 557562
rect 329894 557504 329944 557560
rect 329852 557502 329944 557504
rect 331213 557560 332364 557562
rect 331213 557504 331218 557560
rect 331274 557504 332364 557560
rect 331213 557502 332364 557504
rect 329852 557500 329899 557502
rect 329833 557499 329899 557500
rect 331213 557499 331279 557502
rect 332358 557500 332364 557502
rect 332428 557500 332434 557564
rect 332593 557562 332659 557565
rect 333278 557562 333284 557564
rect 332593 557560 333284 557562
rect 332593 557504 332598 557560
rect 332654 557504 333284 557560
rect 332593 557502 333284 557504
rect 332593 557499 332659 557502
rect 333278 557500 333284 557502
rect 333348 557500 333354 557564
rect 333973 557562 334039 557565
rect 334566 557562 334572 557564
rect 333973 557560 334572 557562
rect 333973 557504 333978 557560
rect 334034 557504 334572 557560
rect 333973 557502 334572 557504
rect 333973 557499 334039 557502
rect 334566 557500 334572 557502
rect 334636 557500 334642 557564
rect 335353 557562 335419 557565
rect 336733 557564 336799 557565
rect 335854 557562 335860 557564
rect 335353 557560 335860 557562
rect 335353 557504 335358 557560
rect 335414 557504 335860 557560
rect 335353 557502 335860 557504
rect 335353 557499 335419 557502
rect 335854 557500 335860 557502
rect 335924 557500 335930 557564
rect 336733 557562 336780 557564
rect 336688 557560 336780 557562
rect 336688 557504 336738 557560
rect 336688 557502 336780 557504
rect 336733 557500 336780 557502
rect 336844 557500 336850 557564
rect 338113 557562 338179 557565
rect 339166 557562 339172 557564
rect 338113 557560 339172 557562
rect 338113 557504 338118 557560
rect 338174 557504 339172 557560
rect 338113 557502 339172 557504
rect 336733 557499 336799 557500
rect 338113 557499 338179 557502
rect 339166 557500 339172 557502
rect 339236 557500 339242 557564
rect 339493 557562 339559 557565
rect 340454 557562 340460 557564
rect 339493 557560 340460 557562
rect 339493 557504 339498 557560
rect 339554 557504 340460 557560
rect 339493 557502 340460 557504
rect 339493 557499 339559 557502
rect 340454 557500 340460 557502
rect 340524 557500 340530 557564
rect 340873 557562 340939 557565
rect 341742 557562 341748 557564
rect 340873 557560 341748 557562
rect 340873 557504 340878 557560
rect 340934 557504 341748 557560
rect 340873 557502 341748 557504
rect 340873 557499 340939 557502
rect 341742 557500 341748 557502
rect 341812 557500 341818 557564
rect 342253 557562 342319 557565
rect 342662 557562 342668 557564
rect 342253 557560 342668 557562
rect 342253 557504 342258 557560
rect 342314 557504 342668 557560
rect 342253 557502 342668 557504
rect 342253 557499 342319 557502
rect 342662 557500 342668 557502
rect 342732 557500 342738 557564
rect 343633 557562 343699 557565
rect 343950 557562 343956 557564
rect 343633 557560 343956 557562
rect 343633 557504 343638 557560
rect 343694 557504 343956 557560
rect 343633 557502 343956 557504
rect 343633 557499 343699 557502
rect 343950 557500 343956 557502
rect 344020 557500 344026 557564
rect 345013 557562 345079 557565
rect 346158 557562 346164 557564
rect 345013 557560 346164 557562
rect 345013 557504 345018 557560
rect 345074 557504 346164 557560
rect 345013 557502 346164 557504
rect 345013 557499 345079 557502
rect 346158 557500 346164 557502
rect 346228 557500 346234 557564
rect 346393 557562 346459 557565
rect 347446 557562 347452 557564
rect 346393 557560 347452 557562
rect 346393 557504 346398 557560
rect 346454 557504 347452 557560
rect 346393 557502 347452 557504
rect 346393 557499 346459 557502
rect 347446 557500 347452 557502
rect 347516 557500 347522 557564
rect 347773 557562 347839 557565
rect 348734 557562 348740 557564
rect 347773 557560 348740 557562
rect 347773 557504 347778 557560
rect 347834 557504 348740 557560
rect 347773 557502 348740 557504
rect 347773 557499 347839 557502
rect 348734 557500 348740 557502
rect 348804 557500 348810 557564
rect 349153 557562 349219 557565
rect 349654 557562 349660 557564
rect 349153 557560 349660 557562
rect 349153 557504 349158 557560
rect 349214 557504 349660 557560
rect 349153 557502 349660 557504
rect 349153 557499 349219 557502
rect 349654 557500 349660 557502
rect 349724 557500 349730 557564
rect 350533 557562 350599 557565
rect 350942 557562 350948 557564
rect 350533 557560 350948 557562
rect 350533 557504 350538 557560
rect 350594 557504 350948 557560
rect 350533 557502 350948 557504
rect 350533 557499 350599 557502
rect 350942 557500 350948 557502
rect 351012 557500 351018 557564
rect 353293 557562 353359 557565
rect 354438 557562 354444 557564
rect 353293 557560 354444 557562
rect 353293 557504 353298 557560
rect 353354 557504 354444 557560
rect 353293 557502 354444 557504
rect 353293 557499 353359 557502
rect 354438 557500 354444 557502
rect 354508 557500 354514 557564
rect 354673 557562 354739 557565
rect 355726 557562 355732 557564
rect 354673 557560 355732 557562
rect 354673 557504 354678 557560
rect 354734 557504 355732 557560
rect 354673 557502 355732 557504
rect 354673 557499 354739 557502
rect 355726 557500 355732 557502
rect 355796 557500 355802 557564
rect 356053 557562 356119 557565
rect 356646 557562 356652 557564
rect 356053 557560 356652 557562
rect 356053 557504 356058 557560
rect 356114 557504 356652 557560
rect 356053 557502 356652 557504
rect 356053 557499 356119 557502
rect 356646 557500 356652 557502
rect 356716 557500 356722 557564
rect 357525 557562 357591 557565
rect 357934 557562 357940 557564
rect 357525 557560 357940 557562
rect 357525 557504 357530 557560
rect 357586 557504 357940 557560
rect 357525 557502 357940 557504
rect 357525 557499 357591 557502
rect 357934 557500 357940 557502
rect 358004 557500 358010 557564
rect 452653 557562 452719 557565
rect 452878 557562 452884 557564
rect 452653 557560 452884 557562
rect 452653 557504 452658 557560
rect 452714 557504 452884 557560
rect 452653 557502 452884 557504
rect 452653 557499 452719 557502
rect 452878 557500 452884 557502
rect 452948 557500 452954 557564
rect 453389 557562 453455 557565
rect 455270 557562 455276 557564
rect 453389 557560 455276 557562
rect 453389 557504 453394 557560
rect 453450 557504 455276 557560
rect 453389 557502 455276 557504
rect 453389 557499 453455 557502
rect 455270 557500 455276 557502
rect 455340 557500 455346 557564
rect 455413 557562 455479 557565
rect 456558 557562 456564 557564
rect 455413 557560 456564 557562
rect 455413 557504 455418 557560
rect 455474 557504 456564 557560
rect 455413 557502 456564 557504
rect 455413 557499 455479 557502
rect 456558 557500 456564 557502
rect 456628 557500 456634 557564
rect 456793 557562 456859 557565
rect 457478 557562 457484 557564
rect 456793 557560 457484 557562
rect 456793 557504 456798 557560
rect 456854 557504 457484 557560
rect 456793 557502 457484 557504
rect 456793 557499 456859 557502
rect 457478 557500 457484 557502
rect 457548 557500 457554 557564
rect 458173 557562 458239 557565
rect 458766 557562 458772 557564
rect 458173 557560 458772 557562
rect 458173 557504 458178 557560
rect 458234 557504 458772 557560
rect 458173 557502 458772 557504
rect 458173 557499 458239 557502
rect 458766 557500 458772 557502
rect 458836 557500 458842 557564
rect 459553 557562 459619 557565
rect 460933 557564 460999 557565
rect 460054 557562 460060 557564
rect 459553 557560 460060 557562
rect 459553 557504 459558 557560
rect 459614 557504 460060 557560
rect 459553 557502 460060 557504
rect 459553 557499 459619 557502
rect 460054 557500 460060 557502
rect 460124 557500 460130 557564
rect 460933 557562 460980 557564
rect 460888 557560 460980 557562
rect 460888 557504 460938 557560
rect 460888 557502 460980 557504
rect 460933 557500 460980 557502
rect 461044 557500 461050 557564
rect 462313 557562 462379 557565
rect 463550 557562 463556 557564
rect 462313 557560 463556 557562
rect 462313 557504 462318 557560
rect 462374 557504 463556 557560
rect 462313 557502 463556 557504
rect 460933 557499 460999 557500
rect 462313 557499 462379 557502
rect 463550 557500 463556 557502
rect 463620 557500 463626 557564
rect 463693 557562 463759 557565
rect 464470 557562 464476 557564
rect 463693 557560 464476 557562
rect 463693 557504 463698 557560
rect 463754 557504 464476 557560
rect 463693 557502 464476 557504
rect 463693 557499 463759 557502
rect 464470 557500 464476 557502
rect 464540 557500 464546 557564
rect 465073 557562 465139 557565
rect 465758 557562 465764 557564
rect 465073 557560 465764 557562
rect 465073 557504 465078 557560
rect 465134 557504 465764 557560
rect 465073 557502 465764 557504
rect 465073 557499 465139 557502
rect 465758 557500 465764 557502
rect 465828 557500 465834 557564
rect 474641 557562 474707 557565
rect 476389 557562 476455 557565
rect 474641 557560 476455 557562
rect 474641 557504 474646 557560
rect 474702 557504 476394 557560
rect 476450 557504 476455 557560
rect 474641 557502 476455 557504
rect 474641 557499 474707 557502
rect 476389 557499 476455 557502
rect 583520 557140 584960 557380
rect 352189 555524 352255 555525
rect 352189 555522 352236 555524
rect 352144 555520 352236 555522
rect 352144 555464 352194 555520
rect 352144 555462 352236 555464
rect 352189 555460 352236 555462
rect 352300 555460 352306 555524
rect 358905 555522 358971 555525
rect 359222 555522 359228 555524
rect 358905 555520 359228 555522
rect 358905 555464 358910 555520
rect 358966 555464 359228 555520
rect 358905 555462 359228 555464
rect 352189 555459 352255 555460
rect 358905 555459 358971 555462
rect 359222 555460 359228 555462
rect 359292 555460 359298 555524
rect -960 552924 480 553164
rect 583520 545444 584960 545684
rect 140037 543690 140103 543693
rect 200021 543690 200087 543693
rect 140037 543688 200087 543690
rect 140037 543632 140042 543688
rect 140098 543632 200026 543688
rect 200082 543632 200087 543688
rect 140037 543630 200087 543632
rect 140037 543627 140103 543630
rect 200021 543627 200087 543630
rect 148317 543554 148383 543557
rect 210417 543554 210483 543557
rect 148317 543552 210483 543554
rect 148317 543496 148322 543552
rect 148378 543496 210422 543552
rect 210478 543496 210483 543552
rect 148317 543494 210483 543496
rect 148317 543491 148383 543494
rect 210417 543491 210483 543494
rect 141417 543418 141483 543421
rect 208301 543418 208367 543421
rect 141417 543416 208367 543418
rect 141417 543360 141422 543416
rect 141478 543360 208306 543416
rect 208362 543360 208367 543416
rect 141417 543358 208367 543360
rect 141417 543355 141483 543358
rect 208301 543355 208367 543358
rect 96245 543282 96311 543285
rect 188337 543282 188403 543285
rect 96245 543280 188403 543282
rect 96245 543224 96250 543280
rect 96306 543224 188342 543280
rect 188398 543224 188403 543280
rect 96245 543222 188403 543224
rect 96245 543219 96311 543222
rect 188337 543219 188403 543222
rect 103421 543146 103487 543149
rect 202045 543146 202111 543149
rect 103421 543144 202111 543146
rect 103421 543088 103426 543144
rect 103482 543088 202050 543144
rect 202106 543088 202111 543144
rect 103421 543086 202111 543088
rect 103421 543083 103487 543086
rect 202045 543083 202111 543086
rect 77569 543010 77635 543013
rect 188981 543010 189047 543013
rect 77569 543008 189047 543010
rect 77569 542952 77574 543008
rect 77630 542952 188986 543008
rect 189042 542952 189047 543008
rect 77569 542950 189047 542952
rect 77569 542947 77635 542950
rect 188981 542947 189047 542950
rect 281717 539066 281783 539069
rect 279956 539064 281783 539066
rect 279956 539008 281722 539064
rect 281778 539008 281783 539064
rect 279956 539006 281783 539008
rect 281717 539003 281783 539006
rect -960 538508 480 538748
rect 281717 537026 281783 537029
rect 279956 537024 281783 537026
rect 279956 536968 281722 537024
rect 281778 536968 281783 537024
rect 279956 536966 281783 536968
rect 281717 536963 281783 536966
rect 281717 534986 281783 534989
rect 279956 534984 281783 534986
rect 279956 534928 281722 534984
rect 281778 534928 281783 534984
rect 279956 534926 281783 534928
rect 281717 534923 281783 534926
rect 583520 533748 584960 533988
rect 281717 532946 281783 532949
rect 279956 532944 281783 532946
rect 279956 532888 281722 532944
rect 281778 532888 281783 532944
rect 279956 532886 281783 532888
rect 281717 532883 281783 532886
rect 281717 530906 281783 530909
rect 279956 530904 281783 530906
rect 279956 530848 281722 530904
rect 281778 530848 281783 530904
rect 279956 530846 281783 530848
rect 281717 530843 281783 530846
rect 281717 528866 281783 528869
rect 279956 528864 281783 528866
rect 279956 528808 281722 528864
rect 281778 528808 281783 528864
rect 279956 528806 281783 528808
rect 281717 528803 281783 528806
rect 281717 526826 281783 526829
rect 279956 526824 281783 526826
rect 279956 526768 281722 526824
rect 281778 526768 281783 526824
rect 279956 526766 281783 526768
rect 281717 526763 281783 526766
rect 281717 524786 281783 524789
rect 279956 524784 281783 524786
rect 279956 524728 281722 524784
rect 281778 524728 281783 524784
rect 279956 524726 281783 524728
rect 281717 524723 281783 524726
rect -960 524092 480 524332
rect 281717 522746 281783 522749
rect 279956 522744 281783 522746
rect 279956 522688 281722 522744
rect 281778 522688 281783 522744
rect 279956 522686 281783 522688
rect 281717 522683 281783 522686
rect 583520 521916 584960 522156
rect 281717 520706 281783 520709
rect 279956 520704 281783 520706
rect 279956 520648 281722 520704
rect 281778 520648 281783 520704
rect 279956 520646 281783 520648
rect 281717 520643 281783 520646
rect 281717 518666 281783 518669
rect 279956 518664 281783 518666
rect 279956 518608 281722 518664
rect 281778 518608 281783 518664
rect 279956 518606 281783 518608
rect 281717 518603 281783 518606
rect 281717 516626 281783 516629
rect 279956 516624 281783 516626
rect 279956 516568 281722 516624
rect 281778 516568 281783 516624
rect 279956 516566 281783 516568
rect 281717 516563 281783 516566
rect 281717 514586 281783 514589
rect 279956 514584 281783 514586
rect 279956 514528 281722 514584
rect 281778 514528 281783 514584
rect 279956 514526 281783 514528
rect 281717 514523 281783 514526
rect 281717 512546 281783 512549
rect 279956 512544 281783 512546
rect 279956 512488 281722 512544
rect 281778 512488 281783 512544
rect 279956 512486 281783 512488
rect 281717 512483 281783 512486
rect 281717 510506 281783 510509
rect 279956 510504 281783 510506
rect 279956 510448 281722 510504
rect 281778 510448 281783 510504
rect 279956 510446 281783 510448
rect 281717 510443 281783 510446
rect 583520 510220 584960 510460
rect -960 509812 480 510052
rect 281717 508466 281783 508469
rect 279956 508464 281783 508466
rect 279956 508408 281722 508464
rect 281778 508408 281783 508464
rect 279956 508406 281783 508408
rect 281717 508403 281783 508406
rect 281717 506426 281783 506429
rect 279956 506424 281783 506426
rect 279956 506368 281722 506424
rect 281778 506368 281783 506424
rect 279956 506366 281783 506368
rect 281717 506363 281783 506366
rect 281717 504386 281783 504389
rect 279956 504384 281783 504386
rect 279956 504328 281722 504384
rect 281778 504328 281783 504384
rect 279956 504326 281783 504328
rect 281717 504323 281783 504326
rect 281717 502346 281783 502349
rect 279956 502344 281783 502346
rect 279956 502288 281722 502344
rect 281778 502288 281783 502344
rect 279956 502286 281783 502288
rect 281717 502283 281783 502286
rect 281717 500306 281783 500309
rect 279956 500304 281783 500306
rect 279956 500248 281722 500304
rect 281778 500248 281783 500304
rect 279956 500246 281783 500248
rect 281717 500243 281783 500246
rect 583520 498524 584960 498764
rect 281717 498266 281783 498269
rect 279956 498264 281783 498266
rect 279956 498208 281722 498264
rect 281778 498208 281783 498264
rect 279956 498206 281783 498208
rect 281717 498203 281783 498206
rect 281717 496226 281783 496229
rect 279956 496224 281783 496226
rect 279956 496168 281722 496224
rect 281778 496168 281783 496224
rect 279956 496166 281783 496168
rect 281717 496163 281783 496166
rect -960 495396 480 495636
rect 281717 494186 281783 494189
rect 279956 494184 281783 494186
rect 279956 494128 281722 494184
rect 281778 494128 281783 494184
rect 279956 494126 281783 494128
rect 281717 494123 281783 494126
rect 281717 492146 281783 492149
rect 279956 492144 281783 492146
rect 279956 492088 281722 492144
rect 281778 492088 281783 492144
rect 279956 492086 281783 492088
rect 281717 492083 281783 492086
rect 281717 490106 281783 490109
rect 279956 490104 281783 490106
rect 279956 490048 281722 490104
rect 281778 490048 281783 490104
rect 279956 490046 281783 490048
rect 281717 490043 281783 490046
rect 281717 488066 281783 488069
rect 279956 488064 281783 488066
rect 279956 488008 281722 488064
rect 281778 488008 281783 488064
rect 279956 488006 281783 488008
rect 281717 488003 281783 488006
rect 583520 486692 584960 486932
rect 281717 486026 281783 486029
rect 279956 486024 281783 486026
rect 279956 485968 281722 486024
rect 281778 485968 281783 486024
rect 279956 485966 281783 485968
rect 281717 485963 281783 485966
rect 281717 483986 281783 483989
rect 279956 483984 281783 483986
rect 279956 483928 281722 483984
rect 281778 483928 281783 483984
rect 279956 483926 281783 483928
rect 281717 483923 281783 483926
rect 281717 481946 281783 481949
rect 279956 481944 281783 481946
rect 279956 481888 281722 481944
rect 281778 481888 281783 481944
rect 279956 481886 281783 481888
rect 281717 481883 281783 481886
rect -960 480980 480 481220
rect 281717 479906 281783 479909
rect 279956 479904 281783 479906
rect 279956 479848 281722 479904
rect 281778 479848 281783 479904
rect 279956 479846 281783 479848
rect 281717 479843 281783 479846
rect 281717 477866 281783 477869
rect 279956 477864 281783 477866
rect 279956 477808 281722 477864
rect 281778 477808 281783 477864
rect 279956 477806 281783 477808
rect 281717 477803 281783 477806
rect 281717 475826 281783 475829
rect 279956 475824 281783 475826
rect 279956 475768 281722 475824
rect 281778 475768 281783 475824
rect 279956 475766 281783 475768
rect 281717 475763 281783 475766
rect 583520 474996 584960 475236
rect 281717 473786 281783 473789
rect 279956 473784 281783 473786
rect 279956 473728 281722 473784
rect 281778 473728 281783 473784
rect 279956 473726 281783 473728
rect 281717 473723 281783 473726
rect 281717 471746 281783 471749
rect 279956 471744 281783 471746
rect 279956 471688 281722 471744
rect 281778 471688 281783 471744
rect 279956 471686 281783 471688
rect 281717 471683 281783 471686
rect 281717 469706 281783 469709
rect 279956 469704 281783 469706
rect 279956 469648 281722 469704
rect 281778 469648 281783 469704
rect 279956 469646 281783 469648
rect 281717 469643 281783 469646
rect 281717 467666 281783 467669
rect 279956 467664 281783 467666
rect 279956 467608 281722 467664
rect 281778 467608 281783 467664
rect 279956 467606 281783 467608
rect 281717 467603 281783 467606
rect -960 466700 480 466940
rect 281717 465626 281783 465629
rect 279956 465624 281783 465626
rect 279956 465568 281722 465624
rect 281778 465568 281783 465624
rect 279956 465566 281783 465568
rect 281717 465563 281783 465566
rect 281717 463586 281783 463589
rect 279956 463584 281783 463586
rect 279956 463528 281722 463584
rect 281778 463528 281783 463584
rect 279956 463526 281783 463528
rect 281717 463523 281783 463526
rect 583520 463300 584960 463540
rect 281717 461546 281783 461549
rect 279956 461544 281783 461546
rect 279956 461488 281722 461544
rect 281778 461488 281783 461544
rect 279956 461486 281783 461488
rect 281717 461483 281783 461486
rect 281717 459506 281783 459509
rect 279956 459504 281783 459506
rect 279956 459448 281722 459504
rect 281778 459448 281783 459504
rect 279956 459446 281783 459448
rect 281717 459443 281783 459446
rect 281717 457466 281783 457469
rect 279956 457464 281783 457466
rect 279956 457408 281722 457464
rect 281778 457408 281783 457464
rect 279956 457406 281783 457408
rect 281717 457403 281783 457406
rect 281717 455426 281783 455429
rect 279956 455424 281783 455426
rect 279956 455368 281722 455424
rect 281778 455368 281783 455424
rect 279956 455366 281783 455368
rect 281717 455363 281783 455366
rect 281717 453386 281783 453389
rect 279956 453384 281783 453386
rect 279956 453328 281722 453384
rect 281778 453328 281783 453384
rect 279956 453326 281783 453328
rect 281717 453323 281783 453326
rect -960 452284 480 452524
rect 583520 451604 584960 451844
rect 281717 451346 281783 451349
rect 279956 451344 281783 451346
rect 279956 451288 281722 451344
rect 281778 451288 281783 451344
rect 279956 451286 281783 451288
rect 281717 451283 281783 451286
rect 281717 449306 281783 449309
rect 279956 449304 281783 449306
rect 279956 449248 281722 449304
rect 281778 449248 281783 449304
rect 279956 449246 281783 449248
rect 281717 449243 281783 449246
rect 281717 447266 281783 447269
rect 279956 447264 281783 447266
rect 279956 447208 281722 447264
rect 281778 447208 281783 447264
rect 279956 447206 281783 447208
rect 281717 447203 281783 447206
rect 281717 445226 281783 445229
rect 279956 445224 281783 445226
rect 279956 445168 281722 445224
rect 281778 445168 281783 445224
rect 279956 445166 281783 445168
rect 281717 445163 281783 445166
rect 281717 443186 281783 443189
rect 279956 443184 281783 443186
rect 279956 443128 281722 443184
rect 281778 443128 281783 443184
rect 279956 443126 281783 443128
rect 281717 443123 281783 443126
rect 281717 441146 281783 441149
rect 279956 441144 281783 441146
rect 279956 441088 281722 441144
rect 281778 441088 281783 441144
rect 279956 441086 281783 441088
rect 281717 441083 281783 441086
rect 583520 439772 584960 440012
rect 281717 439106 281783 439109
rect 279956 439104 281783 439106
rect 279956 439048 281722 439104
rect 281778 439048 281783 439104
rect 279956 439046 281783 439048
rect 281717 439043 281783 439046
rect -960 437868 480 438108
rect 281717 437066 281783 437069
rect 279956 437064 281783 437066
rect 279956 437008 281722 437064
rect 281778 437008 281783 437064
rect 279956 437006 281783 437008
rect 281717 437003 281783 437006
rect 281717 435026 281783 435029
rect 279956 435024 281783 435026
rect 279956 434968 281722 435024
rect 281778 434968 281783 435024
rect 279956 434966 281783 434968
rect 281717 434963 281783 434966
rect 281717 432986 281783 432989
rect 279956 432984 281783 432986
rect 279956 432928 281722 432984
rect 281778 432928 281783 432984
rect 279956 432926 281783 432928
rect 281717 432923 281783 432926
rect 281717 431082 281783 431085
rect 279956 431080 281783 431082
rect 279956 431024 281722 431080
rect 281778 431024 281783 431080
rect 279956 431022 281783 431024
rect 281717 431019 281783 431022
rect 281717 429042 281783 429045
rect 279956 429040 281783 429042
rect 279956 428984 281722 429040
rect 281778 428984 281783 429040
rect 279956 428982 281783 428984
rect 281717 428979 281783 428982
rect 583520 428076 584960 428316
rect 281717 427002 281783 427005
rect 279956 427000 281783 427002
rect 279956 426944 281722 427000
rect 281778 426944 281783 427000
rect 279956 426942 281783 426944
rect 281717 426939 281783 426942
rect 281717 424962 281783 424965
rect 279956 424960 281783 424962
rect 279956 424904 281722 424960
rect 281778 424904 281783 424960
rect 279956 424902 281783 424904
rect 281717 424899 281783 424902
rect -960 423588 480 423828
rect 281717 422922 281783 422925
rect 279956 422920 281783 422922
rect 279956 422864 281722 422920
rect 281778 422864 281783 422920
rect 279956 422862 281783 422864
rect 281717 422859 281783 422862
rect 281717 420882 281783 420885
rect 279956 420880 281783 420882
rect 279956 420824 281722 420880
rect 281778 420824 281783 420880
rect 279956 420822 281783 420824
rect 281717 420819 281783 420822
rect 281717 418842 281783 418845
rect 279956 418840 281783 418842
rect 279956 418784 281722 418840
rect 281778 418784 281783 418840
rect 279956 418782 281783 418784
rect 281717 418779 281783 418782
rect 281717 416802 281783 416805
rect 279956 416800 281783 416802
rect 279956 416744 281722 416800
rect 281778 416744 281783 416800
rect 279956 416742 281783 416744
rect 281717 416739 281783 416742
rect 583520 416380 584960 416620
rect 281717 414762 281783 414765
rect 279956 414760 281783 414762
rect 279956 414704 281722 414760
rect 281778 414704 281783 414760
rect 279956 414702 281783 414704
rect 281717 414699 281783 414702
rect 383561 413268 383627 413269
rect 383510 413266 383516 413268
rect 383470 413206 383516 413266
rect 383580 413264 383627 413268
rect 383622 413208 383627 413264
rect 383510 413204 383516 413206
rect 383580 413204 383627 413208
rect 383561 413203 383627 413204
rect 281717 412722 281783 412725
rect 513373 412724 513439 412725
rect 513373 412722 513420 412724
rect 279956 412720 281783 412722
rect 279956 412664 281722 412720
rect 281778 412664 281783 412720
rect 279956 412662 281783 412664
rect 513328 412720 513420 412722
rect 513328 412664 513378 412720
rect 513328 412662 513420 412664
rect 281717 412659 281783 412662
rect 513373 412660 513420 412662
rect 513484 412660 513490 412724
rect 513373 412659 513439 412660
rect 281993 410682 282059 410685
rect 279956 410680 282059 410682
rect 279956 410624 281998 410680
rect 282054 410624 282059 410680
rect 279956 410622 282059 410624
rect 281993 410619 282059 410622
rect -960 409172 480 409412
rect 281809 408642 281875 408645
rect 279956 408640 281875 408642
rect 279956 408584 281814 408640
rect 281870 408584 281875 408640
rect 279956 408582 281875 408584
rect 281809 408579 281875 408582
rect 281901 406602 281967 406605
rect 279956 406600 281967 406602
rect 279956 406544 281906 406600
rect 281962 406544 281967 406600
rect 279956 406542 281967 406544
rect 281901 406539 281967 406542
rect 583520 404684 584960 404924
rect 281717 404562 281783 404565
rect 279956 404560 281783 404562
rect 279956 404504 281722 404560
rect 281778 404504 281783 404560
rect 279956 404502 281783 404504
rect 281717 404499 281783 404502
rect 281533 402522 281599 402525
rect 279956 402520 281599 402522
rect 279956 402464 281538 402520
rect 281594 402464 281599 402520
rect 279956 402462 281599 402464
rect 281533 402459 281599 402462
rect 281625 400482 281691 400485
rect 279956 400480 281691 400482
rect 279956 400424 281630 400480
rect 281686 400424 281691 400480
rect 279956 400422 281691 400424
rect 281625 400419 281691 400422
rect 281717 398442 281783 398445
rect 279956 398440 281783 398442
rect 279956 398384 281722 398440
rect 281778 398384 281783 398440
rect 279956 398382 281783 398384
rect 281717 398379 281783 398382
rect 281533 396402 281599 396405
rect 279956 396400 281599 396402
rect 279956 396344 281538 396400
rect 281594 396344 281599 396400
rect 279956 396342 281599 396344
rect 281533 396339 281599 396342
rect -960 394892 480 395132
rect 282085 394362 282151 394365
rect 279956 394360 282151 394362
rect 279956 394304 282090 394360
rect 282146 394304 282151 394360
rect 279956 394302 282151 394304
rect 282085 394299 282151 394302
rect 583520 392852 584960 393092
rect 282821 392322 282887 392325
rect 279956 392320 282887 392322
rect 279956 392264 282826 392320
rect 282882 392264 282887 392320
rect 279956 392262 282887 392264
rect 282821 392259 282887 392262
rect 282729 390282 282795 390285
rect 279956 390280 282795 390282
rect 279956 390224 282734 390280
rect 282790 390224 282795 390280
rect 279956 390222 282795 390224
rect 282729 390219 282795 390222
rect 282637 388242 282703 388245
rect 279956 388240 282703 388242
rect 279956 388184 282642 388240
rect 282698 388184 282703 388240
rect 279956 388182 282703 388184
rect 282637 388179 282703 388182
rect 282545 386202 282611 386205
rect 279956 386200 282611 386202
rect 279956 386144 282550 386200
rect 282606 386144 282611 386200
rect 279956 386142 282611 386144
rect 282545 386139 282611 386142
rect 282453 384162 282519 384165
rect 279956 384160 282519 384162
rect 279956 384104 282458 384160
rect 282514 384104 282519 384160
rect 279956 384102 282519 384104
rect 282453 384099 282519 384102
rect 282361 382122 282427 382125
rect 279956 382120 282427 382122
rect 279956 382064 282366 382120
rect 282422 382064 282427 382120
rect 279956 382062 282427 382064
rect 282361 382059 282427 382062
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 282269 380082 282335 380085
rect 279956 380080 282335 380082
rect 279956 380024 282274 380080
rect 282330 380024 282335 380080
rect 279956 380022 282335 380024
rect 282269 380019 282335 380022
rect 281901 378042 281967 378045
rect 279956 378040 281967 378042
rect 279956 377984 281906 378040
rect 281962 377984 281967 378040
rect 279956 377982 281967 377984
rect 281901 377979 281967 377982
rect 282821 376002 282887 376005
rect 279956 376000 282887 376002
rect 279956 375944 282826 376000
rect 282882 375944 282887 376000
rect 279956 375942 282887 375944
rect 282821 375939 282887 375942
rect 282821 373962 282887 373965
rect 279956 373960 282887 373962
rect 279956 373904 282826 373960
rect 282882 373904 282887 373960
rect 279956 373902 282887 373904
rect 282821 373899 282887 373902
rect 282821 371922 282887 371925
rect 279956 371920 282887 371922
rect 279956 371864 282826 371920
rect 282882 371864 282887 371920
rect 279956 371862 282887 371864
rect 282821 371859 282887 371862
rect 282361 369882 282427 369885
rect 279956 369880 282427 369882
rect 279956 369824 282366 369880
rect 282422 369824 282427 369880
rect 279956 369822 282427 369824
rect 282361 369819 282427 369822
rect 583520 369460 584960 369700
rect 282269 367842 282335 367845
rect 279956 367840 282335 367842
rect 279956 367784 282274 367840
rect 282330 367784 282335 367840
rect 279956 367782 282335 367784
rect 282269 367779 282335 367782
rect -960 366060 480 366300
rect 281717 365802 281783 365805
rect 279956 365800 281783 365802
rect 279956 365744 281722 365800
rect 281778 365744 281783 365800
rect 279956 365742 281783 365744
rect 281717 365739 281783 365742
rect 282821 363762 282887 363765
rect 279956 363760 282887 363762
rect 279956 363704 282826 363760
rect 282882 363704 282887 363760
rect 279956 363702 282887 363704
rect 282821 363699 282887 363702
rect 281901 361722 281967 361725
rect 279956 361720 281967 361722
rect 279956 361664 281906 361720
rect 281962 361664 281967 361720
rect 279956 361662 281967 361664
rect 281901 361659 281967 361662
rect 281901 359682 281967 359685
rect 279956 359680 281967 359682
rect 279956 359624 281906 359680
rect 281962 359624 281967 359680
rect 279956 359622 281967 359624
rect 281901 359619 281967 359622
rect 583520 357764 584960 358004
rect 281717 357642 281783 357645
rect 279956 357640 281783 357642
rect 279956 357584 281722 357640
rect 281778 357584 281783 357640
rect 279956 357582 281783 357584
rect 281717 357579 281783 357582
rect 282085 355602 282151 355605
rect 279956 355600 282151 355602
rect 279956 355544 282090 355600
rect 282146 355544 282151 355600
rect 279956 355542 282151 355544
rect 282085 355539 282151 355542
rect 282821 353562 282887 353565
rect 279956 353560 282887 353562
rect 279956 353504 282826 353560
rect 282882 353504 282887 353560
rect 279956 353502 282887 353504
rect 282821 353499 282887 353502
rect -960 351780 480 352020
rect 282821 351522 282887 351525
rect 279956 351520 282887 351522
rect 279956 351464 282826 351520
rect 282882 351464 282887 351520
rect 279956 351462 282887 351464
rect 282821 351459 282887 351462
rect 282821 349482 282887 349485
rect 279956 349480 282887 349482
rect 279956 349424 282826 349480
rect 282882 349424 282887 349480
rect 279956 349422 282887 349424
rect 282821 349419 282887 349422
rect 282821 347714 282887 347717
rect 279926 347712 282887 347714
rect 279926 347656 282826 347712
rect 282882 347656 282887 347712
rect 279926 347654 282887 347656
rect 279926 347412 279986 347654
rect 282821 347651 282887 347654
rect 583520 345932 584960 346172
rect 281533 345402 281599 345405
rect 279956 345400 281599 345402
rect 279956 345344 281538 345400
rect 281594 345344 281599 345400
rect 279956 345342 281599 345344
rect 281533 345339 281599 345342
rect 282821 343362 282887 343365
rect 279956 343360 282887 343362
rect 279956 343304 282826 343360
rect 282882 343304 282887 343360
rect 279956 343302 282887 343304
rect 282821 343299 282887 343302
rect 281533 341322 281599 341325
rect 279956 341320 281599 341322
rect 279956 341264 281538 341320
rect 281594 341264 281599 341320
rect 279956 341262 281599 341264
rect 281533 341259 281599 341262
rect 281717 339282 281783 339285
rect 279956 339280 281783 339282
rect 279956 339224 281722 339280
rect 281778 339224 281783 339280
rect 279956 339222 281783 339224
rect 281717 339219 281783 339222
rect -960 337364 480 337604
rect 281533 337242 281599 337245
rect 279956 337240 281599 337242
rect 279956 337184 281538 337240
rect 281594 337184 281599 337240
rect 279956 337182 281599 337184
rect 281533 337179 281599 337182
rect 281625 335202 281691 335205
rect 279956 335200 281691 335202
rect 279956 335144 281630 335200
rect 281686 335144 281691 335200
rect 279956 335142 281691 335144
rect 281625 335139 281691 335142
rect 583520 334236 584960 334476
rect 281533 333162 281599 333165
rect 279956 333160 281599 333162
rect 279956 333104 281538 333160
rect 281594 333104 281599 333160
rect 279956 333102 281599 333104
rect 281533 333099 281599 333102
rect 281533 331122 281599 331125
rect 279956 331120 281599 331122
rect 279956 331064 281538 331120
rect 281594 331064 281599 331120
rect 279956 331062 281599 331064
rect 281533 331059 281599 331062
rect 281533 329082 281599 329085
rect 279956 329080 281599 329082
rect 279956 329024 281538 329080
rect 281594 329024 281599 329080
rect 279956 329022 281599 329024
rect 281533 329019 281599 329022
rect 281533 327042 281599 327045
rect 279956 327040 281599 327042
rect 279956 326984 281538 327040
rect 281594 326984 281599 327040
rect 279956 326982 281599 326984
rect 281533 326979 281599 326982
rect 281533 325002 281599 325005
rect 279956 325000 281599 325002
rect 279956 324944 281538 325000
rect 281594 324944 281599 325000
rect 279956 324942 281599 324944
rect 281533 324939 281599 324942
rect -960 322948 480 323188
rect 282310 322962 282316 322964
rect 279956 322902 282316 322962
rect 282310 322900 282316 322902
rect 282380 322900 282386 322964
rect 583520 322540 584960 322780
rect 282177 321058 282243 321061
rect 279956 321056 282243 321058
rect 279956 321000 282182 321056
rect 282238 321000 282243 321056
rect 279956 320998 282243 321000
rect 282177 320995 282243 320998
rect 313273 318746 313339 318749
rect 443085 318748 443151 318749
rect 313406 318746 313412 318748
rect 313273 318744 313412 318746
rect 313273 318688 313278 318744
rect 313334 318688 313412 318744
rect 313273 318686 313412 318688
rect 313273 318683 313339 318686
rect 313406 318684 313412 318686
rect 313476 318684 313482 318748
rect 443085 318744 443132 318748
rect 443196 318746 443202 318748
rect 443085 318688 443090 318744
rect 443085 318684 443132 318688
rect 443196 318686 443242 318746
rect 443196 318684 443202 318686
rect 443085 318683 443151 318684
rect 12341 318474 12407 318477
rect 64137 318474 64203 318477
rect 12341 318472 64203 318474
rect 12341 318416 12346 318472
rect 12402 318416 64142 318472
rect 64198 318416 64203 318472
rect 12341 318414 64203 318416
rect 12341 318411 12407 318414
rect 64137 318411 64203 318414
rect 144862 318412 144868 318476
rect 144932 318474 144938 318476
rect 149697 318474 149763 318477
rect 144932 318472 149763 318474
rect 144932 318416 149702 318472
rect 149758 318416 149763 318472
rect 144932 318414 149763 318416
rect 144932 318412 144938 318414
rect 149697 318411 149763 318414
rect 13629 318338 13695 318341
rect 65057 318338 65123 318341
rect 13629 318336 65123 318338
rect 13629 318280 13634 318336
rect 13690 318280 65062 318336
rect 65118 318280 65123 318336
rect 13629 318278 65123 318280
rect 13629 318275 13695 318278
rect 65057 318275 65123 318278
rect 279693 318338 279759 318341
rect 320766 318338 320772 318340
rect 279693 318336 320772 318338
rect 279693 318280 279698 318336
rect 279754 318280 320772 318336
rect 279693 318278 320772 318280
rect 279693 318275 279759 318278
rect 320766 318276 320772 318278
rect 320836 318276 320842 318340
rect 9581 318202 9647 318205
rect 63309 318202 63375 318205
rect 9581 318200 63375 318202
rect 9581 318144 9586 318200
rect 9642 318144 63314 318200
rect 63370 318144 63375 318200
rect 9581 318142 63375 318144
rect 9581 318139 9647 318142
rect 63309 318139 63375 318142
rect 136449 318202 136515 318205
rect 144862 318202 144868 318204
rect 136449 318200 144868 318202
rect 136449 318144 136454 318200
rect 136510 318144 144868 318200
rect 136449 318142 144868 318144
rect 136449 318139 136515 318142
rect 144862 318140 144868 318142
rect 144932 318140 144938 318204
rect 149697 318202 149763 318205
rect 157885 318202 157951 318205
rect 149697 318200 154498 318202
rect 149697 318144 149702 318200
rect 149758 318144 154498 318200
rect 149697 318142 154498 318144
rect 149697 318139 149763 318142
rect 154438 318100 154498 318142
rect 154622 318200 157951 318202
rect 154622 318144 157890 318200
rect 157946 318144 157951 318200
rect 154622 318142 157951 318144
rect 154622 318100 154682 318142
rect 157885 318139 157951 318142
rect 178677 318202 178743 318205
rect 311198 318202 311204 318204
rect 178677 318200 311204 318202
rect 178677 318144 178682 318200
rect 178738 318144 311204 318200
rect 178677 318142 311204 318144
rect 178677 318139 178743 318142
rect 311198 318140 311204 318142
rect 311268 318140 311274 318204
rect 5441 318066 5507 318069
rect 61929 318066 61995 318069
rect 5441 318064 61995 318066
rect 5441 318008 5446 318064
rect 5502 318008 61934 318064
rect 61990 318008 61995 318064
rect 154438 318040 154682 318100
rect 181345 318066 181411 318069
rect 321502 318066 321508 318068
rect 181345 318064 321508 318066
rect 5441 318006 61995 318008
rect 5441 318003 5507 318006
rect 61929 318003 61995 318006
rect 181345 318008 181350 318064
rect 181406 318008 321508 318064
rect 181345 318006 321508 318008
rect 181345 318003 181411 318006
rect 321502 318004 321508 318006
rect 321572 318004 321578 318068
rect 134609 317930 134675 317933
rect 137921 317930 137987 317933
rect 134609 317928 137987 317930
rect 134609 317872 134614 317928
rect 134670 317872 137926 317928
rect 137982 317872 137987 317928
rect 134609 317870 137987 317872
rect 134609 317867 134675 317870
rect 137921 317867 137987 317870
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 583520 299012 584960 299252
rect -960 294252 480 294492
rect 583520 287316 584960 287556
rect -960 279972 480 280212
rect 134977 280122 135043 280125
rect 135110 280122 135116 280124
rect 134977 280120 135116 280122
rect 134977 280064 134982 280120
rect 135038 280064 135116 280120
rect 134977 280062 135116 280064
rect 134977 280059 135043 280062
rect 135110 280060 135116 280062
rect 135180 280060 135186 280124
rect 74257 278762 74323 278765
rect 74441 278762 74507 278765
rect 74257 278760 74507 278762
rect 74257 278704 74262 278760
rect 74318 278704 74446 278760
rect 74502 278704 74507 278760
rect 74257 278702 74507 278704
rect 74257 278699 74323 278702
rect 74441 278699 74507 278702
rect 81709 278764 81775 278765
rect 81709 278760 81756 278764
rect 81820 278762 81826 278764
rect 81709 278704 81714 278760
rect 81709 278700 81756 278704
rect 81820 278702 81866 278762
rect 81820 278700 81826 278702
rect 81709 278699 81775 278700
rect 583520 275620 584960 275860
rect 134977 270602 135043 270605
rect 135110 270602 135116 270604
rect 134977 270600 135116 270602
rect 134977 270544 134982 270600
rect 135038 270544 135116 270600
rect 134977 270542 135116 270544
rect 134977 270539 135043 270542
rect 135110 270540 135116 270542
rect 135180 270540 135186 270604
rect 81750 270404 81756 270468
rect 81820 270466 81826 270468
rect 81893 270466 81959 270469
rect 81820 270464 81959 270466
rect 81820 270408 81898 270464
rect 81954 270408 81959 270464
rect 81820 270406 81959 270408
rect 81820 270404 81826 270406
rect 81893 270403 81959 270406
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 134977 260810 135043 260813
rect 135110 260810 135116 260812
rect 134977 260808 135116 260810
rect 134977 260752 134982 260808
rect 135038 260752 135116 260808
rect 134977 260750 135116 260752
rect 134977 260747 135043 260750
rect 135110 260748 135116 260750
rect 135180 260748 135186 260812
rect 74257 259450 74323 259453
rect 74441 259450 74507 259453
rect 74257 259448 74507 259450
rect 74257 259392 74262 259448
rect 74318 259392 74446 259448
rect 74502 259392 74507 259448
rect 74257 259390 74507 259392
rect 74257 259387 74323 259390
rect 74441 259387 74507 259390
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 134977 251290 135043 251293
rect 135110 251290 135116 251292
rect 134977 251288 135116 251290
rect 134977 251232 134982 251288
rect 135038 251232 135116 251288
rect 134977 251230 135116 251232
rect 134977 251227 135043 251230
rect 135110 251228 135116 251230
rect 135180 251228 135186 251292
rect 66345 241498 66411 241501
rect 66529 241498 66595 241501
rect 66345 241496 66595 241498
rect 66345 241440 66350 241496
rect 66406 241440 66534 241496
rect 66590 241440 66595 241496
rect 66345 241438 66595 241440
rect 66345 241435 66411 241438
rect 66529 241435 66595 241438
rect 72049 241498 72115 241501
rect 72233 241498 72299 241501
rect 72049 241496 72299 241498
rect 72049 241440 72054 241496
rect 72110 241440 72238 241496
rect 72294 241440 72299 241496
rect 72049 241438 72299 241440
rect 72049 241435 72115 241438
rect 72233 241435 72299 241438
rect 74809 241498 74875 241501
rect 74993 241498 75059 241501
rect 74809 241496 75059 241498
rect 74809 241440 74814 241496
rect 74870 241440 74998 241496
rect 75054 241440 75059 241496
rect 74809 241438 75059 241440
rect 74809 241435 74875 241438
rect 74993 241435 75059 241438
rect 95417 241498 95483 241501
rect 95601 241498 95667 241501
rect 95417 241496 95667 241498
rect 95417 241440 95422 241496
rect 95478 241440 95606 241496
rect 95662 241440 95667 241496
rect 95417 241438 95667 241440
rect 95417 241435 95483 241438
rect 95601 241435 95667 241438
rect 583520 240396 584960 240636
rect 74257 240138 74323 240141
rect 74441 240138 74507 240141
rect 74257 240136 74507 240138
rect 74257 240080 74262 240136
rect 74318 240080 74446 240136
rect 74502 240080 74507 240136
rect 74257 240078 74507 240080
rect 74257 240075 74323 240078
rect 74441 240075 74507 240078
rect -960 236860 480 237100
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 66345 222186 66411 222189
rect 66529 222186 66595 222189
rect 66345 222184 66595 222186
rect 66345 222128 66350 222184
rect 66406 222128 66534 222184
rect 66590 222128 66595 222184
rect 66345 222126 66595 222128
rect 66345 222123 66411 222126
rect 66529 222123 66595 222126
rect 72049 222186 72115 222189
rect 72233 222186 72299 222189
rect 72049 222184 72299 222186
rect 72049 222128 72054 222184
rect 72110 222128 72238 222184
rect 72294 222128 72299 222184
rect 72049 222126 72299 222128
rect 72049 222123 72115 222126
rect 72233 222123 72299 222126
rect 74809 222186 74875 222189
rect 74993 222186 75059 222189
rect 74809 222184 75059 222186
rect 74809 222128 74814 222184
rect 74870 222128 74998 222184
rect 75054 222128 75059 222184
rect 74809 222126 75059 222128
rect 74809 222123 74875 222126
rect 74993 222123 75059 222126
rect 77569 222186 77635 222189
rect 77753 222186 77819 222189
rect 77569 222184 77819 222186
rect 77569 222128 77574 222184
rect 77630 222128 77758 222184
rect 77814 222128 77819 222184
rect 77569 222126 77819 222128
rect 77569 222123 77635 222126
rect 77753 222123 77819 222126
rect 95417 222186 95483 222189
rect 95601 222186 95667 222189
rect 95417 222184 95667 222186
rect 95417 222128 95422 222184
rect 95478 222128 95606 222184
rect 95662 222128 95667 222184
rect 95417 222126 95667 222128
rect 95417 222123 95483 222126
rect 95601 222123 95667 222126
rect 74257 220826 74323 220829
rect 74441 220826 74507 220829
rect 74257 220824 74507 220826
rect 74257 220768 74262 220824
rect 74318 220768 74446 220824
rect 74502 220768 74507 220824
rect 74257 220766 74507 220768
rect 74257 220763 74323 220766
rect 74441 220763 74507 220766
rect 583520 216868 584960 217108
rect 85849 212530 85915 212533
rect 86125 212530 86191 212533
rect 85849 212528 86191 212530
rect 85849 212472 85854 212528
rect 85910 212472 86130 212528
rect 86186 212472 86191 212528
rect 85849 212470 86191 212472
rect 85849 212467 85915 212470
rect 86125 212467 86191 212470
rect 74257 211170 74323 211173
rect 74441 211170 74507 211173
rect 74257 211168 74507 211170
rect 74257 211112 74262 211168
rect 74318 211112 74446 211168
rect 74502 211112 74507 211168
rect 74257 211110 74507 211112
rect 74257 211107 74323 211110
rect 74441 211107 74507 211110
rect -960 208028 480 208268
rect 583520 205172 584960 205412
rect 66345 202874 66411 202877
rect 66529 202874 66595 202877
rect 66345 202872 66595 202874
rect 66345 202816 66350 202872
rect 66406 202816 66534 202872
rect 66590 202816 66595 202872
rect 66345 202814 66595 202816
rect 66345 202811 66411 202814
rect 66529 202811 66595 202814
rect 72049 202874 72115 202877
rect 72233 202874 72299 202877
rect 72049 202872 72299 202874
rect 72049 202816 72054 202872
rect 72110 202816 72238 202872
rect 72294 202816 72299 202872
rect 72049 202814 72299 202816
rect 72049 202811 72115 202814
rect 72233 202811 72299 202814
rect 74809 202874 74875 202877
rect 74993 202874 75059 202877
rect 74809 202872 75059 202874
rect 74809 202816 74814 202872
rect 74870 202816 74998 202872
rect 75054 202816 75059 202872
rect 74809 202814 75059 202816
rect 74809 202811 74875 202814
rect 74993 202811 75059 202814
rect 95417 202874 95483 202877
rect 95601 202874 95667 202877
rect 95417 202872 95667 202874
rect 95417 202816 95422 202872
rect 95478 202816 95606 202872
rect 95662 202816 95667 202872
rect 95417 202814 95667 202816
rect 95417 202811 95483 202814
rect 95601 202811 95667 202814
rect 160553 202874 160619 202877
rect 160737 202874 160803 202877
rect 160553 202872 160803 202874
rect 160553 202816 160558 202872
rect 160614 202816 160742 202872
rect 160798 202816 160803 202872
rect 160553 202814 160803 202816
rect 160553 202811 160619 202814
rect 160737 202811 160803 202814
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 85849 193218 85915 193221
rect 86125 193218 86191 193221
rect 85849 193216 86191 193218
rect 85849 193160 85854 193216
rect 85910 193160 86130 193216
rect 86186 193160 86191 193216
rect 85849 193158 86191 193160
rect 85849 193155 85915 193158
rect 86125 193155 86191 193158
rect 134793 193218 134859 193221
rect 134977 193218 135043 193221
rect 134793 193216 135043 193218
rect 134793 193160 134798 193216
rect 134854 193160 134982 193216
rect 135038 193160 135043 193216
rect 134793 193158 135043 193160
rect 134793 193155 134859 193158
rect 134977 193155 135043 193158
rect 74257 191858 74323 191861
rect 74441 191858 74507 191861
rect 74257 191856 74507 191858
rect 74257 191800 74262 191856
rect 74318 191800 74446 191856
rect 74502 191800 74507 191856
rect 74257 191798 74507 191800
rect 74257 191795 74323 191798
rect 74441 191795 74507 191798
rect 66345 183562 66411 183565
rect 66529 183562 66595 183565
rect 66345 183560 66595 183562
rect 66345 183504 66350 183560
rect 66406 183504 66534 183560
rect 66590 183504 66595 183560
rect 66345 183502 66595 183504
rect 66345 183499 66411 183502
rect 66529 183499 66595 183502
rect 72049 183562 72115 183565
rect 72233 183562 72299 183565
rect 72049 183560 72299 183562
rect 72049 183504 72054 183560
rect 72110 183504 72238 183560
rect 72294 183504 72299 183560
rect 72049 183502 72299 183504
rect 72049 183499 72115 183502
rect 72233 183499 72299 183502
rect 74809 183562 74875 183565
rect 74993 183562 75059 183565
rect 74809 183560 75059 183562
rect 74809 183504 74814 183560
rect 74870 183504 74998 183560
rect 75054 183504 75059 183560
rect 74809 183502 75059 183504
rect 74809 183499 74875 183502
rect 74993 183499 75059 183502
rect 95417 183562 95483 183565
rect 95601 183562 95667 183565
rect 95417 183560 95667 183562
rect 95417 183504 95422 183560
rect 95478 183504 95606 183560
rect 95662 183504 95667 183560
rect 95417 183502 95667 183504
rect 95417 183499 95483 183502
rect 95601 183499 95667 183502
rect 140865 183562 140931 183565
rect 141141 183562 141207 183565
rect 140865 183560 141207 183562
rect 140865 183504 140870 183560
rect 140926 183504 141146 183560
rect 141202 183504 141207 183560
rect 140865 183502 141207 183504
rect 140865 183499 140931 183502
rect 141141 183499 141207 183502
rect 150065 183562 150131 183565
rect 150249 183562 150315 183565
rect 150065 183560 150315 183562
rect 150065 183504 150070 183560
rect 150126 183504 150254 183560
rect 150310 183504 150315 183560
rect 150065 183502 150315 183504
rect 150065 183499 150131 183502
rect 150249 183499 150315 183502
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 134793 173906 134859 173909
rect 134977 173906 135043 173909
rect 134793 173904 135043 173906
rect 134793 173848 134798 173904
rect 134854 173848 134982 173904
rect 135038 173848 135043 173904
rect 134793 173846 135043 173848
rect 134793 173843 134859 173846
rect 134977 173843 135043 173846
rect 74257 172546 74323 172549
rect 74441 172546 74507 172549
rect 74257 172544 74507 172546
rect 74257 172488 74262 172544
rect 74318 172488 74446 172544
rect 74502 172488 74507 172544
rect 74257 172486 74507 172488
rect 74257 172483 74323 172486
rect 74441 172483 74507 172486
rect 583520 169948 584960 170188
rect -960 164916 480 165156
rect 583520 158252 584960 158492
rect 66345 154594 66411 154597
rect 66621 154594 66687 154597
rect 66345 154592 66687 154594
rect 66345 154536 66350 154592
rect 66406 154536 66626 154592
rect 66682 154536 66687 154592
rect 66345 154534 66687 154536
rect 66345 154531 66411 154534
rect 66621 154531 66687 154534
rect 95417 154594 95483 154597
rect 95693 154594 95759 154597
rect 95417 154592 95759 154594
rect 95417 154536 95422 154592
rect 95478 154536 95698 154592
rect 95754 154536 95759 154592
rect 95417 154534 95759 154536
rect 95417 154531 95483 154534
rect 95693 154531 95759 154534
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect 72233 145074 72299 145077
rect 74441 145074 74507 145077
rect 74993 145074 75059 145077
rect 72233 145072 72434 145074
rect 72233 145016 72238 145072
rect 72294 145016 72434 145072
rect 72233 145014 72434 145016
rect 72233 145011 72299 145014
rect 72233 144938 72299 144941
rect 72374 144938 72434 145014
rect 74441 145072 74642 145074
rect 74441 145016 74446 145072
rect 74502 145016 74642 145072
rect 74441 145014 74642 145016
rect 74441 145011 74507 145014
rect 72233 144936 72434 144938
rect 72233 144880 72238 144936
rect 72294 144880 72434 144936
rect 72233 144878 72434 144880
rect 74441 144938 74507 144941
rect 74582 144938 74642 145014
rect 74993 145072 75194 145074
rect 74993 145016 74998 145072
rect 75054 145016 75194 145072
rect 74993 145014 75194 145016
rect 74993 145011 75059 145014
rect 74441 144936 74642 144938
rect 74441 144880 74446 144936
rect 74502 144880 74642 144936
rect 74441 144878 74642 144880
rect 74993 144938 75059 144941
rect 75134 144938 75194 145014
rect 74993 144936 75194 144938
rect 74993 144880 74998 144936
rect 75054 144880 75194 144936
rect 74993 144878 75194 144880
rect 85941 144938 86007 144941
rect 86125 144938 86191 144941
rect 85941 144936 86191 144938
rect 85941 144880 85946 144936
rect 86002 144880 86130 144936
rect 86186 144880 86191 144936
rect 85941 144878 86191 144880
rect 72233 144875 72299 144878
rect 74441 144875 74507 144878
rect 74993 144875 75059 144878
rect 85941 144875 86007 144878
rect 86125 144875 86191 144878
rect 124305 144938 124371 144941
rect 124581 144938 124647 144941
rect 124305 144936 124647 144938
rect 124305 144880 124310 144936
rect 124366 144880 124586 144936
rect 124642 144880 124647 144936
rect 124305 144878 124647 144880
rect 124305 144875 124371 144878
rect 124581 144875 124647 144878
rect -960 136220 480 136460
rect 66345 135282 66411 135285
rect 66621 135282 66687 135285
rect 66345 135280 66687 135282
rect 66345 135224 66350 135280
rect 66406 135224 66626 135280
rect 66682 135224 66687 135280
rect 66345 135222 66687 135224
rect 66345 135219 66411 135222
rect 66621 135219 66687 135222
rect 85849 135282 85915 135285
rect 86033 135282 86099 135285
rect 85849 135280 86099 135282
rect 85849 135224 85854 135280
rect 85910 135224 86038 135280
rect 86094 135224 86099 135280
rect 85849 135222 86099 135224
rect 85849 135219 85915 135222
rect 86033 135219 86099 135222
rect 95417 135282 95483 135285
rect 95693 135282 95759 135285
rect 95417 135280 95759 135282
rect 95417 135224 95422 135280
rect 95478 135224 95698 135280
rect 95754 135224 95759 135280
rect 95417 135222 95759 135224
rect 95417 135219 95483 135222
rect 95693 135219 95759 135222
rect 583520 134724 584960 134964
rect 72233 125762 72299 125765
rect 74441 125762 74507 125765
rect 74993 125762 75059 125765
rect 78857 125762 78923 125765
rect 72233 125760 72434 125762
rect 72233 125704 72238 125760
rect 72294 125704 72434 125760
rect 72233 125702 72434 125704
rect 72233 125699 72299 125702
rect 72233 125626 72299 125629
rect 72374 125626 72434 125702
rect 74441 125760 74642 125762
rect 74441 125704 74446 125760
rect 74502 125704 74642 125760
rect 74441 125702 74642 125704
rect 74441 125699 74507 125702
rect 72233 125624 72434 125626
rect 72233 125568 72238 125624
rect 72294 125568 72434 125624
rect 72233 125566 72434 125568
rect 74441 125626 74507 125629
rect 74582 125626 74642 125702
rect 74993 125760 75194 125762
rect 74993 125704 74998 125760
rect 75054 125704 75194 125760
rect 74993 125702 75194 125704
rect 74993 125699 75059 125702
rect 74441 125624 74642 125626
rect 74441 125568 74446 125624
rect 74502 125568 74642 125624
rect 74441 125566 74642 125568
rect 74993 125626 75059 125629
rect 75134 125626 75194 125702
rect 78814 125760 78923 125762
rect 78814 125704 78862 125760
rect 78918 125704 78923 125760
rect 78814 125699 78923 125704
rect 78814 125629 78874 125699
rect 74993 125624 75194 125626
rect 74993 125568 74998 125624
rect 75054 125568 75194 125624
rect 74993 125566 75194 125568
rect 78765 125624 78874 125629
rect 78765 125568 78770 125624
rect 78826 125568 78874 125624
rect 78765 125566 78874 125568
rect 85941 125626 86007 125629
rect 86125 125626 86191 125629
rect 85941 125624 86191 125626
rect 85941 125568 85946 125624
rect 86002 125568 86130 125624
rect 86186 125568 86191 125624
rect 85941 125566 86191 125568
rect 72233 125563 72299 125566
rect 74441 125563 74507 125566
rect 74993 125563 75059 125566
rect 78765 125563 78831 125566
rect 85941 125563 86007 125566
rect 86125 125563 86191 125566
rect 124305 125626 124371 125629
rect 124581 125626 124647 125629
rect 124305 125624 124647 125626
rect 124305 125568 124310 125624
rect 124366 125568 124586 125624
rect 124642 125568 124647 125624
rect 124305 125566 124647 125568
rect 124305 125563 124371 125566
rect 124581 125563 124647 125566
rect 77477 124266 77543 124269
rect 77845 124266 77911 124269
rect 77477 124264 77911 124266
rect 77477 124208 77482 124264
rect 77538 124208 77850 124264
rect 77906 124208 77911 124264
rect 77477 124206 77911 124208
rect 77477 124203 77543 124206
rect 77845 124203 77911 124206
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 66345 115970 66411 115973
rect 66621 115970 66687 115973
rect 66345 115968 66687 115970
rect 66345 115912 66350 115968
rect 66406 115912 66626 115968
rect 66682 115912 66687 115968
rect 66345 115910 66687 115912
rect 66345 115907 66411 115910
rect 66621 115907 66687 115910
rect 85849 115970 85915 115973
rect 86033 115970 86099 115973
rect 85849 115968 86099 115970
rect 85849 115912 85854 115968
rect 85910 115912 86038 115968
rect 86094 115912 86099 115968
rect 85849 115910 86099 115912
rect 85849 115907 85915 115910
rect 86033 115907 86099 115910
rect 95417 115970 95483 115973
rect 95693 115970 95759 115973
rect 95417 115968 95759 115970
rect 95417 115912 95422 115968
rect 95478 115912 95698 115968
rect 95754 115912 95759 115968
rect 95417 115910 95759 115912
rect 95417 115907 95483 115910
rect 95693 115907 95759 115910
rect 583520 111332 584960 111572
rect -960 107524 480 107764
rect 78857 106450 78923 106453
rect 78814 106448 78923 106450
rect 78814 106392 78862 106448
rect 78918 106392 78923 106448
rect 78814 106387 78923 106392
rect 78814 106317 78874 106387
rect 78765 106312 78874 106317
rect 78765 106256 78770 106312
rect 78826 106256 78874 106312
rect 78765 106254 78874 106256
rect 124305 106314 124371 106317
rect 124581 106314 124647 106317
rect 124305 106312 124647 106314
rect 124305 106256 124310 106312
rect 124366 106256 124586 106312
rect 124642 106256 124647 106312
rect 124305 106254 124647 106256
rect 78765 106251 78831 106254
rect 124305 106251 124371 106254
rect 124581 106251 124647 106254
rect 583520 99636 584960 99876
rect 66345 96658 66411 96661
rect 66621 96658 66687 96661
rect 66345 96656 66687 96658
rect 66345 96600 66350 96656
rect 66406 96600 66626 96656
rect 66682 96600 66687 96656
rect 66345 96598 66687 96600
rect 66345 96595 66411 96598
rect 66621 96595 66687 96598
rect 95417 96658 95483 96661
rect 95693 96658 95759 96661
rect 95417 96656 95759 96658
rect 95417 96600 95422 96656
rect 95478 96600 95698 96656
rect 95754 96600 95759 96656
rect 95417 96598 95759 96600
rect 95417 96595 95483 96598
rect 95693 96595 95759 96598
rect -960 93108 480 93348
rect 583520 87804 584960 88044
rect 124305 87002 124371 87005
rect 124581 87002 124647 87005
rect 124305 87000 124647 87002
rect 124305 86944 124310 87000
rect 124366 86944 124586 87000
rect 124642 86944 124647 87000
rect 124305 86942 124647 86944
rect 124305 86939 124371 86942
rect 124581 86939 124647 86942
rect -960 78828 480 79068
rect 134701 77346 134767 77349
rect 134885 77346 134951 77349
rect 134701 77344 134951 77346
rect 134701 77288 134706 77344
rect 134762 77288 134890 77344
rect 134946 77288 134951 77344
rect 134701 77286 134951 77288
rect 134701 77283 134767 77286
rect 134885 77283 134951 77286
rect 150157 77210 150223 77213
rect 150341 77210 150407 77213
rect 150157 77208 150407 77210
rect 150157 77152 150162 77208
rect 150218 77152 150346 77208
rect 150402 77152 150407 77208
rect 150157 77150 150407 77152
rect 150157 77147 150223 77150
rect 150341 77147 150407 77150
rect 583520 76108 584960 76348
rect 134885 67824 134951 67829
rect 134885 67768 134890 67824
rect 134946 67768 134951 67824
rect 134885 67763 134951 67768
rect 134888 67693 134948 67763
rect 134885 67688 134951 67693
rect 134885 67632 134890 67688
rect 134946 67632 134951 67688
rect 134885 67627 134951 67632
rect -960 64412 480 64652
rect 583520 64412 584960 64652
rect 135069 61436 135135 61437
rect 135069 61434 135116 61436
rect 135024 61432 135116 61434
rect 135024 61376 135074 61432
rect 135024 61374 135116 61376
rect 135069 61372 135116 61374
rect 135180 61372 135186 61436
rect 135069 61371 135135 61372
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 134977 48378 135043 48381
rect 135110 48378 135116 48380
rect 134977 48376 135116 48378
rect 134977 48320 134982 48376
rect 135038 48320 135116 48376
rect 134977 48318 135116 48320
rect 134977 48315 135043 48318
rect 135110 48316 135116 48318
rect 135180 48316 135186 48380
rect 124489 42124 124555 42125
rect 124438 42060 124444 42124
rect 124508 42122 124555 42124
rect 135069 42124 135135 42125
rect 135069 42122 135116 42124
rect 124508 42120 124600 42122
rect 124550 42064 124600 42120
rect 124508 42062 124600 42064
rect 135024 42120 135116 42122
rect 135024 42064 135074 42120
rect 135024 42062 135116 42064
rect 124508 42060 124555 42062
rect 124489 42059 124555 42060
rect 135069 42060 135116 42062
rect 135180 42060 135186 42124
rect 135069 42059 135135 42060
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 124397 32468 124463 32469
rect 124397 32464 124444 32468
rect 124508 32466 124514 32468
rect 124397 32408 124402 32464
rect 124397 32404 124444 32408
rect 124508 32406 124554 32466
rect 124508 32404 124514 32406
rect 124397 32403 124463 32404
rect 583520 29188 584960 29428
rect 134977 29066 135043 29069
rect 135110 29066 135116 29068
rect 134977 29064 135116 29066
rect 134977 29008 134982 29064
rect 135038 29008 135116 29064
rect 134977 29006 135116 29008
rect 134977 29003 135043 29006
rect 135110 29004 135116 29006
rect 135180 29004 135186 29068
rect -960 21300 480 21540
rect 583520 17492 584960 17732
rect 250989 15058 251055 15061
rect 502333 15058 502399 15061
rect 250989 15056 502399 15058
rect 250989 15000 250994 15056
rect 251050 15000 502338 15056
rect 502394 15000 502399 15056
rect 250989 14998 502399 15000
rect 250989 14995 251055 14998
rect 502333 14995 502399 14998
rect 252369 14922 252435 14925
rect 506473 14922 506539 14925
rect 252369 14920 506539 14922
rect 252369 14864 252374 14920
rect 252430 14864 506478 14920
rect 506534 14864 506539 14920
rect 252369 14862 506539 14864
rect 252369 14859 252435 14862
rect 506473 14859 506539 14862
rect 253657 14786 253723 14789
rect 510613 14786 510679 14789
rect 253657 14784 510679 14786
rect 253657 14728 253662 14784
rect 253718 14728 510618 14784
rect 510674 14728 510679 14784
rect 253657 14726 510679 14728
rect 253657 14723 253723 14726
rect 510613 14723 510679 14726
rect 255037 14650 255103 14653
rect 513373 14650 513439 14653
rect 255037 14648 513439 14650
rect 255037 14592 255042 14648
rect 255098 14592 513378 14648
rect 513434 14592 513439 14648
rect 255037 14590 513439 14592
rect 255037 14587 255103 14590
rect 513373 14587 513439 14590
rect 266077 14514 266143 14517
rect 545113 14514 545179 14517
rect 266077 14512 545179 14514
rect 266077 14456 266082 14512
rect 266138 14456 545118 14512
rect 545174 14456 545179 14512
rect 266077 14454 545179 14456
rect 266077 14451 266143 14454
rect 545113 14451 545179 14454
rect 266169 13562 266235 13565
rect 546493 13562 546559 13565
rect 266169 13560 546559 13562
rect 266169 13504 266174 13560
rect 266230 13504 546498 13560
rect 546554 13504 546559 13560
rect 266169 13502 546559 13504
rect 266169 13499 266235 13502
rect 546493 13499 546559 13502
rect 267457 13426 267523 13429
rect 549253 13426 549319 13429
rect 267457 13424 549319 13426
rect 267457 13368 267462 13424
rect 267518 13368 549258 13424
rect 549314 13368 549319 13424
rect 267457 13366 549319 13368
rect 267457 13363 267523 13366
rect 549253 13363 549319 13366
rect 268837 13290 268903 13293
rect 553393 13290 553459 13293
rect 268837 13288 553459 13290
rect 268837 13232 268842 13288
rect 268898 13232 553398 13288
rect 553454 13232 553459 13288
rect 268837 13230 553459 13232
rect 268837 13227 268903 13230
rect 553393 13227 553459 13230
rect 270217 13154 270283 13157
rect 556153 13154 556219 13157
rect 270217 13152 556219 13154
rect 270217 13096 270222 13152
rect 270278 13096 556158 13152
rect 556214 13096 556219 13152
rect 270217 13094 556219 13096
rect 270217 13091 270283 13094
rect 556153 13091 556219 13094
rect 271597 13018 271663 13021
rect 560293 13018 560359 13021
rect 271597 13016 560359 13018
rect 271597 12960 271602 13016
rect 271658 12960 560298 13016
rect 560354 12960 560359 13016
rect 271597 12958 560359 12960
rect 271597 12955 271663 12958
rect 560293 12955 560359 12958
rect 244181 12202 244247 12205
rect 485865 12202 485931 12205
rect 244181 12200 485931 12202
rect 244181 12144 244186 12200
rect 244242 12144 485870 12200
rect 485926 12144 485931 12200
rect 244181 12142 485931 12144
rect 244181 12139 244247 12142
rect 485865 12139 485931 12142
rect 245561 12066 245627 12069
rect 488533 12066 488599 12069
rect 245561 12064 488599 12066
rect 245561 12008 245566 12064
rect 245622 12008 488538 12064
rect 488594 12008 488599 12064
rect 245561 12006 488599 12008
rect 245561 12003 245627 12006
rect 488533 12003 488599 12006
rect 246941 11930 247007 11933
rect 492673 11930 492739 11933
rect 246941 11928 492739 11930
rect 246941 11872 246946 11928
rect 247002 11872 492678 11928
rect 492734 11872 492739 11928
rect 246941 11870 492739 11872
rect 246941 11867 247007 11870
rect 492673 11867 492739 11870
rect 248229 11794 248295 11797
rect 495433 11794 495499 11797
rect 248229 11792 495499 11794
rect 248229 11736 248234 11792
rect 248290 11736 495438 11792
rect 495494 11736 495499 11792
rect 248229 11734 495499 11736
rect 248229 11731 248295 11734
rect 495433 11731 495499 11734
rect 249609 11658 249675 11661
rect 499573 11658 499639 11661
rect 249609 11656 499639 11658
rect 249609 11600 249614 11656
rect 249670 11600 499578 11656
rect 499634 11600 499639 11656
rect 249609 11598 499639 11600
rect 249609 11595 249675 11598
rect 499573 11595 499639 11598
rect 204069 10842 204135 10845
rect 380893 10842 380959 10845
rect 204069 10840 380959 10842
rect 204069 10784 204074 10840
rect 204130 10784 380898 10840
rect 380954 10784 380959 10840
rect 204069 10782 380959 10784
rect 204069 10779 204135 10782
rect 380893 10779 380959 10782
rect 205449 10706 205515 10709
rect 383653 10706 383719 10709
rect 205449 10704 383719 10706
rect 205449 10648 205454 10704
rect 205510 10648 383658 10704
rect 383714 10648 383719 10704
rect 205449 10646 383719 10648
rect 205449 10643 205515 10646
rect 383653 10643 383719 10646
rect 208301 10570 208367 10573
rect 390645 10570 390711 10573
rect 208301 10568 390711 10570
rect 208301 10512 208306 10568
rect 208362 10512 390650 10568
rect 390706 10512 390711 10568
rect 208301 10510 390711 10512
rect 208301 10507 208367 10510
rect 390645 10507 390711 10510
rect 209497 10434 209563 10437
rect 394693 10434 394759 10437
rect 209497 10432 394759 10434
rect 209497 10376 209502 10432
rect 209558 10376 394698 10432
rect 394754 10376 394759 10432
rect 209497 10374 394759 10376
rect 209497 10371 209563 10374
rect 394693 10371 394759 10374
rect 210969 10298 211035 10301
rect 398833 10298 398899 10301
rect 210969 10296 398899 10298
rect 210969 10240 210974 10296
rect 211030 10240 398838 10296
rect 398894 10240 398899 10296
rect 210969 10238 398899 10240
rect 210969 10235 211035 10238
rect 398833 10235 398899 10238
rect 260649 9618 260715 9621
rect 531037 9618 531103 9621
rect 260649 9616 531103 9618
rect 260649 9560 260654 9616
rect 260710 9560 531042 9616
rect 531098 9560 531103 9616
rect 260649 9558 531103 9560
rect 260649 9555 260715 9558
rect 531037 9555 531103 9558
rect 263409 9482 263475 9485
rect 538121 9482 538187 9485
rect 263409 9480 538187 9482
rect 263409 9424 263414 9480
rect 263470 9424 538126 9480
rect 538182 9424 538187 9480
rect 263409 9422 538187 9424
rect 263409 9419 263475 9422
rect 538121 9419 538187 9422
rect 267549 9346 267615 9349
rect 548885 9346 548951 9349
rect 267549 9344 548951 9346
rect 267549 9288 267554 9344
rect 267610 9288 548890 9344
rect 548946 9288 548951 9344
rect 267549 9286 548951 9288
rect 267549 9283 267615 9286
rect 548885 9283 548951 9286
rect 270309 9210 270375 9213
rect 555969 9210 556035 9213
rect 270309 9208 556035 9210
rect 270309 9152 270314 9208
rect 270370 9152 555974 9208
rect 556030 9152 556035 9208
rect 270309 9150 556035 9152
rect 270309 9147 270375 9150
rect 555969 9147 556035 9150
rect 275829 9074 275895 9077
rect 570229 9074 570295 9077
rect 275829 9072 570295 9074
rect 275829 9016 275834 9072
rect 275890 9016 570234 9072
rect 570290 9016 570295 9072
rect 275829 9014 570295 9016
rect 275829 9011 275895 9014
rect 570229 9011 570295 9014
rect 279969 8938 280035 8941
rect 580993 8938 581059 8941
rect 279969 8936 581059 8938
rect 279969 8880 279974 8936
rect 280030 8880 580998 8936
rect 581054 8880 581059 8936
rect 279969 8878 581059 8880
rect 279969 8875 280035 8878
rect 580993 8875 581059 8878
rect 235809 8258 235875 8261
rect 465625 8258 465691 8261
rect 235809 8256 465691 8258
rect 235809 8200 235814 8256
rect 235870 8200 465630 8256
rect 465686 8200 465691 8256
rect 235809 8198 465691 8200
rect 235809 8195 235875 8198
rect 465625 8195 465691 8198
rect 237281 8122 237347 8125
rect 469121 8122 469187 8125
rect 237281 8120 469187 8122
rect 237281 8064 237286 8120
rect 237342 8064 469126 8120
rect 469182 8064 469187 8120
rect 237281 8062 469187 8064
rect 237281 8059 237347 8062
rect 469121 8059 469187 8062
rect 238569 7986 238635 7989
rect 472709 7986 472775 7989
rect 238569 7984 472775 7986
rect 238569 7928 238574 7984
rect 238630 7928 472714 7984
rect 472770 7928 472775 7984
rect 238569 7926 472775 7928
rect 238569 7923 238635 7926
rect 472709 7923 472775 7926
rect 240041 7850 240107 7853
rect 476297 7850 476363 7853
rect 240041 7848 476363 7850
rect 240041 7792 240046 7848
rect 240102 7792 476302 7848
rect 476358 7792 476363 7848
rect 240041 7790 476363 7792
rect 240041 7787 240107 7790
rect 476297 7787 476363 7790
rect 241329 7714 241395 7717
rect 479885 7714 479951 7717
rect 241329 7712 479951 7714
rect 241329 7656 241334 7712
rect 241390 7656 479890 7712
rect 479946 7656 479951 7712
rect 241329 7654 479951 7656
rect 241329 7651 241395 7654
rect 479885 7651 479951 7654
rect 242801 7578 242867 7581
rect 484577 7578 484643 7581
rect 242801 7576 484643 7578
rect 242801 7520 242806 7576
rect 242862 7520 484582 7576
rect 484638 7520 484643 7576
rect 242801 7518 484643 7520
rect 242801 7515 242867 7518
rect 484577 7515 484643 7518
rect -960 7020 480 7260
rect 197169 6762 197235 6765
rect 362125 6762 362191 6765
rect 197169 6760 362191 6762
rect 197169 6704 197174 6760
rect 197230 6704 362130 6760
rect 362186 6704 362191 6760
rect 197169 6702 362191 6704
rect 197169 6699 197235 6702
rect 362125 6699 362191 6702
rect 198641 6626 198707 6629
rect 365805 6626 365871 6629
rect 198641 6624 365871 6626
rect 198641 6568 198646 6624
rect 198702 6568 365810 6624
rect 365866 6568 365871 6624
rect 198641 6566 365871 6568
rect 198641 6563 198707 6566
rect 365805 6563 365871 6566
rect 201401 6490 201467 6493
rect 372797 6490 372863 6493
rect 201401 6488 372863 6490
rect 201401 6432 201406 6488
rect 201462 6432 372802 6488
rect 372858 6432 372863 6488
rect 201401 6430 372863 6432
rect 201401 6427 201467 6430
rect 372797 6427 372863 6430
rect 204161 6354 204227 6357
rect 379973 6354 380039 6357
rect 204161 6352 380039 6354
rect 204161 6296 204166 6352
rect 204222 6296 379978 6352
rect 380034 6296 380039 6352
rect 204161 6294 380039 6296
rect 204161 6291 204227 6294
rect 379973 6291 380039 6294
rect 206829 6218 206895 6221
rect 387057 6218 387123 6221
rect 206829 6216 387123 6218
rect 206829 6160 206834 6216
rect 206890 6160 387062 6216
rect 387118 6160 387123 6216
rect 206829 6158 387123 6160
rect 206829 6155 206895 6158
rect 387057 6155 387123 6158
rect 583520 5796 584960 6036
rect 168281 5538 168347 5541
rect 283649 5538 283715 5541
rect 168281 5536 283715 5538
rect 168281 5480 168286 5536
rect 168342 5480 283654 5536
rect 283710 5480 283715 5536
rect 168281 5478 283715 5480
rect 168281 5475 168347 5478
rect 283649 5475 283715 5478
rect 169661 5402 169727 5405
rect 290733 5402 290799 5405
rect 169661 5400 290799 5402
rect 169661 5344 169666 5400
rect 169722 5344 290738 5400
rect 290794 5344 290799 5400
rect 169661 5342 290799 5344
rect 169661 5339 169727 5342
rect 290733 5339 290799 5342
rect 191649 5266 191715 5269
rect 347865 5266 347931 5269
rect 191649 5264 347931 5266
rect 191649 5208 191654 5264
rect 191710 5208 347870 5264
rect 347926 5208 347931 5264
rect 191649 5206 347931 5208
rect 191649 5203 191715 5206
rect 347865 5203 347931 5206
rect 164141 5130 164207 5133
rect 272885 5130 272951 5133
rect 164141 5128 272951 5130
rect 164141 5072 164146 5128
rect 164202 5072 272890 5128
rect 272946 5072 272951 5128
rect 164141 5070 272951 5072
rect 164141 5067 164207 5070
rect 272885 5067 272951 5070
rect 277301 5130 277367 5133
rect 572621 5130 572687 5133
rect 277301 5128 572687 5130
rect 277301 5072 277306 5128
rect 277362 5072 572626 5128
rect 572682 5072 572687 5128
rect 277301 5070 572687 5072
rect 277301 5067 277367 5070
rect 572621 5067 572687 5070
rect 165521 4994 165587 4997
rect 276473 4994 276539 4997
rect 165521 4992 276539 4994
rect 165521 4936 165526 4992
rect 165582 4936 276478 4992
rect 276534 4936 276539 4992
rect 165521 4934 276539 4936
rect 165521 4931 165587 4934
rect 276473 4931 276539 4934
rect 278681 4994 278747 4997
rect 576209 4994 576275 4997
rect 278681 4992 576275 4994
rect 278681 4936 278686 4992
rect 278742 4936 576214 4992
rect 576270 4936 576275 4992
rect 278681 4934 576275 4936
rect 278681 4931 278747 4934
rect 576209 4931 576275 4934
rect 166901 4856 166967 4861
rect 172329 4858 172395 4861
rect 166901 4800 166906 4856
rect 166962 4824 166967 4856
rect 167134 4856 172395 4858
rect 167134 4824 172334 4856
rect 166962 4800 172334 4824
rect 172390 4800 172395 4856
rect 166901 4798 172395 4800
rect 166901 4795 167194 4798
rect 172329 4795 172395 4798
rect 172513 4858 172579 4861
rect 180701 4858 180767 4861
rect 172513 4856 180767 4858
rect 172513 4800 172518 4856
rect 172574 4800 180706 4856
rect 180762 4800 180767 4856
rect 172513 4798 180767 4800
rect 172513 4795 172579 4798
rect 180701 4795 180767 4798
rect 182081 4858 182147 4861
rect 205449 4858 205515 4861
rect 212441 4858 212507 4861
rect 182081 4856 186192 4858
rect 182081 4800 182086 4856
rect 182142 4800 186192 4856
rect 182081 4798 186192 4800
rect 182081 4795 182147 4798
rect 166904 4764 167194 4795
rect 186132 4722 186192 4798
rect 205449 4856 212507 4858
rect 205449 4800 205454 4856
rect 205510 4800 212446 4856
rect 212502 4800 212507 4856
rect 205449 4798 212507 4800
rect 205449 4795 205515 4798
rect 212441 4795 212507 4798
rect 280061 4858 280127 4861
rect 579797 4858 579863 4861
rect 280061 4856 579863 4858
rect 280061 4800 280066 4856
rect 280122 4800 579802 4856
rect 579858 4800 579863 4856
rect 280061 4798 579863 4800
rect 280061 4795 280127 4798
rect 579797 4795 579863 4798
rect 186132 4662 193138 4722
rect 180701 4586 180767 4589
rect 182081 4586 182147 4589
rect 180701 4584 182147 4586
rect 180701 4528 180706 4584
rect 180762 4528 182086 4584
rect 182142 4528 182147 4584
rect 180701 4526 182147 4528
rect 180701 4523 180767 4526
rect 182081 4523 182147 4526
rect 193078 4450 193138 4662
rect 205449 4586 205515 4589
rect 202830 4584 205515 4586
rect 202830 4528 205454 4584
rect 205510 4528 205515 4584
rect 202830 4526 205515 4528
rect 202830 4450 202890 4526
rect 205449 4523 205515 4526
rect 212441 4586 212507 4589
rect 231761 4586 231827 4589
rect 234521 4586 234587 4589
rect 249742 4586 249748 4588
rect 212441 4584 215218 4586
rect 212441 4528 212446 4584
rect 212502 4528 215218 4584
rect 212441 4526 215218 4528
rect 212441 4523 212507 4526
rect 193078 4390 193322 4450
rect 176561 4314 176627 4317
rect 176745 4314 176811 4317
rect 176561 4312 176811 4314
rect 176561 4256 176566 4312
rect 176622 4256 176750 4312
rect 176806 4256 176811 4312
rect 176561 4254 176811 4256
rect 193262 4314 193322 4390
rect 196022 4390 202890 4450
rect 215158 4416 215218 4526
rect 231761 4584 234587 4586
rect 231761 4528 231766 4584
rect 231822 4528 234526 4584
rect 234582 4528 234587 4584
rect 231761 4526 234587 4528
rect 231761 4523 231827 4526
rect 234521 4523 234587 4526
rect 246254 4526 249748 4586
rect 222142 4450 222148 4452
rect 215342 4416 222148 4450
rect 215158 4390 222148 4416
rect 196022 4314 196082 4390
rect 215158 4356 215402 4390
rect 222142 4388 222148 4390
rect 222212 4388 222218 4452
rect 234705 4450 234771 4453
rect 244089 4450 244155 4453
rect 234705 4448 244155 4450
rect 234705 4392 234710 4448
rect 234766 4392 244094 4448
rect 244150 4392 244155 4448
rect 234705 4390 244155 4392
rect 234705 4387 234771 4390
rect 244089 4387 244155 4390
rect 244273 4450 244339 4453
rect 246254 4450 246314 4526
rect 249742 4524 249748 4526
rect 249812 4524 249818 4588
rect 259361 4586 259427 4589
rect 269062 4586 269068 4588
rect 259361 4584 269068 4586
rect 259361 4528 259366 4584
rect 259422 4528 269068 4584
rect 259361 4526 269068 4528
rect 259361 4523 259427 4526
rect 269062 4524 269068 4526
rect 269132 4524 269138 4588
rect 244273 4448 246314 4450
rect 244273 4392 244278 4448
rect 244334 4392 246314 4448
rect 244273 4390 246314 4392
rect 244273 4387 244339 4390
rect 193262 4254 196082 4314
rect 176561 4251 176627 4254
rect 176745 4251 176811 4254
rect 249742 4252 249748 4316
rect 249812 4314 249818 4316
rect 259361 4314 259427 4317
rect 249812 4312 259427 4314
rect 249812 4256 259366 4312
rect 259422 4256 259427 4312
rect 249812 4254 259427 4256
rect 249812 4252 249818 4254
rect 259361 4251 259427 4254
rect 269062 4252 269068 4316
rect 269132 4314 269138 4316
rect 273437 4314 273503 4317
rect 269132 4312 273503 4314
rect 269132 4256 273442 4312
rect 273498 4256 273503 4312
rect 269132 4254 273503 4256
rect 269132 4252 269138 4254
rect 273437 4251 273503 4254
rect 176469 4178 176535 4181
rect 176837 4178 176903 4181
rect 176469 4176 176903 4178
rect 176469 4120 176474 4176
rect 176530 4120 176842 4176
rect 176898 4120 176903 4176
rect 176469 4118 176903 4120
rect 176469 4115 176535 4118
rect 176837 4115 176903 4118
rect 178677 4178 178743 4181
rect 181529 4178 181595 4181
rect 178677 4176 181595 4178
rect 178677 4120 178682 4176
rect 178738 4120 181534 4176
rect 181590 4120 181595 4176
rect 178677 4118 181595 4120
rect 178677 4115 178743 4118
rect 181529 4115 181595 4118
rect 222142 4116 222148 4180
rect 222212 4178 222218 4180
rect 231761 4178 231827 4181
rect 222212 4176 231827 4178
rect 222212 4120 231766 4176
rect 231822 4120 231827 4176
rect 222212 4118 231827 4120
rect 222212 4116 222218 4118
rect 231761 4115 231827 4118
rect 40953 4042 41019 4045
rect 74717 4042 74783 4045
rect 40953 4040 74783 4042
rect 40953 3984 40958 4040
rect 41014 3984 74722 4040
rect 74778 3984 74783 4040
rect 40953 3982 74783 3984
rect 40953 3979 41019 3982
rect 74717 3979 74783 3982
rect 140681 4042 140747 4045
rect 211061 4042 211127 4045
rect 140681 4040 211127 4042
rect 140681 3984 140686 4040
rect 140742 3984 211066 4040
rect 211122 3984 211127 4040
rect 140681 3982 211127 3984
rect 140681 3979 140747 3982
rect 211061 3979 211127 3982
rect 230381 4042 230447 4045
rect 450169 4042 450235 4045
rect 230381 4040 450235 4042
rect 230381 3984 230386 4040
rect 230442 3984 450174 4040
rect 450230 3984 450235 4040
rect 230381 3982 450235 3984
rect 230381 3979 230447 3982
rect 450169 3979 450235 3982
rect 39757 3906 39823 3909
rect 74625 3906 74691 3909
rect 39757 3904 74691 3906
rect 39757 3848 39762 3904
rect 39818 3848 74630 3904
rect 74686 3848 74691 3904
rect 39757 3846 74691 3848
rect 39757 3843 39823 3846
rect 74625 3843 74691 3846
rect 142061 3906 142127 3909
rect 214649 3906 214715 3909
rect 142061 3904 214715 3906
rect 142061 3848 142066 3904
rect 142122 3848 214654 3904
rect 214710 3848 214715 3904
rect 142061 3846 214715 3848
rect 142061 3843 142127 3846
rect 214649 3843 214715 3846
rect 233141 3906 233207 3909
rect 457253 3906 457319 3909
rect 233141 3904 457319 3906
rect 233141 3848 233146 3904
rect 233202 3848 457258 3904
rect 457314 3848 457319 3904
rect 233141 3846 457319 3848
rect 233141 3843 233207 3846
rect 457253 3843 457319 3846
rect 34973 3770 35039 3773
rect 73245 3770 73311 3773
rect 34973 3768 73311 3770
rect 34973 3712 34978 3768
rect 35034 3712 73250 3768
rect 73306 3712 73311 3768
rect 34973 3710 73311 3712
rect 34973 3707 35039 3710
rect 73245 3707 73311 3710
rect 143441 3770 143507 3773
rect 218145 3770 218211 3773
rect 143441 3768 218211 3770
rect 143441 3712 143446 3768
rect 143502 3712 218150 3768
rect 218206 3712 218211 3768
rect 143441 3710 218211 3712
rect 143441 3707 143507 3710
rect 218145 3707 218211 3710
rect 235901 3770 235967 3773
rect 464429 3770 464495 3773
rect 235901 3768 464495 3770
rect 235901 3712 235906 3768
rect 235962 3712 464434 3768
rect 464490 3712 464495 3768
rect 235901 3710 464495 3712
rect 235901 3707 235967 3710
rect 464429 3707 464495 3710
rect 24301 3634 24367 3637
rect 69289 3634 69355 3637
rect 24301 3632 69355 3634
rect 24301 3576 24306 3632
rect 24362 3576 69294 3632
rect 69350 3576 69355 3632
rect 24301 3574 69355 3576
rect 24301 3571 24367 3574
rect 69289 3571 69355 3574
rect 121361 3634 121427 3637
rect 162301 3634 162367 3637
rect 238385 3634 238451 3637
rect 121361 3632 162367 3634
rect 121361 3576 121366 3632
rect 121422 3576 162306 3632
rect 162362 3576 162367 3632
rect 121361 3574 162367 3576
rect 121361 3571 121427 3574
rect 162301 3571 162367 3574
rect 162534 3632 238451 3634
rect 162534 3576 238390 3632
rect 238446 3576 238451 3632
rect 162534 3574 238451 3576
rect 4061 3498 4127 3501
rect 60733 3498 60799 3501
rect 4061 3496 60799 3498
rect 4061 3440 4066 3496
rect 4122 3440 60738 3496
rect 60794 3440 60799 3496
rect 4061 3438 60799 3440
rect 4061 3435 4127 3438
rect 60733 3435 60799 3438
rect 119981 3498 120047 3501
rect 158713 3498 158779 3501
rect 119981 3496 158779 3498
rect 119981 3440 119986 3496
rect 120042 3440 158718 3496
rect 158774 3440 158779 3496
rect 119981 3438 158779 3440
rect 119981 3435 120047 3438
rect 158713 3435 158779 3438
rect 162117 3498 162183 3501
rect 162534 3498 162594 3574
rect 238385 3571 238451 3574
rect 238661 3634 238727 3637
rect 471513 3634 471579 3637
rect 238661 3632 471579 3634
rect 238661 3576 238666 3632
rect 238722 3576 471518 3632
rect 471574 3576 471579 3632
rect 238661 3574 471579 3576
rect 238661 3571 238727 3574
rect 471513 3571 471579 3574
rect 162117 3496 162594 3498
rect 162117 3440 162122 3496
rect 162178 3440 162594 3496
rect 162117 3438 162594 3440
rect 162761 3498 162827 3501
rect 234797 3498 234863 3501
rect 162761 3496 234863 3498
rect 162761 3440 162766 3496
rect 162822 3440 234802 3496
rect 234858 3440 234863 3496
rect 162761 3438 234863 3440
rect 162117 3435 162183 3438
rect 162761 3435 162827 3438
rect 234797 3435 234863 3438
rect 241421 3498 241487 3501
rect 478689 3498 478755 3501
rect 241421 3496 478755 3498
rect 241421 3440 241426 3496
rect 241482 3440 478694 3496
rect 478750 3440 478755 3496
rect 241421 3438 478755 3440
rect 241421 3435 241487 3438
rect 478689 3435 478755 3438
rect 2865 3362 2931 3365
rect 60825 3362 60891 3365
rect 2865 3360 60891 3362
rect 2865 3304 2870 3360
rect 2926 3304 60830 3360
rect 60886 3304 60891 3360
rect 2865 3302 60891 3304
rect 2865 3299 2931 3302
rect 60825 3299 60891 3302
rect 114461 3362 114527 3365
rect 144453 3362 144519 3365
rect 114461 3360 144519 3362
rect 114461 3304 114466 3360
rect 114522 3304 144458 3360
rect 144514 3304 144519 3360
rect 114461 3302 144519 3304
rect 114461 3299 114527 3302
rect 144453 3299 144519 3302
rect 144821 3362 144887 3365
rect 221733 3362 221799 3365
rect 144821 3360 221799 3362
rect 144821 3304 144826 3360
rect 144882 3304 221738 3360
rect 221794 3304 221799 3360
rect 144821 3302 221799 3304
rect 144821 3299 144887 3302
rect 221733 3299 221799 3302
rect 311198 3300 311204 3364
rect 311268 3362 311274 3364
rect 314561 3362 314627 3365
rect 311268 3360 314627 3362
rect 311268 3304 314566 3360
rect 314622 3304 314627 3360
rect 311268 3302 314627 3304
rect 311268 3300 311274 3302
rect 314561 3299 314627 3302
rect 321502 3300 321508 3364
rect 321572 3362 321578 3364
rect 321645 3362 321711 3365
rect 321572 3360 321711 3362
rect 321572 3304 321650 3360
rect 321706 3304 321711 3360
rect 321572 3302 321711 3304
rect 321572 3300 321578 3302
rect 321645 3299 321711 3302
rect 321829 3362 321895 3365
rect 582189 3362 582255 3365
rect 321829 3360 582255 3362
rect 321829 3304 321834 3360
rect 321890 3304 582194 3360
rect 582250 3304 582255 3360
rect 321829 3302 582255 3304
rect 321829 3299 321895 3302
rect 582189 3299 582255 3302
rect 124029 3226 124095 3229
rect 169385 3226 169451 3229
rect 124029 3224 169451 3226
rect 124029 3168 124034 3224
rect 124090 3168 169390 3224
rect 169446 3168 169451 3224
rect 124029 3166 169451 3168
rect 124029 3163 124095 3166
rect 169385 3163 169451 3166
rect 186129 3226 186195 3229
rect 186405 3226 186471 3229
rect 186129 3224 186471 3226
rect 186129 3168 186134 3224
rect 186190 3168 186410 3224
rect 186466 3168 186471 3224
rect 186129 3166 186471 3168
rect 186129 3163 186195 3166
rect 186405 3163 186471 3166
rect 296069 3226 296135 3229
rect 435817 3226 435883 3229
rect 296069 3224 435883 3226
rect 296069 3168 296074 3224
rect 296130 3168 435822 3224
rect 435878 3168 435883 3224
rect 296069 3166 435883 3168
rect 296069 3163 296135 3166
rect 435817 3163 435883 3166
rect 118601 3090 118667 3093
rect 153929 3090 153995 3093
rect 118601 3088 153995 3090
rect 118601 3032 118606 3088
rect 118662 3032 153934 3088
rect 153990 3032 153995 3088
rect 118601 3030 153995 3032
rect 118601 3027 118667 3030
rect 153929 3027 153995 3030
rect 159357 3090 159423 3093
rect 162761 3090 162827 3093
rect 159357 3088 162827 3090
rect 159357 3032 159362 3088
rect 159418 3032 162766 3088
rect 162822 3032 162827 3088
rect 159357 3030 162827 3032
rect 159357 3027 159423 3030
rect 162761 3027 162827 3030
rect 171777 3090 171843 3093
rect 176745 3090 176811 3093
rect 171777 3088 176811 3090
rect 171777 3032 171782 3088
rect 171838 3032 176750 3088
rect 176806 3032 176811 3088
rect 171777 3030 176811 3032
rect 171777 3027 171843 3030
rect 176745 3027 176811 3030
rect 320766 3028 320772 3092
rect 320836 3090 320842 3092
rect 321829 3090 321895 3093
rect 320836 3088 321895 3090
rect 320836 3032 321834 3088
rect 321890 3032 321895 3088
rect 320836 3030 321895 3032
rect 320836 3028 320842 3030
rect 321829 3027 321895 3030
rect 115749 2954 115815 2957
rect 146845 2954 146911 2957
rect 115749 2952 146911 2954
rect 115749 2896 115754 2952
rect 115810 2896 146850 2952
rect 146906 2896 146911 2952
rect 115749 2894 146911 2896
rect 115749 2891 115815 2894
rect 146845 2891 146911 2894
rect 129549 2818 129615 2821
rect 133965 2818 134031 2821
rect 129549 2816 134031 2818
rect 129549 2760 129554 2816
rect 129610 2760 133970 2816
rect 134026 2760 134031 2816
rect 129549 2758 134031 2760
rect 129549 2755 129615 2758
rect 133965 2755 134031 2758
<< via3 >>
rect 129228 652896 129292 652900
rect 129228 652840 129278 652896
rect 129278 652840 129292 652896
rect 129228 652836 129292 652840
rect 133644 652896 133708 652900
rect 133644 652840 133694 652896
rect 133694 652840 133708 652896
rect 133644 652836 133708 652840
rect 259132 652896 259196 652900
rect 259132 652840 259182 652896
rect 259182 652840 259196 652896
rect 259132 652836 259196 652840
rect 263548 652896 263612 652900
rect 263548 652840 263598 652896
rect 263598 652840 263612 652896
rect 263548 652836 263612 652840
rect 378180 652896 378244 652900
rect 378180 652840 378194 652896
rect 378194 652840 378244 652896
rect 378180 652836 378244 652840
rect 383516 652896 383580 652900
rect 383516 652840 383566 652896
rect 383566 652840 383580 652896
rect 383516 652836 383580 652840
rect 508452 652896 508516 652900
rect 508452 652840 508466 652896
rect 508466 652840 508516 652896
rect 508452 652836 508516 652840
rect 513420 652896 513484 652900
rect 513420 652840 513434 652896
rect 513434 652840 513484 652896
rect 513420 652836 513484 652840
rect 282316 648680 282380 648684
rect 282316 648624 282330 648680
rect 282330 648624 282380 648680
rect 282316 648620 282380 648624
rect 282684 587148 282748 587212
rect 269068 580892 269132 580956
rect 387564 587148 387628 587212
rect 518940 580892 519004 580956
rect 137508 580348 137572 580412
rect 440004 579124 440068 579188
rect 60596 578988 60660 579052
rect 190132 578988 190196 579052
rect 229324 560008 229388 560012
rect 229324 559952 229374 560008
rect 229374 559952 229388 560008
rect 229324 559948 229388 559952
rect 225828 559812 225892 559876
rect 227116 559268 227180 559332
rect 351868 559268 351932 559332
rect 358860 559268 358924 559332
rect 67404 558860 67468 558924
rect 68508 558860 68572 558924
rect 70164 558920 70228 558924
rect 70164 558864 70214 558920
rect 70214 558864 70228 558920
rect 70164 558860 70228 558864
rect 71636 558920 71700 558924
rect 71636 558864 71686 558920
rect 71686 558864 71700 558920
rect 71636 558860 71700 558864
rect 72372 558860 72436 558924
rect 72924 558860 72988 558924
rect 73660 558920 73724 558924
rect 73660 558864 73710 558920
rect 73710 558864 73724 558920
rect 73660 558860 73724 558864
rect 74212 558920 74276 558924
rect 74212 558864 74262 558920
rect 74262 558864 74276 558920
rect 74212 558860 74276 558864
rect 74948 558920 75012 558924
rect 74948 558864 74998 558920
rect 74998 558864 75012 558920
rect 74948 558860 75012 558864
rect 75684 558860 75748 558924
rect 76788 558920 76852 558924
rect 76788 558864 76838 558920
rect 76838 558864 76852 558920
rect 76788 558860 76852 558864
rect 77340 558920 77404 558924
rect 77340 558864 77390 558920
rect 77390 558864 77404 558920
rect 77340 558860 77404 558864
rect 78076 558860 78140 558924
rect 79180 558860 79244 558924
rect 79916 558920 79980 558924
rect 79916 558864 79966 558920
rect 79966 558864 79980 558920
rect 79916 558860 79980 558864
rect 80652 558860 80716 558924
rect 81204 558920 81268 558924
rect 81204 558864 81254 558920
rect 81254 558864 81268 558920
rect 81204 558860 81268 558864
rect 81940 558920 82004 558924
rect 81940 558864 81990 558920
rect 81990 558864 82004 558920
rect 81940 558860 82004 558864
rect 82676 558920 82740 558924
rect 82676 558864 82726 558920
rect 82726 558864 82740 558920
rect 82676 558860 82740 558864
rect 83780 558920 83844 558924
rect 83780 558864 83830 558920
rect 83830 558864 83844 558920
rect 83780 558860 83844 558864
rect 84148 558920 84212 558924
rect 84148 558864 84198 558920
rect 84198 558864 84212 558920
rect 84148 558860 84212 558864
rect 85068 558860 85132 558924
rect 86724 558920 86788 558924
rect 86724 558864 86774 558920
rect 86774 558864 86788 558920
rect 86724 558860 86788 558864
rect 87828 558920 87892 558924
rect 87828 558864 87878 558920
rect 87878 558864 87892 558920
rect 87828 558860 87892 558864
rect 88196 558920 88260 558924
rect 88196 558864 88246 558920
rect 88246 558864 88260 558920
rect 88196 558860 88260 558864
rect 88932 558920 88996 558924
rect 88932 558864 88946 558920
rect 88946 558864 88996 558920
rect 88932 558860 88996 558864
rect 89116 558860 89180 558924
rect 89852 558920 89916 558924
rect 89852 558864 89866 558920
rect 89866 558864 89916 558920
rect 89852 558860 89916 558864
rect 90956 558920 91020 558924
rect 90956 558864 91006 558920
rect 91006 558864 91020 558920
rect 90956 558860 91020 558864
rect 92060 558860 92124 558924
rect 92428 558920 92492 558924
rect 92428 558864 92478 558920
rect 92478 558864 92492 558920
rect 92428 558860 92492 558864
rect 93164 558860 93228 558924
rect 94820 558920 94884 558924
rect 94820 558864 94870 558920
rect 94870 558864 94884 558920
rect 94820 558860 94884 558864
rect 95004 558920 95068 558924
rect 95004 558864 95054 558920
rect 95054 558864 95068 558920
rect 95004 558860 95068 558864
rect 95740 558920 95804 558924
rect 95740 558864 95754 558920
rect 95754 558864 95804 558920
rect 95740 558860 95804 558864
rect 96476 558920 96540 558924
rect 96476 558864 96526 558920
rect 96526 558864 96540 558920
rect 96476 558860 96540 558864
rect 97028 558920 97092 558924
rect 97028 558864 97078 558920
rect 97078 558864 97092 558920
rect 97028 558860 97092 558864
rect 97580 558920 97644 558924
rect 97580 558864 97630 558920
rect 97630 558864 97644 558920
rect 97580 558860 97644 558864
rect 98316 558860 98380 558924
rect 99052 558860 99116 558924
rect 100156 558860 100220 558924
rect 101996 558920 102060 558924
rect 101996 558864 102046 558920
rect 102046 558864 102060 558920
rect 101996 558860 102060 558864
rect 104756 558920 104820 558924
rect 104756 558864 104806 558920
rect 104806 558864 104820 558920
rect 104756 558860 104820 558864
rect 107148 558860 107212 558924
rect 108436 558920 108500 558924
rect 108436 558864 108486 558920
rect 108486 558864 108500 558920
rect 108436 558860 108500 558864
rect 194364 558920 194428 558924
rect 194364 558864 194414 558920
rect 194414 558864 194428 558920
rect 194364 558860 194428 558864
rect 196204 558860 196268 558924
rect 200252 558920 200316 558924
rect 200252 558864 200266 558920
rect 200266 558864 200316 558920
rect 200252 558860 200316 558864
rect 201540 558920 201604 558924
rect 201540 558864 201554 558920
rect 201554 558864 201604 558920
rect 201540 558860 201604 558864
rect 202644 558860 202708 558924
rect 203748 558920 203812 558924
rect 203748 558864 203798 558920
rect 203798 558864 203812 558920
rect 203748 558860 203812 558864
rect 203932 558860 203996 558924
rect 205404 558860 205468 558924
rect 206140 558860 206204 558924
rect 208348 558860 208412 558924
rect 211844 558920 211908 558924
rect 211844 558864 211894 558920
rect 211894 558864 211908 558920
rect 211844 558860 211908 558864
rect 213132 558920 213196 558924
rect 213132 558864 213146 558920
rect 213146 558864 213196 558920
rect 213132 558860 213196 558864
rect 214052 558860 214116 558924
rect 215340 558920 215404 558924
rect 215340 558864 215354 558920
rect 215354 558864 215404 558920
rect 215340 558860 215404 558864
rect 218836 558920 218900 558924
rect 218836 558864 218850 558920
rect 218850 558864 218900 558920
rect 218836 558860 218900 558864
rect 220124 558920 220188 558924
rect 220124 558864 220138 558920
rect 220138 558864 220188 558920
rect 220124 558860 220188 558864
rect 221044 558920 221108 558924
rect 221044 558864 221094 558920
rect 221094 558864 221108 558920
rect 221044 558860 221108 558864
rect 222332 558920 222396 558924
rect 222332 558864 222346 558920
rect 222346 558864 222396 558920
rect 222332 558860 222396 558864
rect 223620 558920 223684 558924
rect 223620 558864 223634 558920
rect 223634 558864 223684 558920
rect 223620 558860 223684 558864
rect 224540 558860 224604 558924
rect 228036 558920 228100 558924
rect 228036 558864 228086 558920
rect 228086 558864 228100 558920
rect 228036 558860 228100 558864
rect 235764 558860 235828 558924
rect 237236 558920 237300 558924
rect 237236 558864 237286 558920
rect 237286 558864 237300 558920
rect 237236 558860 237300 558864
rect 239628 558860 239692 558924
rect 313780 558920 313844 558924
rect 313780 558864 313794 558920
rect 313794 558864 313844 558920
rect 313780 558860 313844 558864
rect 316172 558860 316236 558924
rect 317460 558920 317524 558924
rect 317460 558864 317474 558920
rect 317474 558864 317524 558920
rect 317460 558860 317524 558864
rect 320956 558860 321020 558924
rect 322612 558860 322676 558924
rect 323532 558920 323596 558924
rect 323532 558864 323546 558920
rect 323546 558864 323596 558920
rect 323532 558860 323596 558864
rect 328500 558920 328564 558924
rect 328500 558864 328550 558920
rect 328550 558864 328564 558920
rect 328500 558860 328564 558864
rect 329604 558920 329668 558924
rect 329604 558864 329618 558920
rect 329618 558864 329668 558920
rect 329604 558860 329668 558864
rect 330524 558920 330588 558924
rect 330524 558864 330538 558920
rect 330538 558864 330588 558920
rect 330524 558860 330588 558864
rect 331812 558860 331876 558924
rect 333100 558920 333164 558924
rect 333100 558864 333150 558920
rect 333150 558864 333164 558920
rect 333100 558860 333164 558864
rect 334020 558860 334084 558924
rect 335492 558860 335556 558924
rect 336412 558860 336476 558924
rect 337700 558920 337764 558924
rect 337700 558864 337750 558920
rect 337750 558864 337764 558920
rect 337700 558860 337764 558864
rect 338988 558920 339052 558924
rect 338988 558864 339038 558920
rect 339038 558864 339052 558920
rect 338988 558860 339052 558864
rect 339908 558920 339972 558924
rect 339908 558864 339922 558920
rect 339922 558864 339972 558920
rect 339908 558860 339972 558864
rect 341196 558920 341260 558924
rect 341196 558864 341246 558920
rect 341246 558864 341260 558920
rect 341196 558860 341260 558864
rect 342484 558920 342548 558924
rect 342484 558864 342534 558920
rect 342534 558864 342548 558920
rect 342484 558860 342548 558864
rect 343588 558920 343652 558924
rect 343588 558864 343638 558920
rect 343638 558864 343652 558920
rect 343588 558860 343652 558864
rect 344692 558860 344756 558924
rect 345796 558920 345860 558924
rect 345796 558864 345810 558920
rect 345810 558864 345860 558920
rect 345796 558860 345860 558864
rect 346532 558920 346596 558924
rect 346532 558864 346546 558920
rect 346546 558864 346596 558920
rect 346532 558860 346596 558864
rect 348188 558920 348252 558924
rect 348188 558864 348238 558920
rect 348238 558864 348252 558920
rect 348188 558860 348252 558864
rect 349476 558860 349540 558924
rect 350580 558920 350644 558924
rect 350580 558864 350594 558920
rect 350594 558864 350644 558920
rect 350580 558860 350644 558864
rect 352420 558860 352484 558924
rect 353524 558860 353588 558924
rect 443132 558920 443196 558924
rect 443132 558864 443146 558920
rect 443146 558864 443196 558920
rect 443132 558860 443196 558864
rect 446260 558860 446324 558924
rect 447732 558860 447796 558924
rect 453620 558920 453684 558924
rect 453620 558864 453670 558920
rect 453670 558864 453684 558920
rect 453620 558860 453684 558864
rect 454724 558920 454788 558924
rect 454724 558864 454738 558920
rect 454738 558864 454788 558920
rect 454724 558860 454788 558864
rect 456012 558920 456076 558924
rect 456012 558864 456026 558920
rect 456026 558864 456076 558920
rect 456012 558860 456076 558864
rect 457300 558920 457364 558924
rect 457300 558864 457350 558920
rect 457350 558864 457364 558920
rect 457300 558860 457364 558864
rect 458220 558920 458284 558924
rect 458220 558864 458270 558920
rect 458270 558864 458284 558920
rect 458220 558860 458284 558864
rect 460796 558920 460860 558924
rect 460796 558864 460846 558920
rect 460846 558864 460860 558920
rect 460796 558860 460860 558864
rect 461716 558920 461780 558924
rect 461716 558864 461730 558920
rect 461730 558864 461780 558920
rect 461716 558860 461780 558864
rect 462636 558920 462700 558924
rect 462636 558864 462650 558920
rect 462650 558864 462700 558920
rect 462636 558860 462700 558864
rect 464292 558920 464356 558924
rect 464292 558864 464306 558920
rect 464306 558864 464356 558920
rect 464292 558860 464356 558864
rect 465212 558920 465276 558924
rect 465212 558864 465262 558920
rect 465262 558864 465276 558920
rect 465212 558860 465276 558864
rect 466868 558860 466932 558924
rect 467972 558860 468036 558924
rect 468708 558920 468772 558924
rect 468708 558864 468722 558920
rect 468722 558864 468772 558920
rect 468708 558860 468772 558864
rect 470364 558860 470428 558924
rect 471468 558860 471532 558924
rect 472756 558860 472820 558924
rect 474044 558860 474108 558924
rect 474780 558920 474844 558924
rect 474780 558864 474830 558920
rect 474830 558864 474844 558920
rect 474780 558860 474844 558864
rect 475516 558920 475580 558924
rect 475516 558864 475530 558920
rect 475530 558864 475580 558920
rect 475516 558860 475580 558864
rect 477172 558920 477236 558924
rect 477172 558864 477186 558920
rect 477186 558864 477236 558920
rect 477172 558860 477236 558864
rect 478276 558920 478340 558924
rect 478276 558864 478290 558920
rect 478290 558864 478340 558920
rect 478276 558860 478340 558864
rect 479012 558920 479076 558924
rect 479012 558864 479026 558920
rect 479026 558864 479076 558920
rect 479012 558860 479076 558864
rect 480852 558860 480916 558924
rect 483612 558860 483676 558924
rect 69796 558724 69860 558788
rect 75868 558784 75932 558788
rect 75868 558728 75918 558784
rect 75918 558728 75932 558784
rect 75868 558724 75932 558728
rect 78444 558784 78508 558788
rect 78444 558728 78494 558784
rect 78494 558728 78508 558784
rect 78444 558724 78508 558728
rect 79364 558724 79428 558788
rect 82860 558784 82924 558788
rect 82860 558728 82910 558784
rect 82910 558728 82924 558784
rect 82860 558724 82924 558728
rect 85436 558784 85500 558788
rect 85436 558728 85450 558784
rect 85450 558728 85500 558784
rect 85436 558724 85500 558728
rect 86172 558724 86236 558788
rect 91140 558784 91204 558788
rect 91140 558728 91154 558784
rect 91154 558728 91204 558784
rect 91140 558724 91204 558728
rect 93716 558784 93780 558788
rect 93716 558728 93766 558784
rect 93766 558728 93780 558784
rect 93716 558724 93780 558728
rect 105308 558724 105372 558788
rect 202460 558724 202524 558788
rect 216628 558724 216692 558788
rect 232820 558724 232884 558788
rect 233556 558724 233620 558788
rect 234660 558784 234724 558788
rect 234660 558728 234674 558784
rect 234674 558728 234724 558784
rect 234660 558724 234724 558728
rect 236132 558724 236196 558788
rect 320220 558784 320284 558788
rect 320220 558728 320234 558784
rect 320234 558728 320284 558784
rect 320220 558724 320284 558728
rect 354812 558724 354876 558788
rect 356100 558784 356164 558788
rect 356100 558728 356114 558784
rect 356114 558728 356164 558784
rect 356100 558724 356164 558728
rect 453804 558724 453868 558788
rect 466500 558784 466564 558788
rect 466500 558728 466550 558784
rect 466550 558728 466564 558784
rect 466500 558724 466564 558728
rect 469076 558724 469140 558788
rect 469996 558784 470060 558788
rect 469996 558728 470046 558784
rect 470046 558728 470060 558784
rect 469996 558724 470060 558728
rect 471284 558784 471348 558788
rect 471284 558728 471334 558784
rect 471334 558728 471348 558784
rect 471284 558724 471348 558728
rect 472204 558784 472268 558788
rect 472204 558728 472218 558784
rect 472218 558728 472268 558784
rect 472204 558724 472268 558728
rect 480484 558724 480548 558788
rect 481588 558784 481652 558788
rect 481588 558728 481638 558784
rect 481638 558728 481652 558784
rect 481588 558724 481652 558728
rect 86356 558588 86420 558652
rect 93532 558648 93596 558652
rect 93532 558592 93582 558648
rect 93582 558592 93596 558648
rect 93532 558588 93596 558592
rect 204852 558648 204916 558652
rect 204852 558592 204902 558648
rect 204902 558592 204916 558648
rect 204852 558588 204916 558592
rect 210556 558648 210620 558652
rect 210556 558592 210570 558648
rect 210570 558592 210620 558648
rect 210556 558588 210620 558592
rect 217548 558588 217612 558652
rect 231900 558648 231964 558652
rect 231900 558592 231914 558648
rect 231914 558592 231964 558648
rect 231900 558588 231964 558592
rect 237420 558648 237484 558652
rect 237420 558592 237434 558648
rect 237434 558592 237484 558648
rect 237420 558588 237484 558592
rect 318932 558588 318996 558652
rect 452700 558588 452764 558652
rect 459508 558588 459572 558652
rect 467788 558588 467852 558652
rect 473492 558648 473556 558652
rect 473492 558592 473506 558648
rect 473506 558592 473556 558648
rect 473492 558588 473556 558592
rect 484716 558588 484780 558652
rect 488580 558648 488644 558652
rect 488580 558592 488594 558648
rect 488594 558592 488644 558648
rect 488580 558588 488644 558592
rect 99420 558512 99484 558516
rect 99420 558456 99434 558512
rect 99434 558456 99484 558512
rect 99420 558452 99484 558456
rect 108620 558452 108684 558516
rect 230612 558452 230676 558516
rect 357572 558452 357636 558516
rect 449940 558512 450004 558516
rect 449940 558456 449954 558512
rect 449954 558456 450004 558512
rect 449940 558452 450004 558456
rect 477356 558452 477420 558516
rect 482140 558452 482204 558516
rect 486004 558452 486068 558516
rect 487292 558452 487356 558516
rect 197308 558316 197372 558380
rect 238708 558376 238772 558380
rect 238708 558320 238758 558376
rect 238758 558320 238772 558376
rect 238708 558316 238772 558320
rect 474964 558316 475028 558380
rect 476252 558376 476316 558380
rect 476252 558320 476266 558376
rect 476266 558320 476316 558376
rect 476252 558316 476316 558320
rect 478460 558316 478524 558380
rect 198780 558180 198844 558244
rect 448468 558180 448532 558244
rect 479748 558180 479812 558244
rect 483428 558180 483492 558244
rect 485636 558180 485700 558244
rect 486924 558180 486988 558244
rect 64276 558044 64340 558108
rect 238340 558044 238404 558108
rect 451412 558044 451476 558108
rect 484164 558044 484228 558108
rect 489132 558044 489196 558108
rect 487844 557908 487908 557972
rect 100340 557772 100404 557836
rect 101628 557636 101692 557700
rect 106228 557696 106292 557700
rect 106228 557640 106278 557696
rect 106278 557640 106292 557696
rect 106228 557636 106292 557640
rect 207060 557636 207124 557700
rect 209636 557636 209700 557700
rect 210372 557636 210436 557700
rect 217364 557636 217428 557700
rect 225644 557636 225708 557700
rect 232636 557636 232700 557700
rect 324820 557636 324884 557700
rect 326108 557636 326172 557700
rect 327028 557636 327092 557700
rect 331076 557636 331140 557700
rect 337884 557636 337948 557700
rect 344876 557636 344940 557700
rect 353156 557636 353220 557700
rect 462084 557636 462148 557700
rect 483060 557696 483124 557700
rect 483060 557640 483074 557696
rect 483074 557640 483124 557696
rect 483060 557636 483124 557640
rect 101444 557500 101508 557564
rect 102732 557560 102796 557564
rect 102732 557504 102782 557560
rect 102782 557504 102796 557560
rect 102732 557500 102796 557504
rect 103284 557500 103348 557564
rect 104020 557500 104084 557564
rect 105308 557500 105372 557564
rect 106044 557500 106108 557564
rect 107700 557560 107764 557564
rect 107700 557504 107714 557560
rect 107714 557504 107764 557560
rect 107700 557500 107764 557504
rect 108988 557500 109052 557564
rect 206876 557560 206940 557564
rect 206876 557504 206926 557560
rect 206926 557504 206940 557560
rect 206876 557500 206940 557504
rect 207980 557500 208044 557564
rect 209268 557500 209332 557564
rect 210924 557500 210988 557564
rect 212396 557560 212460 557564
rect 212396 557504 212446 557560
rect 212446 557504 212460 557560
rect 212396 557500 212460 557504
rect 213500 557500 213564 557564
rect 214788 557500 214852 557564
rect 216260 557500 216324 557564
rect 217916 557560 217980 557564
rect 217916 557504 217966 557560
rect 217966 557504 217980 557560
rect 217916 557500 217980 557504
rect 219204 557500 219268 557564
rect 220676 557560 220740 557564
rect 220676 557504 220726 557560
rect 220726 557504 220740 557560
rect 220676 557500 220740 557504
rect 221964 557500 222028 557564
rect 223252 557500 223316 557564
rect 224356 557500 224420 557564
rect 226196 557560 226260 557564
rect 226196 557504 226210 557560
rect 226210 557504 226260 557560
rect 226196 557500 226260 557504
rect 227484 557500 227548 557564
rect 228772 557500 228836 557564
rect 230244 557500 230308 557564
rect 230796 557500 230860 557564
rect 233004 557560 233068 557564
rect 233004 557504 233054 557560
rect 233054 557504 233068 557560
rect 233004 557500 233068 557504
rect 234476 557560 234540 557564
rect 234476 557504 234526 557560
rect 234526 557504 234540 557560
rect 234476 557500 234540 557504
rect 322796 557500 322860 557564
rect 324084 557500 324148 557564
rect 325372 557500 325436 557564
rect 326292 557500 326356 557564
rect 327580 557500 327644 557564
rect 328868 557500 328932 557564
rect 329788 557560 329852 557564
rect 329788 557504 329838 557560
rect 329838 557504 329852 557560
rect 329788 557500 329852 557504
rect 332364 557500 332428 557564
rect 333284 557500 333348 557564
rect 334572 557500 334636 557564
rect 335860 557500 335924 557564
rect 336780 557560 336844 557564
rect 336780 557504 336794 557560
rect 336794 557504 336844 557560
rect 336780 557500 336844 557504
rect 339172 557500 339236 557564
rect 340460 557500 340524 557564
rect 341748 557500 341812 557564
rect 342668 557500 342732 557564
rect 343956 557500 344020 557564
rect 346164 557500 346228 557564
rect 347452 557500 347516 557564
rect 348740 557500 348804 557564
rect 349660 557500 349724 557564
rect 350948 557500 351012 557564
rect 354444 557500 354508 557564
rect 355732 557500 355796 557564
rect 356652 557500 356716 557564
rect 357940 557500 358004 557564
rect 452884 557500 452948 557564
rect 455276 557500 455340 557564
rect 456564 557500 456628 557564
rect 457484 557500 457548 557564
rect 458772 557500 458836 557564
rect 460060 557500 460124 557564
rect 460980 557560 461044 557564
rect 460980 557504 460994 557560
rect 460994 557504 461044 557560
rect 460980 557500 461044 557504
rect 463556 557500 463620 557564
rect 464476 557500 464540 557564
rect 465764 557500 465828 557564
rect 352236 555520 352300 555524
rect 352236 555464 352250 555520
rect 352250 555464 352300 555520
rect 352236 555460 352300 555464
rect 359228 555460 359292 555524
rect 383516 413264 383580 413268
rect 383516 413208 383566 413264
rect 383566 413208 383580 413264
rect 383516 413204 383580 413208
rect 513420 412720 513484 412724
rect 513420 412664 513434 412720
rect 513434 412664 513484 412720
rect 513420 412660 513484 412664
rect 282316 322900 282380 322964
rect 313412 318684 313476 318748
rect 443132 318744 443196 318748
rect 443132 318688 443146 318744
rect 443146 318688 443196 318744
rect 443132 318684 443196 318688
rect 144868 318412 144932 318476
rect 320772 318276 320836 318340
rect 144868 318140 144932 318204
rect 311204 318140 311268 318204
rect 321508 318004 321572 318068
rect 135116 280060 135180 280124
rect 81756 278760 81820 278764
rect 81756 278704 81770 278760
rect 81770 278704 81820 278760
rect 81756 278700 81820 278704
rect 135116 270540 135180 270604
rect 81756 270404 81820 270468
rect 135116 260748 135180 260812
rect 135116 251228 135180 251292
rect 135116 61432 135180 61436
rect 135116 61376 135130 61432
rect 135130 61376 135180 61432
rect 135116 61372 135180 61376
rect 135116 48316 135180 48380
rect 124444 42120 124508 42124
rect 124444 42064 124494 42120
rect 124494 42064 124508 42120
rect 124444 42060 124508 42064
rect 135116 42120 135180 42124
rect 135116 42064 135130 42120
rect 135130 42064 135180 42120
rect 135116 42060 135180 42064
rect 124444 32464 124508 32468
rect 124444 32408 124458 32464
rect 124458 32408 124508 32464
rect 124444 32404 124508 32408
rect 135116 29004 135180 29068
rect 222148 4388 222212 4452
rect 249748 4524 249812 4588
rect 269068 4524 269132 4588
rect 249748 4252 249812 4316
rect 269068 4252 269132 4316
rect 222148 4116 222212 4180
rect 311204 3300 311268 3364
rect 321508 3300 321572 3364
rect 320772 3028 320836 3092
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 654247 59004 671498
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 654247 62604 675098
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 654247 66204 678698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 654247 73404 685898
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654247 77004 689498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 654247 80604 657098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 654247 84204 660698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 654247 91404 667898
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 654247 95004 671498
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 654247 98604 675098
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 654247 102204 678698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 654247 109404 685898
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654247 113004 689498
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 654247 116604 657098
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 654247 120204 660698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 654247 127404 667898
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 654247 131004 671498
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 654247 134604 675098
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 654247 138204 678698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 129227 652900 129293 652901
rect 129227 652836 129228 652900
rect 129292 652836 129293 652900
rect 129227 652835 129293 652836
rect 133643 652900 133709 652901
rect 133643 652836 133644 652900
rect 133708 652836 133709 652900
rect 133643 652835 133709 652836
rect 129230 651130 129290 652835
rect 133646 651810 133706 652835
rect 128608 651070 129290 651130
rect 133573 651750 133706 651810
rect 133573 651100 133633 651750
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 136938 643254 137262 643276
rect 136938 643018 136982 643254
rect 137218 643018 137262 643254
rect 136938 642934 137262 643018
rect 136938 642698 136982 642934
rect 137218 642698 137262 642934
rect 136938 642676 137262 642698
rect 136938 639654 137262 639676
rect 136938 639418 136982 639654
rect 137218 639418 137262 639654
rect 136938 639334 137262 639418
rect 136938 639098 136982 639334
rect 137218 639098 137262 639334
rect 136938 639076 137262 639098
rect 136938 636054 137262 636076
rect 136938 635818 136982 636054
rect 137218 635818 137262 636054
rect 136938 635734 137262 635818
rect 136938 635498 136982 635734
rect 137218 635498 137262 635734
rect 136938 635476 137262 635498
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 136938 632454 137262 632476
rect 136938 632218 136982 632454
rect 137218 632218 137262 632454
rect 136938 632134 137262 632218
rect 136938 631898 136982 632134
rect 137218 631898 137262 632134
rect 136938 631876 137262 631898
rect 136494 625254 136814 625276
rect 136494 625018 136536 625254
rect 136772 625018 136814 625254
rect 136494 624934 136814 625018
rect 136494 624698 136536 624934
rect 136772 624698 136814 624934
rect 136494 624676 136814 624698
rect 136494 621654 136814 621676
rect 136494 621418 136536 621654
rect 136772 621418 136814 621654
rect 136494 621334 136814 621418
rect 136494 621098 136536 621334
rect 136772 621098 136814 621334
rect 136494 621076 136814 621098
rect 136494 618054 136814 618076
rect 136494 617818 136536 618054
rect 136772 617818 136814 618054
rect 136494 617734 136814 617818
rect 136494 617498 136536 617734
rect 136772 617498 136814 617734
rect 136494 617476 136814 617498
rect 136494 614454 136814 614476
rect 136494 614218 136536 614454
rect 136772 614218 136814 614454
rect 136494 614134 136814 614218
rect 136494 613898 136536 614134
rect 136772 613898 136814 614134
rect 136494 613876 136814 613898
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 136938 607254 137262 607276
rect 136938 607018 136982 607254
rect 137218 607018 137262 607254
rect 136938 606934 137262 607018
rect 136938 606698 136982 606934
rect 137218 606698 137262 606934
rect 136938 606676 137262 606698
rect 136938 603654 137262 603676
rect 136938 603418 136982 603654
rect 137218 603418 137262 603654
rect 136938 603334 137262 603418
rect 136938 603098 136982 603334
rect 137218 603098 137262 603334
rect 136938 603076 137262 603098
rect 136938 600054 137262 600076
rect 136938 599818 136982 600054
rect 137218 599818 137262 600054
rect 136938 599734 137262 599818
rect 136938 599498 136982 599734
rect 137218 599498 137262 599734
rect 136938 599476 137262 599498
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 136938 596454 137262 596476
rect 136938 596218 136982 596454
rect 137218 596218 137262 596454
rect 136938 596134 137262 596218
rect 136938 595898 136982 596134
rect 137218 595898 137262 596134
rect 136938 595876 137262 595898
rect 136494 589254 136814 589276
rect 136494 589018 136536 589254
rect 136772 589018 136814 589254
rect 136494 588934 136814 589018
rect 136494 588698 136536 588934
rect 136772 588698 136814 588934
rect 136494 588676 136814 588698
rect 136494 585654 136814 585676
rect 136494 585418 136536 585654
rect 136772 585418 136814 585654
rect 136494 585334 136814 585418
rect 136494 585098 136536 585334
rect 136772 585098 136814 585334
rect 136494 585076 136814 585098
rect 136494 582054 136814 582076
rect 136494 581818 136536 582054
rect 136772 581818 136814 582054
rect 136494 581734 136814 581818
rect 136494 581498 136536 581734
rect 136772 581498 136814 581734
rect 136494 581476 136814 581498
rect 137507 580412 137573 580413
rect 137507 580348 137508 580412
rect 137572 580348 137573 580412
rect 137507 580347 137573 580348
rect 137510 579138 137570 580347
rect 136494 578454 136814 578476
rect 136494 578218 136536 578454
rect 136772 578218 136814 578454
rect 136494 578134 136814 578218
rect 136494 577898 136536 578134
rect 136772 577898 136814 578134
rect 136494 577876 136814 577898
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 136938 571254 137262 571276
rect 136938 571018 136982 571254
rect 137218 571018 137262 571254
rect 136938 570934 137262 571018
rect 136938 570698 136982 570934
rect 137218 570698 137262 570934
rect 136938 570676 137262 570698
rect 136938 567654 137262 567676
rect 136938 567418 136982 567654
rect 137218 567418 137262 567654
rect 136938 567334 137262 567418
rect 136938 567098 136982 567334
rect 137218 567098 137262 567334
rect 136938 567076 137262 567098
rect 136938 564054 137262 564076
rect 136938 563818 136982 564054
rect 137218 563818 137262 564054
rect 136938 563734 137262 563818
rect 136938 563498 136982 563734
rect 137218 563498 137262 563734
rect 136938 563476 137262 563498
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 72374 560430 72672 560490
rect 79366 560430 79680 560490
rect 82862 560430 83184 560490
rect 86358 560430 86688 560490
rect 102734 560430 103040 560490
rect 106230 560430 106544 560490
rect 63833 560290 64338 560350
rect 66832 560290 67466 560350
rect 68000 560290 68570 560350
rect 69168 560290 69858 560350
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 64278 558109 64338 560290
rect 67406 558925 67466 560290
rect 68510 558925 68570 560290
rect 67403 558924 67469 558925
rect 67403 558860 67404 558924
rect 67468 558860 67469 558924
rect 67403 558859 67469 558860
rect 68507 558924 68573 558925
rect 68507 558860 68508 558924
rect 68572 558860 68573 558924
rect 68507 558859 68573 558860
rect 69798 558789 69858 560290
rect 70166 560290 70336 560350
rect 71504 560290 71698 560350
rect 70166 558925 70226 560290
rect 71638 558925 71698 560290
rect 72374 558925 72434 560430
rect 72796 560290 72986 560350
rect 72926 558925 72986 560290
rect 73662 560290 73840 560350
rect 73964 560290 74274 560350
rect 73662 558925 73722 560290
rect 74214 558925 74274 560290
rect 74950 558925 75010 560350
rect 75132 560290 75746 560350
rect 75686 558925 75746 560290
rect 75870 560290 76176 560350
rect 76300 560290 76850 560350
rect 70163 558924 70229 558925
rect 70163 558860 70164 558924
rect 70228 558860 70229 558924
rect 70163 558859 70229 558860
rect 71635 558924 71701 558925
rect 71635 558860 71636 558924
rect 71700 558860 71701 558924
rect 71635 558859 71701 558860
rect 72371 558924 72437 558925
rect 72371 558860 72372 558924
rect 72436 558860 72437 558924
rect 72371 558859 72437 558860
rect 72923 558924 72989 558925
rect 72923 558860 72924 558924
rect 72988 558860 72989 558924
rect 72923 558859 72989 558860
rect 73659 558924 73725 558925
rect 73659 558860 73660 558924
rect 73724 558860 73725 558924
rect 73659 558859 73725 558860
rect 74211 558924 74277 558925
rect 74211 558860 74212 558924
rect 74276 558860 74277 558924
rect 74211 558859 74277 558860
rect 74947 558924 75013 558925
rect 74947 558860 74948 558924
rect 75012 558860 75013 558924
rect 74947 558859 75013 558860
rect 75683 558924 75749 558925
rect 75683 558860 75684 558924
rect 75748 558860 75749 558924
rect 75683 558859 75749 558860
rect 75870 558789 75930 560290
rect 76790 558925 76850 560290
rect 77314 559330 77374 560320
rect 77468 560290 78138 560350
rect 77314 559270 77402 559330
rect 77342 558925 77402 559270
rect 78078 558925 78138 560290
rect 78446 560290 78512 560350
rect 78636 560290 79242 560350
rect 76787 558924 76853 558925
rect 76787 558860 76788 558924
rect 76852 558860 76853 558924
rect 76787 558859 76853 558860
rect 77339 558924 77405 558925
rect 77339 558860 77340 558924
rect 77404 558860 77405 558924
rect 77339 558859 77405 558860
rect 78075 558924 78141 558925
rect 78075 558860 78076 558924
rect 78140 558860 78141 558924
rect 78075 558859 78141 558860
rect 78446 558789 78506 560290
rect 79182 558925 79242 560290
rect 79179 558924 79245 558925
rect 79179 558860 79180 558924
rect 79244 558860 79245 558924
rect 79179 558859 79245 558860
rect 79366 558789 79426 560430
rect 79804 560290 79978 560350
rect 79918 558925 79978 560290
rect 80654 560290 80848 560350
rect 80972 560290 81266 560350
rect 80654 558925 80714 560290
rect 81206 558925 81266 560290
rect 81942 560290 82016 560350
rect 82140 560290 82738 560350
rect 81942 558925 82002 560290
rect 82678 558925 82738 560290
rect 79915 558924 79981 558925
rect 79915 558860 79916 558924
rect 79980 558860 79981 558924
rect 79915 558859 79981 558860
rect 80651 558924 80717 558925
rect 80651 558860 80652 558924
rect 80716 558860 80717 558924
rect 80651 558859 80717 558860
rect 81203 558924 81269 558925
rect 81203 558860 81204 558924
rect 81268 558860 81269 558924
rect 81203 558859 81269 558860
rect 81939 558924 82005 558925
rect 81939 558860 81940 558924
rect 82004 558860 82005 558924
rect 81939 558859 82005 558860
rect 82675 558924 82741 558925
rect 82675 558860 82676 558924
rect 82740 558860 82741 558924
rect 82675 558859 82741 558860
rect 82862 558789 82922 560430
rect 83308 560290 83842 560350
rect 83782 558925 83842 560290
rect 84150 560290 84352 560350
rect 84476 560290 85130 560350
rect 84150 558925 84210 560290
rect 85070 558925 85130 560290
rect 85438 560290 85520 560350
rect 85644 560290 86234 560350
rect 83779 558924 83845 558925
rect 83779 558860 83780 558924
rect 83844 558860 83845 558924
rect 83779 558859 83845 558860
rect 84147 558924 84213 558925
rect 84147 558860 84148 558924
rect 84212 558860 84213 558924
rect 84147 558859 84213 558860
rect 85067 558924 85133 558925
rect 85067 558860 85068 558924
rect 85132 558860 85133 558924
rect 85067 558859 85133 558860
rect 85438 558789 85498 560290
rect 86174 558789 86234 560290
rect 69795 558788 69861 558789
rect 69795 558724 69796 558788
rect 69860 558724 69861 558788
rect 69795 558723 69861 558724
rect 75867 558788 75933 558789
rect 75867 558724 75868 558788
rect 75932 558724 75933 558788
rect 75867 558723 75933 558724
rect 78443 558788 78509 558789
rect 78443 558724 78444 558788
rect 78508 558724 78509 558788
rect 78443 558723 78509 558724
rect 79363 558788 79429 558789
rect 79363 558724 79364 558788
rect 79428 558724 79429 558788
rect 79363 558723 79429 558724
rect 82859 558788 82925 558789
rect 82859 558724 82860 558788
rect 82924 558724 82925 558788
rect 82859 558723 82925 558724
rect 85435 558788 85501 558789
rect 85435 558724 85436 558788
rect 85500 558724 85501 558788
rect 85435 558723 85501 558724
rect 86171 558788 86237 558789
rect 86171 558724 86172 558788
rect 86236 558724 86237 558788
rect 86171 558723 86237 558724
rect 86358 558653 86418 560430
rect 86782 559330 86842 560320
rect 87826 560010 87886 560320
rect 87980 560290 88258 560350
rect 87826 559950 87890 560010
rect 86726 559270 86842 559330
rect 86726 558925 86786 559270
rect 87830 558925 87890 559950
rect 88198 558925 88258 560290
rect 88934 560290 89024 560350
rect 88934 558925 88994 560290
rect 89118 558925 89178 560320
rect 89854 560290 90192 560350
rect 90316 560290 91018 560350
rect 89854 558925 89914 560290
rect 90958 558925 91018 560290
rect 91142 560290 91360 560350
rect 91484 560290 92122 560350
rect 86723 558924 86789 558925
rect 86723 558860 86724 558924
rect 86788 558860 86789 558924
rect 86723 558859 86789 558860
rect 87827 558924 87893 558925
rect 87827 558860 87828 558924
rect 87892 558860 87893 558924
rect 87827 558859 87893 558860
rect 88195 558924 88261 558925
rect 88195 558860 88196 558924
rect 88260 558860 88261 558924
rect 88195 558859 88261 558860
rect 88931 558924 88997 558925
rect 88931 558860 88932 558924
rect 88996 558860 88997 558924
rect 88931 558859 88997 558860
rect 89115 558924 89181 558925
rect 89115 558860 89116 558924
rect 89180 558860 89181 558924
rect 89115 558859 89181 558860
rect 89851 558924 89917 558925
rect 89851 558860 89852 558924
rect 89916 558860 89917 558924
rect 89851 558859 89917 558860
rect 90955 558924 91021 558925
rect 90955 558860 90956 558924
rect 91020 558860 91021 558924
rect 90955 558859 91021 558860
rect 91142 558789 91202 560290
rect 92062 558925 92122 560290
rect 92498 560010 92558 560320
rect 92652 560290 93226 560350
rect 92430 559950 92558 560010
rect 92430 558925 92490 559950
rect 93166 558925 93226 560290
rect 93534 560290 93696 560350
rect 92059 558924 92125 558925
rect 92059 558860 92060 558924
rect 92124 558860 92125 558924
rect 92059 558859 92125 558860
rect 92427 558924 92493 558925
rect 92427 558860 92428 558924
rect 92492 558860 92493 558924
rect 92427 558859 92493 558860
rect 93163 558924 93229 558925
rect 93163 558860 93164 558924
rect 93228 558860 93229 558924
rect 93163 558859 93229 558860
rect 91139 558788 91205 558789
rect 91139 558724 91140 558788
rect 91204 558724 91205 558788
rect 91139 558723 91205 558724
rect 93534 558653 93594 560290
rect 93790 559330 93850 560320
rect 93718 559270 93850 559330
rect 93718 558789 93778 559270
rect 94822 558925 94882 560350
rect 94988 560290 95066 560350
rect 95006 558925 95066 560290
rect 95742 560290 96032 560350
rect 96156 560290 96538 560350
rect 95742 558925 95802 560290
rect 96478 558925 96538 560290
rect 97030 560290 97200 560350
rect 97324 560290 97642 560350
rect 97030 558925 97090 560290
rect 97582 558925 97642 560290
rect 98318 558925 98378 560350
rect 98492 560290 99114 560350
rect 99054 558925 99114 560290
rect 99506 560010 99566 560320
rect 99660 560290 100218 560350
rect 99422 559950 99566 560010
rect 94819 558924 94885 558925
rect 94819 558860 94820 558924
rect 94884 558860 94885 558924
rect 94819 558859 94885 558860
rect 95003 558924 95069 558925
rect 95003 558860 95004 558924
rect 95068 558860 95069 558924
rect 95003 558859 95069 558860
rect 95739 558924 95805 558925
rect 95739 558860 95740 558924
rect 95804 558860 95805 558924
rect 95739 558859 95805 558860
rect 96475 558924 96541 558925
rect 96475 558860 96476 558924
rect 96540 558860 96541 558924
rect 96475 558859 96541 558860
rect 97027 558924 97093 558925
rect 97027 558860 97028 558924
rect 97092 558860 97093 558924
rect 97027 558859 97093 558860
rect 97579 558924 97645 558925
rect 97579 558860 97580 558924
rect 97644 558860 97645 558924
rect 97579 558859 97645 558860
rect 98315 558924 98381 558925
rect 98315 558860 98316 558924
rect 98380 558860 98381 558924
rect 98315 558859 98381 558860
rect 99051 558924 99117 558925
rect 99051 558860 99052 558924
rect 99116 558860 99117 558924
rect 99051 558859 99117 558860
rect 93715 558788 93781 558789
rect 93715 558724 93716 558788
rect 93780 558724 93781 558788
rect 93715 558723 93781 558724
rect 86355 558652 86421 558653
rect 86355 558588 86356 558652
rect 86420 558588 86421 558652
rect 86355 558587 86421 558588
rect 93531 558652 93597 558653
rect 93531 558588 93532 558652
rect 93596 558588 93597 558652
rect 93531 558587 93597 558588
rect 99422 558517 99482 559950
rect 100158 558925 100218 560290
rect 100342 560290 100704 560350
rect 100828 560290 101506 560350
rect 100155 558924 100221 558925
rect 100155 558860 100156 558924
rect 100220 558860 100221 558924
rect 100155 558859 100221 558860
rect 99419 558516 99485 558517
rect 99419 558452 99420 558516
rect 99484 558452 99485 558516
rect 99419 558451 99485 558452
rect 64275 558108 64341 558109
rect 64275 558044 64276 558108
rect 64340 558044 64341 558108
rect 64275 558043 64341 558044
rect 100342 557837 100402 560290
rect 100339 557836 100405 557837
rect 100339 557772 100340 557836
rect 100404 557772 100405 557836
rect 100339 557771 100405 557772
rect 101446 557565 101506 560290
rect 101630 560290 101872 560350
rect 101996 560290 102058 560350
rect 101630 557701 101690 560290
rect 101998 558925 102058 560290
rect 101995 558924 102061 558925
rect 101995 558860 101996 558924
rect 102060 558860 102061 558924
rect 101995 558859 102061 558860
rect 101627 557700 101693 557701
rect 101627 557636 101628 557700
rect 101692 557636 101693 557700
rect 101627 557635 101693 557636
rect 102734 557565 102794 560430
rect 103164 560290 103346 560350
rect 103286 557565 103346 560290
rect 104022 560290 104208 560350
rect 104332 560290 104818 560350
rect 104022 557565 104082 560290
rect 104758 558925 104818 560290
rect 105310 560290 105376 560350
rect 105500 560290 106106 560350
rect 104755 558924 104821 558925
rect 104755 558860 104756 558924
rect 104820 558860 104821 558924
rect 104755 558859 104821 558860
rect 105310 558789 105370 560290
rect 105307 558788 105373 558789
rect 105307 558724 105308 558788
rect 105372 558724 105373 558788
rect 105307 558723 105373 558724
rect 105310 557565 105370 558723
rect 106046 557565 106106 560290
rect 106230 557701 106290 560430
rect 106668 560290 107210 560350
rect 107150 558925 107210 560290
rect 107682 559330 107742 560320
rect 107836 560290 108498 560350
rect 107682 559270 107762 559330
rect 107147 558924 107213 558925
rect 107147 558860 107148 558924
rect 107212 558860 107213 558924
rect 107147 558859 107213 558860
rect 106227 557700 106293 557701
rect 106227 557636 106228 557700
rect 106292 557636 106293 557700
rect 106227 557635 106293 557636
rect 107702 557565 107762 559270
rect 108438 558925 108498 560290
rect 108622 560290 108880 560350
rect 108435 558924 108501 558925
rect 108435 558860 108436 558924
rect 108500 558860 108501 558924
rect 108435 558859 108501 558860
rect 108622 558517 108682 560290
rect 108619 558516 108685 558517
rect 108619 558452 108620 558516
rect 108684 558452 108685 558516
rect 108619 558451 108685 558452
rect 108990 557565 109050 560350
rect 101443 557564 101509 557565
rect 101443 557500 101444 557564
rect 101508 557500 101509 557564
rect 101443 557499 101509 557500
rect 102731 557564 102797 557565
rect 102731 557500 102732 557564
rect 102796 557500 102797 557564
rect 102731 557499 102797 557500
rect 103283 557564 103349 557565
rect 103283 557500 103284 557564
rect 103348 557500 103349 557564
rect 103283 557499 103349 557500
rect 104019 557564 104085 557565
rect 104019 557500 104020 557564
rect 104084 557500 104085 557564
rect 104019 557499 104085 557500
rect 105307 557564 105373 557565
rect 105307 557500 105308 557564
rect 105372 557500 105373 557564
rect 105307 557499 105373 557500
rect 106043 557564 106109 557565
rect 106043 557500 106044 557564
rect 106108 557500 106109 557564
rect 106043 557499 106109 557500
rect 107699 557564 107765 557565
rect 107699 557500 107700 557564
rect 107764 557500 107765 557564
rect 107699 557499 107765 557500
rect 108987 557564 109053 557565
rect 108987 557500 108988 557564
rect 109052 557500 109053 557564
rect 108987 557499 109053 557500
rect 58404 543000 59004 557000
rect 62004 543000 62604 557000
rect 65604 543000 66204 557000
rect 72804 543000 73404 557000
rect 76404 546054 77004 557000
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 543000 77004 545498
rect 80004 549654 80604 557000
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 543000 80604 549098
rect 83604 553254 84204 557000
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 543000 84204 552698
rect 90804 543000 91404 557000
rect 94404 543000 95004 557000
rect 98004 543000 98604 557000
rect 101604 543000 102204 557000
rect 108804 543000 109404 557000
rect 112404 546054 113004 557000
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 543000 113004 545498
rect 116004 549654 116604 557000
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 543000 116604 549098
rect 119604 553254 120204 557000
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 543000 120204 552698
rect 126804 543000 127404 557000
rect 130404 543000 131004 557000
rect 134004 543000 134604 557000
rect 137604 543000 138204 557000
rect 144804 543000 145404 577898
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 543000 149004 545498
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 543000 152604 549098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 543000 156204 552698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 543000 163404 559898
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 543000 167004 563498
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 543000 170604 567098
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 543000 174204 570698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 543000 181404 577898
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 654247 188604 657098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 654247 192204 660698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 654247 199404 667898
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 654247 203004 671498
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 654247 206604 675098
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 654247 210204 678698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 654247 217404 685898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654247 221004 689498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 654247 224604 657098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 654247 228204 660698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 654247 235404 667898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 654247 239004 671498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 654247 242604 675098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 654247 246204 678698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 654247 253404 685898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654247 257004 689498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 654247 260604 657098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 654247 264204 660698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 259131 652900 259197 652901
rect 259131 652836 259132 652900
rect 259196 652836 259197 652900
rect 259131 652835 259197 652836
rect 263547 652900 263613 652901
rect 263547 652836 263548 652900
rect 263612 652836 263613 652900
rect 263547 652835 263613 652836
rect 259134 651130 259194 652835
rect 258608 651070 259194 651130
rect 263550 651070 263610 652835
rect 266938 643254 267262 643276
rect 266938 643018 266982 643254
rect 267218 643018 267262 643254
rect 266938 642934 267262 643018
rect 266938 642698 266982 642934
rect 267218 642698 267262 642934
rect 266938 642676 267262 642698
rect 266938 639654 267262 639676
rect 266938 639418 266982 639654
rect 267218 639418 267262 639654
rect 266938 639334 267262 639418
rect 266938 639098 266982 639334
rect 267218 639098 267262 639334
rect 266938 639076 267262 639098
rect 266938 636054 267262 636076
rect 266938 635818 266982 636054
rect 267218 635818 267262 636054
rect 266938 635734 267262 635818
rect 266938 635498 266982 635734
rect 267218 635498 267262 635734
rect 266938 635476 267262 635498
rect 266938 632454 267262 632476
rect 266938 632218 266982 632454
rect 267218 632218 267262 632454
rect 266938 632134 267262 632218
rect 266938 631898 266982 632134
rect 267218 631898 267262 632134
rect 266938 631876 267262 631898
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 266494 625254 266814 625276
rect 266494 625018 266536 625254
rect 266772 625018 266814 625254
rect 266494 624934 266814 625018
rect 266494 624698 266536 624934
rect 266772 624698 266814 624934
rect 266494 624676 266814 624698
rect 266494 621654 266814 621676
rect 266494 621418 266536 621654
rect 266772 621418 266814 621654
rect 266494 621334 266814 621418
rect 266494 621098 266536 621334
rect 266772 621098 266814 621334
rect 266494 621076 266814 621098
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 266494 618054 266814 618076
rect 266494 617818 266536 618054
rect 266772 617818 266814 618054
rect 266494 617734 266814 617818
rect 266494 617498 266536 617734
rect 266772 617498 266814 617734
rect 266494 617476 266814 617498
rect 266494 614454 266814 614476
rect 266494 614218 266536 614454
rect 266772 614218 266814 614454
rect 266494 614134 266814 614218
rect 266494 613898 266536 614134
rect 266772 613898 266814 614134
rect 266494 613876 266814 613898
rect 266938 607254 267262 607276
rect 266938 607018 266982 607254
rect 267218 607018 267262 607254
rect 266938 606934 267262 607018
rect 266938 606698 266982 606934
rect 267218 606698 267262 606934
rect 266938 606676 267262 606698
rect 266938 603654 267262 603676
rect 266938 603418 266982 603654
rect 267218 603418 267262 603654
rect 266938 603334 267262 603418
rect 266938 603098 266982 603334
rect 267218 603098 267262 603334
rect 266938 603076 267262 603098
rect 266938 600054 267262 600076
rect 266938 599818 266982 600054
rect 267218 599818 267262 600054
rect 266938 599734 267262 599818
rect 266938 599498 266982 599734
rect 267218 599498 267262 599734
rect 266938 599476 267262 599498
rect 266938 596454 267262 596476
rect 266938 596218 266982 596454
rect 267218 596218 267262 596454
rect 266938 596134 267262 596218
rect 266938 595898 266982 596134
rect 267218 595898 267262 596134
rect 266938 595876 267262 595898
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 266494 589254 266814 589276
rect 266494 589018 266536 589254
rect 266772 589018 266814 589254
rect 266494 588934 266814 589018
rect 266494 588698 266536 588934
rect 266772 588698 266814 588934
rect 266494 588676 266814 588698
rect 266494 585654 266814 585676
rect 266494 585418 266536 585654
rect 266772 585418 266814 585654
rect 266494 585334 266814 585418
rect 266494 585098 266536 585334
rect 266772 585098 266814 585334
rect 266494 585076 266814 585098
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 266494 582054 266814 582076
rect 266494 581818 266536 582054
rect 266772 581818 266814 582054
rect 266494 581734 266814 581818
rect 266494 581498 266536 581734
rect 266772 581498 266814 581734
rect 266494 581476 266814 581498
rect 269067 580956 269133 580957
rect 269067 580892 269068 580956
rect 269132 580892 269133 580956
rect 269067 580891 269133 580892
rect 269070 579138 269130 580891
rect 266494 578454 266814 578476
rect 266494 578218 266536 578454
rect 266772 578218 266814 578454
rect 266494 578134 266814 578218
rect 266494 577898 266536 578134
rect 266772 577898 266814 578134
rect 266494 577876 266814 577898
rect 266938 571254 267262 571276
rect 266938 571018 266982 571254
rect 267218 571018 267262 571254
rect 266938 570934 267262 571018
rect 266938 570698 266982 570934
rect 267218 570698 267262 570934
rect 266938 570676 267262 570698
rect 266938 567654 267262 567676
rect 266938 567418 266982 567654
rect 267218 567418 267262 567654
rect 266938 567334 267262 567418
rect 266938 567098 266982 567334
rect 267218 567098 267262 567334
rect 266938 567076 267262 567098
rect 266938 564054 267262 564076
rect 266938 563818 266982 564054
rect 267218 563818 267262 564054
rect 266938 563734 267262 563818
rect 266938 563498 266982 563734
rect 267218 563498 267262 563734
rect 266938 563476 267262 563498
rect 207062 560430 207344 560490
rect 221046 560430 221360 560490
rect 228038 560430 228368 560490
rect 270804 560454 271404 595898
rect 193833 560290 194426 560350
rect 194366 558925 194426 560290
rect 196206 560290 196832 560350
rect 197310 560290 198000 560350
rect 198782 560290 199168 560350
rect 200254 560290 200336 560350
rect 196206 558925 196266 560290
rect 194363 558924 194429 558925
rect 194363 558860 194364 558924
rect 194428 558860 194429 558924
rect 194363 558859 194429 558860
rect 196203 558924 196269 558925
rect 196203 558860 196204 558924
rect 196268 558860 196269 558924
rect 196203 558859 196269 558860
rect 197310 558381 197370 560290
rect 197307 558380 197373 558381
rect 197307 558316 197308 558380
rect 197372 558316 197373 558380
rect 197307 558315 197373 558316
rect 198782 558245 198842 560290
rect 200254 558925 200314 560290
rect 201474 560010 201534 560320
rect 202462 560290 202672 560350
rect 201474 559950 201602 560010
rect 201542 558925 201602 559950
rect 200251 558924 200317 558925
rect 200251 558860 200252 558924
rect 200316 558860 200317 558924
rect 200251 558859 200317 558860
rect 201539 558924 201605 558925
rect 201539 558860 201540 558924
rect 201604 558860 201605 558924
rect 201539 558859 201605 558860
rect 202462 558789 202522 560290
rect 202766 559330 202826 560320
rect 202646 559270 202826 559330
rect 203750 560290 203840 560350
rect 202646 558925 202706 559270
rect 203750 558925 203810 560290
rect 203934 558925 203994 560320
rect 204854 560290 205008 560350
rect 205132 560290 205466 560350
rect 202643 558924 202709 558925
rect 202643 558860 202644 558924
rect 202708 558860 202709 558924
rect 202643 558859 202709 558860
rect 203747 558924 203813 558925
rect 203747 558860 203748 558924
rect 203812 558860 203813 558924
rect 203747 558859 203813 558860
rect 203931 558924 203997 558925
rect 203931 558860 203932 558924
rect 203996 558860 203997 558924
rect 203931 558859 203997 558860
rect 202459 558788 202525 558789
rect 202459 558724 202460 558788
rect 202524 558724 202525 558788
rect 202459 558723 202525 558724
rect 204854 558653 204914 560290
rect 205406 558925 205466 560290
rect 206142 558925 206202 560350
rect 206300 560290 206938 560350
rect 205403 558924 205469 558925
rect 205403 558860 205404 558924
rect 205468 558860 205469 558924
rect 205403 558859 205469 558860
rect 206139 558924 206205 558925
rect 206139 558860 206140 558924
rect 206204 558860 206205 558924
rect 206139 558859 206205 558860
rect 204851 558652 204917 558653
rect 204851 558588 204852 558652
rect 204916 558588 204917 558652
rect 204851 558587 204917 558588
rect 198779 558244 198845 558245
rect 198779 558180 198780 558244
rect 198844 558180 198845 558244
rect 198779 558179 198845 558180
rect 206878 557565 206938 560290
rect 207062 557701 207122 560430
rect 207468 560290 208042 560350
rect 207059 557700 207125 557701
rect 207059 557636 207060 557700
rect 207124 557636 207125 557700
rect 207059 557635 207125 557636
rect 207982 557565 208042 560290
rect 208350 560290 208512 560350
rect 208636 560290 209330 560350
rect 208350 558925 208410 560290
rect 208347 558924 208413 558925
rect 208347 558860 208348 558924
rect 208412 558860 208413 558924
rect 208347 558859 208413 558860
rect 209270 557565 209330 560290
rect 209638 557701 209698 560350
rect 209804 560290 210434 560350
rect 210374 557701 210434 560290
rect 210558 560290 210848 560350
rect 210558 558653 210618 560290
rect 210942 559330 211002 560320
rect 210926 559270 211002 559330
rect 211846 560290 212016 560350
rect 212140 560290 212458 560350
rect 210555 558652 210621 558653
rect 210555 558588 210556 558652
rect 210620 558588 210621 558652
rect 210555 558587 210621 558588
rect 209635 557700 209701 557701
rect 209635 557636 209636 557700
rect 209700 557636 209701 557700
rect 209635 557635 209701 557636
rect 210371 557700 210437 557701
rect 210371 557636 210372 557700
rect 210436 557636 210437 557700
rect 210371 557635 210437 557636
rect 210926 557565 210986 559270
rect 211846 558925 211906 560290
rect 211843 558924 211909 558925
rect 211843 558860 211844 558924
rect 211908 558860 211909 558924
rect 211843 558859 211909 558860
rect 212398 557565 212458 560290
rect 213134 558925 213194 560350
rect 213308 560290 213562 560350
rect 213131 558924 213197 558925
rect 213131 558860 213132 558924
rect 213196 558860 213197 558924
rect 213131 558859 213197 558860
rect 213502 557565 213562 560290
rect 214054 560290 214352 560350
rect 214476 560290 214850 560350
rect 214054 558925 214114 560290
rect 214051 558924 214117 558925
rect 214051 558860 214052 558924
rect 214116 558860 214117 558924
rect 214051 558859 214117 558860
rect 214790 557565 214850 560290
rect 215342 560290 215520 560350
rect 215644 560290 216322 560350
rect 215342 558925 215402 560290
rect 215339 558924 215405 558925
rect 215339 558860 215340 558924
rect 215404 558860 215405 558924
rect 215339 558859 215405 558860
rect 216262 557565 216322 560290
rect 216630 558789 216690 560350
rect 216812 560290 217426 560350
rect 216627 558788 216693 558789
rect 216627 558724 216628 558788
rect 216692 558724 216693 558788
rect 216627 558723 216693 558724
rect 217366 557701 217426 560290
rect 217550 560290 217856 560350
rect 217550 558653 217610 560290
rect 217950 559330 218010 560320
rect 217918 559270 218010 559330
rect 218838 560290 219024 560350
rect 217547 558652 217613 558653
rect 217547 558588 217548 558652
rect 217612 558588 217613 558652
rect 217547 558587 217613 558588
rect 217363 557700 217429 557701
rect 217363 557636 217364 557700
rect 217428 557636 217429 557700
rect 217363 557635 217429 557636
rect 217918 557565 217978 559270
rect 218838 558925 218898 560290
rect 219118 560010 219178 560320
rect 220126 560290 220192 560350
rect 220316 560290 220738 560350
rect 219118 559950 219266 560010
rect 218835 558924 218901 558925
rect 218835 558860 218836 558924
rect 218900 558860 218901 558924
rect 218835 558859 218901 558860
rect 219206 557565 219266 559950
rect 220126 558925 220186 560290
rect 220123 558924 220189 558925
rect 220123 558860 220124 558924
rect 220188 558860 220189 558924
rect 220123 558859 220189 558860
rect 220678 557565 220738 560290
rect 221046 558925 221106 560430
rect 221484 560290 222026 560350
rect 221043 558924 221109 558925
rect 221043 558860 221044 558924
rect 221108 558860 221109 558924
rect 221043 558859 221109 558860
rect 221966 557565 222026 560290
rect 222334 560290 222528 560350
rect 222652 560290 223314 560350
rect 222334 558925 222394 560290
rect 222331 558924 222397 558925
rect 222331 558860 222332 558924
rect 222396 558860 222397 558924
rect 222331 558859 222397 558860
rect 223254 557565 223314 560290
rect 223622 560290 223696 560350
rect 223820 560290 224418 560350
rect 223622 558925 223682 560290
rect 223619 558924 223685 558925
rect 223619 558860 223620 558924
rect 223684 558860 223685 558924
rect 223619 558859 223685 558860
rect 224358 557565 224418 560290
rect 224542 560290 224864 560350
rect 224988 560290 225706 560350
rect 224542 558925 224602 560290
rect 224539 558924 224605 558925
rect 224539 558860 224540 558924
rect 224604 558860 224605 558924
rect 224539 558859 224605 558860
rect 225646 557701 225706 560290
rect 225830 560290 226032 560350
rect 225830 559877 225890 560290
rect 226126 560010 226186 560320
rect 227118 560290 227200 560350
rect 227324 560290 227546 560350
rect 226126 559950 226258 560010
rect 225827 559876 225893 559877
rect 225827 559812 225828 559876
rect 225892 559812 225893 559876
rect 225827 559811 225893 559812
rect 225643 557700 225709 557701
rect 225643 557636 225644 557700
rect 225708 557636 225709 557700
rect 225643 557635 225709 557636
rect 226198 557565 226258 559950
rect 227118 559333 227178 560290
rect 227115 559332 227181 559333
rect 227115 559268 227116 559332
rect 227180 559268 227181 559332
rect 227115 559267 227181 559268
rect 227486 557565 227546 560290
rect 228038 558925 228098 560430
rect 228492 560290 228834 560350
rect 228035 558924 228101 558925
rect 228035 558860 228036 558924
rect 228100 558860 228101 558924
rect 228035 558859 228101 558860
rect 228774 557565 228834 560290
rect 229323 560012 229389 560013
rect 229323 559948 229324 560012
rect 229388 560010 229389 560012
rect 229506 560010 229566 560320
rect 229660 560290 230306 560350
rect 229388 559950 229566 560010
rect 229388 559948 229389 559950
rect 229323 559947 229389 559948
rect 230246 557565 230306 560290
rect 230614 560290 230704 560350
rect 230614 558517 230674 560290
rect 230611 558516 230677 558517
rect 230611 558452 230612 558516
rect 230676 558452 230677 558516
rect 230611 558451 230677 558452
rect 230798 557565 230858 560320
rect 231842 559330 231902 560320
rect 231996 560290 232698 560350
rect 231842 559270 231962 559330
rect 231902 558653 231962 559270
rect 231899 558652 231965 558653
rect 231899 558588 231900 558652
rect 231964 558588 231965 558652
rect 231899 558587 231965 558588
rect 232638 557701 232698 560290
rect 232822 560290 233040 560350
rect 232822 558789 232882 560290
rect 233134 559330 233194 560320
rect 233006 559270 233194 559330
rect 233558 560290 234208 560350
rect 234332 560290 234538 560350
rect 232819 558788 232885 558789
rect 232819 558724 232820 558788
rect 232884 558724 232885 558788
rect 232819 558723 232885 558724
rect 232635 557700 232701 557701
rect 232635 557636 232636 557700
rect 232700 557636 232701 557700
rect 232635 557635 232701 557636
rect 233006 557565 233066 559270
rect 233558 558789 233618 560290
rect 233555 558788 233621 558789
rect 233555 558724 233556 558788
rect 233620 558724 233621 558788
rect 233555 558723 233621 558724
rect 234478 557565 234538 560290
rect 234662 560290 235376 560350
rect 235500 560290 235826 560350
rect 234662 558789 234722 560290
rect 235766 558925 235826 560290
rect 236134 560290 236544 560350
rect 236668 560290 237298 560350
rect 235763 558924 235829 558925
rect 235763 558860 235764 558924
rect 235828 558860 235829 558924
rect 235763 558859 235829 558860
rect 236134 558789 236194 560290
rect 237238 558925 237298 560290
rect 237422 560290 237712 560350
rect 237836 560290 238402 560350
rect 237235 558924 237301 558925
rect 237235 558860 237236 558924
rect 237300 558860 237301 558924
rect 237235 558859 237301 558860
rect 234659 558788 234725 558789
rect 234659 558724 234660 558788
rect 234724 558724 234725 558788
rect 234659 558723 234725 558724
rect 236131 558788 236197 558789
rect 236131 558724 236132 558788
rect 236196 558724 236197 558788
rect 236131 558723 236197 558724
rect 237422 558653 237482 560290
rect 237419 558652 237485 558653
rect 237419 558588 237420 558652
rect 237484 558588 237485 558652
rect 237419 558587 237485 558588
rect 238342 558109 238402 560290
rect 238710 560290 238880 560350
rect 239004 560290 239690 560350
rect 238710 558381 238770 560290
rect 239630 558925 239690 560290
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 239627 558924 239693 558925
rect 239627 558860 239628 558924
rect 239692 558860 239693 558924
rect 239627 558859 239693 558860
rect 238707 558380 238773 558381
rect 238707 558316 238708 558380
rect 238772 558316 238773 558380
rect 238707 558315 238773 558316
rect 238339 558108 238405 558109
rect 238339 558044 238340 558108
rect 238404 558044 238405 558108
rect 238339 558043 238405 558044
rect 206875 557564 206941 557565
rect 206875 557500 206876 557564
rect 206940 557500 206941 557564
rect 206875 557499 206941 557500
rect 207979 557564 208045 557565
rect 207979 557500 207980 557564
rect 208044 557500 208045 557564
rect 207979 557499 208045 557500
rect 209267 557564 209333 557565
rect 209267 557500 209268 557564
rect 209332 557500 209333 557564
rect 209267 557499 209333 557500
rect 210923 557564 210989 557565
rect 210923 557500 210924 557564
rect 210988 557500 210989 557564
rect 210923 557499 210989 557500
rect 212395 557564 212461 557565
rect 212395 557500 212396 557564
rect 212460 557500 212461 557564
rect 212395 557499 212461 557500
rect 213499 557564 213565 557565
rect 213499 557500 213500 557564
rect 213564 557500 213565 557564
rect 213499 557499 213565 557500
rect 214787 557564 214853 557565
rect 214787 557500 214788 557564
rect 214852 557500 214853 557564
rect 214787 557499 214853 557500
rect 216259 557564 216325 557565
rect 216259 557500 216260 557564
rect 216324 557500 216325 557564
rect 216259 557499 216325 557500
rect 217915 557564 217981 557565
rect 217915 557500 217916 557564
rect 217980 557500 217981 557564
rect 217915 557499 217981 557500
rect 219203 557564 219269 557565
rect 219203 557500 219204 557564
rect 219268 557500 219269 557564
rect 219203 557499 219269 557500
rect 220675 557564 220741 557565
rect 220675 557500 220676 557564
rect 220740 557500 220741 557564
rect 220675 557499 220741 557500
rect 221963 557564 222029 557565
rect 221963 557500 221964 557564
rect 222028 557500 222029 557564
rect 221963 557499 222029 557500
rect 223251 557564 223317 557565
rect 223251 557500 223252 557564
rect 223316 557500 223317 557564
rect 223251 557499 223317 557500
rect 224355 557564 224421 557565
rect 224355 557500 224356 557564
rect 224420 557500 224421 557564
rect 224355 557499 224421 557500
rect 226195 557564 226261 557565
rect 226195 557500 226196 557564
rect 226260 557500 226261 557564
rect 226195 557499 226261 557500
rect 227483 557564 227549 557565
rect 227483 557500 227484 557564
rect 227548 557500 227549 557564
rect 227483 557499 227549 557500
rect 228771 557564 228837 557565
rect 228771 557500 228772 557564
rect 228836 557500 228837 557564
rect 228771 557499 228837 557500
rect 230243 557564 230309 557565
rect 230243 557500 230244 557564
rect 230308 557500 230309 557564
rect 230243 557499 230309 557500
rect 230795 557564 230861 557565
rect 230795 557500 230796 557564
rect 230860 557500 230861 557564
rect 230795 557499 230861 557500
rect 233003 557564 233069 557565
rect 233003 557500 233004 557564
rect 233068 557500 233069 557564
rect 233003 557499 233069 557500
rect 234475 557564 234541 557565
rect 234475 557500 234476 557564
rect 234540 557500 234541 557564
rect 234475 557499 234541 557500
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 543000 185004 545498
rect 188004 549654 188604 557000
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 543000 188604 549098
rect 191604 553254 192204 557000
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 543000 192204 552698
rect 198804 543000 199404 557000
rect 202404 543000 203004 557000
rect 206004 543000 206604 557000
rect 209604 543000 210204 557000
rect 216804 543000 217404 557000
rect 220404 546054 221004 557000
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 543000 221004 545498
rect 224004 549654 224604 557000
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 543000 224604 549098
rect 227604 553254 228204 557000
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 543000 228204 552698
rect 234804 543000 235404 557000
rect 238404 543000 239004 557000
rect 242004 543000 242604 557000
rect 245604 543000 246204 557000
rect 252804 543000 253404 557000
rect 256404 546054 257004 557000
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 543000 257004 545498
rect 260004 549654 260604 557000
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 543000 260604 549098
rect 263604 553254 264204 557000
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 543000 264204 552698
rect 270804 543000 271404 559898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 543000 275004 563498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 543000 278604 567098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 282315 648684 282381 648685
rect 282315 648620 282316 648684
rect 282380 648620 282381 648684
rect 282315 648619 282381 648620
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 543000 282204 570698
rect 79554 535254 79874 535276
rect 79554 535018 79596 535254
rect 79832 535018 79874 535254
rect 79554 534934 79874 535018
rect 79554 534698 79596 534934
rect 79832 534698 79874 534934
rect 79554 534676 79874 534698
rect 79554 531654 79874 531676
rect 79554 531418 79596 531654
rect 79832 531418 79874 531654
rect 79554 531334 79874 531418
rect 79554 531098 79596 531334
rect 79832 531098 79874 531334
rect 79554 531076 79874 531098
rect 79554 528054 79874 528076
rect 79554 527818 79596 528054
rect 79832 527818 79874 528054
rect 79554 527734 79874 527818
rect 79554 527498 79596 527734
rect 79832 527498 79874 527734
rect 79554 527476 79874 527498
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 79554 524454 79874 524476
rect 79554 524218 79596 524454
rect 79832 524218 79874 524454
rect 79554 524134 79874 524218
rect 79554 523898 79596 524134
rect 79832 523898 79874 524134
rect 79554 523876 79874 523898
rect 64194 517254 64514 517276
rect 64194 517018 64236 517254
rect 64472 517018 64514 517254
rect 64194 516934 64514 517018
rect 64194 516698 64236 516934
rect 64472 516698 64514 516934
rect 64194 516676 64514 516698
rect 64194 513654 64514 513676
rect 64194 513418 64236 513654
rect 64472 513418 64514 513654
rect 64194 513334 64514 513418
rect 64194 513098 64236 513334
rect 64472 513098 64514 513334
rect 64194 513076 64514 513098
rect 64194 510054 64514 510076
rect 64194 509818 64236 510054
rect 64472 509818 64514 510054
rect 64194 509734 64514 509818
rect 64194 509498 64236 509734
rect 64472 509498 64514 509734
rect 64194 509476 64514 509498
rect 64194 506454 64514 506476
rect 64194 506218 64236 506454
rect 64472 506218 64514 506454
rect 64194 506134 64514 506218
rect 64194 505898 64236 506134
rect 64472 505898 64514 506134
rect 64194 505876 64514 505898
rect 79554 499254 79874 499276
rect 79554 499018 79596 499254
rect 79832 499018 79874 499254
rect 79554 498934 79874 499018
rect 79554 498698 79596 498934
rect 79832 498698 79874 498934
rect 79554 498676 79874 498698
rect 79554 495654 79874 495676
rect 79554 495418 79596 495654
rect 79832 495418 79874 495654
rect 79554 495334 79874 495418
rect 79554 495098 79596 495334
rect 79832 495098 79874 495334
rect 79554 495076 79874 495098
rect 79554 492054 79874 492076
rect 79554 491818 79596 492054
rect 79832 491818 79874 492054
rect 79554 491734 79874 491818
rect 79554 491498 79596 491734
rect 79832 491498 79874 491734
rect 79554 491476 79874 491498
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 79554 488454 79874 488476
rect 79554 488218 79596 488454
rect 79832 488218 79874 488454
rect 79554 488134 79874 488218
rect 79554 487898 79596 488134
rect 79832 487898 79874 488134
rect 79554 487876 79874 487898
rect 64194 481254 64514 481276
rect 64194 481018 64236 481254
rect 64472 481018 64514 481254
rect 64194 480934 64514 481018
rect 64194 480698 64236 480934
rect 64472 480698 64514 480934
rect 64194 480676 64514 480698
rect 64194 477654 64514 477676
rect 64194 477418 64236 477654
rect 64472 477418 64514 477654
rect 64194 477334 64514 477418
rect 64194 477098 64236 477334
rect 64472 477098 64514 477334
rect 64194 477076 64514 477098
rect 64194 474054 64514 474076
rect 64194 473818 64236 474054
rect 64472 473818 64514 474054
rect 64194 473734 64514 473818
rect 64194 473498 64236 473734
rect 64472 473498 64514 473734
rect 64194 473476 64514 473498
rect 64194 470454 64514 470476
rect 64194 470218 64236 470454
rect 64472 470218 64514 470454
rect 64194 470134 64514 470218
rect 64194 469898 64236 470134
rect 64472 469898 64514 470134
rect 64194 469876 64514 469898
rect 79554 463254 79874 463276
rect 79554 463018 79596 463254
rect 79832 463018 79874 463254
rect 79554 462934 79874 463018
rect 79554 462698 79596 462934
rect 79832 462698 79874 462934
rect 79554 462676 79874 462698
rect 79554 459654 79874 459676
rect 79554 459418 79596 459654
rect 79832 459418 79874 459654
rect 79554 459334 79874 459418
rect 79554 459098 79596 459334
rect 79832 459098 79874 459334
rect 79554 459076 79874 459098
rect 79554 456054 79874 456076
rect 79554 455818 79596 456054
rect 79832 455818 79874 456054
rect 79554 455734 79874 455818
rect 79554 455498 79596 455734
rect 79832 455498 79874 455734
rect 79554 455476 79874 455498
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 79554 452454 79874 452476
rect 79554 452218 79596 452454
rect 79832 452218 79874 452454
rect 79554 452134 79874 452218
rect 79554 451898 79596 452134
rect 79832 451898 79874 452134
rect 79554 451876 79874 451898
rect 64194 445254 64514 445276
rect 64194 445018 64236 445254
rect 64472 445018 64514 445254
rect 64194 444934 64514 445018
rect 64194 444698 64236 444934
rect 64472 444698 64514 444934
rect 64194 444676 64514 444698
rect 64194 441654 64514 441676
rect 64194 441418 64236 441654
rect 64472 441418 64514 441654
rect 64194 441334 64514 441418
rect 64194 441098 64236 441334
rect 64472 441098 64514 441334
rect 64194 441076 64514 441098
rect 64194 438054 64514 438076
rect 64194 437818 64236 438054
rect 64472 437818 64514 438054
rect 64194 437734 64514 437818
rect 64194 437498 64236 437734
rect 64472 437498 64514 437734
rect 64194 437476 64514 437498
rect 64194 434454 64514 434476
rect 64194 434218 64236 434454
rect 64472 434218 64514 434454
rect 64194 434134 64514 434218
rect 64194 433898 64236 434134
rect 64472 433898 64514 434134
rect 64194 433876 64514 433898
rect 79554 427254 79874 427276
rect 79554 427018 79596 427254
rect 79832 427018 79874 427254
rect 79554 426934 79874 427018
rect 79554 426698 79596 426934
rect 79832 426698 79874 426934
rect 79554 426676 79874 426698
rect 79554 423654 79874 423676
rect 79554 423418 79596 423654
rect 79832 423418 79874 423654
rect 79554 423334 79874 423418
rect 79554 423098 79596 423334
rect 79832 423098 79874 423334
rect 79554 423076 79874 423098
rect 79554 420054 79874 420076
rect 79554 419818 79596 420054
rect 79832 419818 79874 420054
rect 79554 419734 79874 419818
rect 79554 419498 79596 419734
rect 79832 419498 79874 419734
rect 79554 419476 79874 419498
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 79554 416454 79874 416476
rect 79554 416218 79596 416454
rect 79832 416218 79874 416454
rect 79554 416134 79874 416218
rect 79554 415898 79596 416134
rect 79832 415898 79874 416134
rect 79554 415876 79874 415898
rect 64194 409254 64514 409276
rect 64194 409018 64236 409254
rect 64472 409018 64514 409254
rect 64194 408934 64514 409018
rect 64194 408698 64236 408934
rect 64472 408698 64514 408934
rect 64194 408676 64514 408698
rect 64194 405654 64514 405676
rect 64194 405418 64236 405654
rect 64472 405418 64514 405654
rect 64194 405334 64514 405418
rect 64194 405098 64236 405334
rect 64472 405098 64514 405334
rect 64194 405076 64514 405098
rect 64194 402054 64514 402076
rect 64194 401818 64236 402054
rect 64472 401818 64514 402054
rect 64194 401734 64514 401818
rect 64194 401498 64236 401734
rect 64472 401498 64514 401734
rect 64194 401476 64514 401498
rect 64194 398454 64514 398476
rect 64194 398218 64236 398454
rect 64472 398218 64514 398454
rect 64194 398134 64514 398218
rect 64194 397898 64236 398134
rect 64472 397898 64514 398134
rect 64194 397876 64514 397898
rect 79554 391254 79874 391276
rect 79554 391018 79596 391254
rect 79832 391018 79874 391254
rect 79554 390934 79874 391018
rect 79554 390698 79596 390934
rect 79832 390698 79874 390934
rect 79554 390676 79874 390698
rect 79554 387654 79874 387676
rect 79554 387418 79596 387654
rect 79832 387418 79874 387654
rect 79554 387334 79874 387418
rect 79554 387098 79596 387334
rect 79832 387098 79874 387334
rect 79554 387076 79874 387098
rect 79554 384054 79874 384076
rect 79554 383818 79596 384054
rect 79832 383818 79874 384054
rect 79554 383734 79874 383818
rect 79554 383498 79596 383734
rect 79832 383498 79874 383734
rect 79554 383476 79874 383498
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 79554 380454 79874 380476
rect 79554 380218 79596 380454
rect 79832 380218 79874 380454
rect 79554 380134 79874 380218
rect 79554 379898 79596 380134
rect 79832 379898 79874 380134
rect 79554 379876 79874 379898
rect 64194 373254 64514 373276
rect 64194 373018 64236 373254
rect 64472 373018 64514 373254
rect 64194 372934 64514 373018
rect 64194 372698 64236 372934
rect 64472 372698 64514 372934
rect 64194 372676 64514 372698
rect 64194 369654 64514 369676
rect 64194 369418 64236 369654
rect 64472 369418 64514 369654
rect 64194 369334 64514 369418
rect 64194 369098 64236 369334
rect 64472 369098 64514 369334
rect 64194 369076 64514 369098
rect 64194 366054 64514 366076
rect 64194 365818 64236 366054
rect 64472 365818 64514 366054
rect 64194 365734 64514 365818
rect 64194 365498 64236 365734
rect 64472 365498 64514 365734
rect 64194 365476 64514 365498
rect 64194 362454 64514 362476
rect 64194 362218 64236 362454
rect 64472 362218 64514 362454
rect 64194 362134 64514 362218
rect 64194 361898 64236 362134
rect 64472 361898 64514 362134
rect 64194 361876 64514 361898
rect 79554 355254 79874 355276
rect 79554 355018 79596 355254
rect 79832 355018 79874 355254
rect 79554 354934 79874 355018
rect 79554 354698 79596 354934
rect 79832 354698 79874 354934
rect 79554 354676 79874 354698
rect 79554 351654 79874 351676
rect 79554 351418 79596 351654
rect 79832 351418 79874 351654
rect 79554 351334 79874 351418
rect 79554 351098 79596 351334
rect 79832 351098 79874 351334
rect 79554 351076 79874 351098
rect 79554 348054 79874 348076
rect 79554 347818 79596 348054
rect 79832 347818 79874 348054
rect 79554 347734 79874 347818
rect 79554 347498 79596 347734
rect 79832 347498 79874 347734
rect 79554 347476 79874 347498
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 79554 344454 79874 344476
rect 79554 344218 79596 344454
rect 79832 344218 79874 344454
rect 79554 344134 79874 344218
rect 79554 343898 79596 344134
rect 79832 343898 79874 344134
rect 79554 343876 79874 343898
rect 64194 337254 64514 337276
rect 64194 337018 64236 337254
rect 64472 337018 64514 337254
rect 64194 336934 64514 337018
rect 64194 336698 64236 336934
rect 64472 336698 64514 336934
rect 64194 336676 64514 336698
rect 64194 333654 64514 333676
rect 64194 333418 64236 333654
rect 64472 333418 64514 333654
rect 64194 333334 64514 333418
rect 64194 333098 64236 333334
rect 64472 333098 64514 333334
rect 64194 333076 64514 333098
rect 64194 330054 64514 330076
rect 64194 329818 64236 330054
rect 64472 329818 64514 330054
rect 64194 329734 64514 329818
rect 64194 329498 64236 329734
rect 64472 329498 64514 329734
rect 64194 329476 64514 329498
rect 64194 326454 64514 326476
rect 64194 326218 64236 326454
rect 64472 326218 64514 326454
rect 64194 326134 64514 326218
rect 64194 325898 64236 326134
rect 64472 325898 64514 326134
rect 64194 325876 64514 325898
rect 282318 322965 282378 648619
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 282315 322964 282381 322965
rect 282315 322900 282316 322964
rect 282380 322900 282381 322964
rect 282315 322899 282381 322900
rect 144867 318476 144933 318477
rect 144867 318412 144868 318476
rect 144932 318412 144933 318476
rect 144867 318411 144933 318412
rect 144870 318205 144930 318411
rect 144867 318204 144933 318205
rect 144867 318140 144868 318204
rect 144932 318140 144933 318204
rect 144867 318139 144933 318140
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 312054 59004 317000
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 315654 62604 317000
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 283254 66204 317000
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 290454 73404 317000
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 294054 77004 317000
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 297654 80604 317000
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 83604 301254 84204 317000
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 81755 278764 81821 278765
rect 81755 278700 81756 278764
rect 81820 278700 81821 278764
rect 81755 278699 81821 278700
rect 81758 270469 81818 278699
rect 81755 270468 81821 270469
rect 81755 270404 81756 270468
rect 81820 270404 81821 270468
rect 81755 270403 81821 270404
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 308454 91404 317000
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 312054 95004 317000
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 315654 98604 317000
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 283254 102204 317000
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 290454 109404 317000
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 294054 113004 317000
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 297654 116604 317000
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 301254 120204 317000
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 126804 308454 127404 317000
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 124443 42124 124509 42125
rect 124443 42060 124444 42124
rect 124508 42060 124509 42124
rect 124443 42059 124509 42060
rect 124446 32469 124506 42059
rect 124443 32468 124509 32469
rect 124443 32404 124444 32468
rect 124508 32404 124509 32468
rect 124443 32403 124509 32404
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 312054 131004 317000
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 315654 134604 317000
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 137604 283254 138204 317000
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 135115 280124 135181 280125
rect 135115 280060 135116 280124
rect 135180 280060 135181 280124
rect 135115 280059 135181 280060
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 135118 270605 135178 280059
rect 135115 270604 135181 270605
rect 135115 270540 135116 270604
rect 135180 270540 135181 270604
rect 135115 270539 135181 270540
rect 135115 260812 135181 260813
rect 135115 260748 135116 260812
rect 135180 260748 135181 260812
rect 135115 260747 135181 260748
rect 135118 251293 135178 260747
rect 135115 251292 135181 251293
rect 135115 251228 135116 251292
rect 135180 251228 135181 251292
rect 135115 251227 135181 251228
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 135115 61436 135181 61437
rect 135115 61372 135116 61436
rect 135180 61372 135181 61436
rect 135115 61371 135181 61372
rect 135118 48381 135178 61371
rect 135115 48380 135181 48381
rect 135115 48316 135116 48380
rect 135180 48316 135181 48380
rect 135115 48315 135181 48316
rect 135115 42124 135181 42125
rect 135115 42060 135116 42124
rect 135180 42060 135181 42124
rect 135115 42059 135181 42060
rect 135118 29069 135178 42059
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 135115 29068 135181 29069
rect 135115 29004 135116 29068
rect 135180 29004 135181 29068
rect 135115 29003 135181 29004
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 290454 145404 317000
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 294054 149004 317000
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 297654 152604 317000
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 301254 156204 317000
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 308454 163404 317000
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 312054 167004 317000
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 315654 170604 317000
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 283254 174204 317000
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 290454 181404 317000
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 294054 185004 317000
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 297654 188604 317000
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 301254 192204 317000
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 308454 199404 317000
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 312054 203004 317000
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 315654 206604 317000
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 283254 210204 317000
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 290454 217404 317000
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 294054 221004 317000
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 224004 297654 224604 317000
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 222147 4452 222213 4453
rect 222147 4388 222148 4452
rect 222212 4388 222213 4452
rect 222147 4387 222213 4388
rect 222150 4181 222210 4387
rect 222147 4180 222213 4181
rect 222147 4116 222148 4180
rect 222212 4116 222213 4180
rect 222147 4115 222213 4116
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 301254 228204 317000
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 308454 235404 317000
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 312054 239004 317000
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 315654 242604 317000
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 283254 246204 317000
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 290454 253404 317000
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 249747 4588 249813 4589
rect 249747 4524 249748 4588
rect 249812 4524 249813 4588
rect 249747 4523 249813 4524
rect 249750 4317 249810 4523
rect 249747 4316 249813 4317
rect 249747 4252 249748 4316
rect 249812 4252 249813 4316
rect 249747 4251 249813 4252
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 294054 257004 317000
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 297654 260604 317000
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 301254 264204 317000
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 308454 271404 317000
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 269067 4588 269133 4589
rect 269067 4524 269068 4588
rect 269132 4524 269133 4588
rect 269067 4523 269133 4524
rect 269070 4317 269130 4523
rect 269067 4316 269133 4317
rect 269067 4252 269068 4316
rect 269132 4252 269133 4316
rect 269067 4251 269133 4252
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 312054 275004 317000
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 315654 278604 317000
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 283254 282204 317000
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 654247 307404 667898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 654247 311004 671498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 654247 314604 675098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 654247 318204 678698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 654247 325404 685898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654247 329004 689498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 654247 332604 657098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 654247 336204 660698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 654247 343404 667898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 654247 347004 671498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 654247 350604 675098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 654247 354204 678698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 654247 361404 685898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654247 365004 689498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 654247 368604 657098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 654247 372204 660698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 654247 379404 667898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 654247 383004 671498
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 654247 386604 675098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 654247 390204 678698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 378179 652900 378245 652901
rect 378179 652836 378180 652900
rect 378244 652836 378245 652900
rect 378179 652835 378245 652836
rect 383515 652900 383581 652901
rect 383515 652836 383516 652900
rect 383580 652836 383581 652900
rect 383515 652835 383581 652836
rect 378182 651130 378242 652835
rect 383518 651130 383578 652835
rect 378182 651070 378608 651130
rect 383518 651070 383603 651130
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 386938 643254 387262 643276
rect 386938 643018 386982 643254
rect 387218 643018 387262 643254
rect 386938 642934 387262 643018
rect 386938 642698 386982 642934
rect 387218 642698 387262 642934
rect 386938 642676 387262 642698
rect 386938 639654 387262 639676
rect 386938 639418 386982 639654
rect 387218 639418 387262 639654
rect 386938 639334 387262 639418
rect 386938 639098 386982 639334
rect 387218 639098 387262 639334
rect 386938 639076 387262 639098
rect 386938 636054 387262 636076
rect 386938 635818 386982 636054
rect 387218 635818 387262 636054
rect 386938 635734 387262 635818
rect 386938 635498 386982 635734
rect 387218 635498 387262 635734
rect 386938 635476 387262 635498
rect 386938 632454 387262 632476
rect 386938 632218 386982 632454
rect 387218 632218 387262 632454
rect 386938 632134 387262 632218
rect 386938 631898 386982 632134
rect 387218 631898 387262 632134
rect 386938 631876 387262 631898
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 386494 625254 386814 625276
rect 386494 625018 386536 625254
rect 386772 625018 386814 625254
rect 386494 624934 386814 625018
rect 386494 624698 386536 624934
rect 386772 624698 386814 624934
rect 386494 624676 386814 624698
rect 386494 621654 386814 621676
rect 386494 621418 386536 621654
rect 386772 621418 386814 621654
rect 386494 621334 386814 621418
rect 386494 621098 386536 621334
rect 386772 621098 386814 621334
rect 386494 621076 386814 621098
rect 386494 618054 386814 618076
rect 386494 617818 386536 618054
rect 386772 617818 386814 618054
rect 386494 617734 386814 617818
rect 386494 617498 386536 617734
rect 386772 617498 386814 617734
rect 386494 617476 386814 617498
rect 386494 614454 386814 614476
rect 386494 614218 386536 614454
rect 386772 614218 386814 614454
rect 386494 614134 386814 614218
rect 386494 613898 386536 614134
rect 386772 613898 386814 614134
rect 386494 613876 386814 613898
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 386938 607254 387262 607276
rect 386938 607018 386982 607254
rect 387218 607018 387262 607254
rect 386938 606934 387262 607018
rect 386938 606698 386982 606934
rect 387218 606698 387262 606934
rect 386938 606676 387262 606698
rect 386938 603654 387262 603676
rect 386938 603418 386982 603654
rect 387218 603418 387262 603654
rect 386938 603334 387262 603418
rect 386938 603098 386982 603334
rect 387218 603098 387262 603334
rect 386938 603076 387262 603098
rect 386938 600054 387262 600076
rect 386938 599818 386982 600054
rect 387218 599818 387262 600054
rect 386938 599734 387262 599818
rect 386938 599498 386982 599734
rect 387218 599498 387262 599734
rect 386938 599476 387262 599498
rect 386938 596454 387262 596476
rect 386938 596218 386982 596454
rect 387218 596218 387262 596454
rect 386938 596134 387262 596218
rect 386938 595898 386982 596134
rect 387218 595898 387262 596134
rect 386938 595876 387262 595898
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 386494 589254 386814 589276
rect 386494 589018 386536 589254
rect 386772 589018 386814 589254
rect 386494 588934 386814 589018
rect 386494 588698 386536 588934
rect 386772 588698 386814 588934
rect 386494 588676 386814 588698
rect 386494 585654 386814 585676
rect 386494 585418 386536 585654
rect 386772 585418 386814 585654
rect 386494 585334 386814 585418
rect 386494 585098 386536 585334
rect 386772 585098 386814 585334
rect 386494 585076 386814 585098
rect 386494 582054 386814 582076
rect 386494 581818 386536 582054
rect 386772 581818 386814 582054
rect 386494 581734 386814 581818
rect 386494 581498 386536 581734
rect 386772 581498 386814 581734
rect 386494 581476 386814 581498
rect 386494 578454 386814 578476
rect 386494 578218 386536 578454
rect 386772 578218 386814 578454
rect 386494 578134 386814 578218
rect 386494 577898 386536 578134
rect 386772 577898 386814 578134
rect 386494 577876 386814 577898
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 386938 571254 387262 571276
rect 386938 571018 386982 571254
rect 387218 571018 387262 571254
rect 386938 570934 387262 571018
rect 386938 570698 386982 570934
rect 387218 570698 387262 570934
rect 386938 570676 387262 570698
rect 386938 567654 387262 567676
rect 386938 567418 386982 567654
rect 387218 567418 387262 567654
rect 386938 567334 387262 567418
rect 386938 567098 386982 567334
rect 387218 567098 387262 567334
rect 386938 567076 387262 567098
rect 386938 564054 387262 564076
rect 386938 563818 386982 564054
rect 387218 563818 387262 564054
rect 386938 563734 387262 563818
rect 386938 563498 386982 563734
rect 387218 563498 387262 563734
rect 386938 563476 387262 563498
rect 323534 560430 323840 560490
rect 325132 560430 325434 560490
rect 313782 558925 313842 560350
rect 316174 560290 316832 560350
rect 317462 560290 318000 560350
rect 318934 560290 319168 560350
rect 316174 558925 316234 560290
rect 317462 558925 317522 560290
rect 313779 558924 313845 558925
rect 313779 558860 313780 558924
rect 313844 558860 313845 558924
rect 313779 558859 313845 558860
rect 316171 558924 316237 558925
rect 316171 558860 316172 558924
rect 316236 558860 316237 558924
rect 316171 558859 316237 558860
rect 317459 558924 317525 558925
rect 317459 558860 317460 558924
rect 317524 558860 317525 558924
rect 317459 558859 317525 558860
rect 318934 558653 318994 560290
rect 320306 560010 320366 560320
rect 320222 559950 320366 560010
rect 320958 560290 321504 560350
rect 320222 558789 320282 559950
rect 320958 558925 321018 560290
rect 322614 558925 322674 560350
rect 322796 560290 322858 560350
rect 320955 558924 321021 558925
rect 320955 558860 320956 558924
rect 321020 558860 321021 558924
rect 320955 558859 321021 558860
rect 322611 558924 322677 558925
rect 322611 558860 322612 558924
rect 322676 558860 322677 558924
rect 322611 558859 322677 558860
rect 320219 558788 320285 558789
rect 320219 558724 320220 558788
rect 320284 558724 320285 558788
rect 320219 558723 320285 558724
rect 318931 558652 318997 558653
rect 318931 558588 318932 558652
rect 318996 558588 318997 558652
rect 318931 558587 318997 558588
rect 322798 557565 322858 560290
rect 323534 558925 323594 560430
rect 323964 560290 324146 560350
rect 323531 558924 323597 558925
rect 323531 558860 323532 558924
rect 323596 558860 323597 558924
rect 323531 558859 323597 558860
rect 324086 557565 324146 560290
rect 324822 560290 325008 560350
rect 324822 557701 324882 560290
rect 324819 557700 324885 557701
rect 324819 557636 324820 557700
rect 324884 557636 324885 557700
rect 324819 557635 324885 557636
rect 325374 557565 325434 560430
rect 327030 560430 327344 560490
rect 328636 560430 328930 560490
rect 326110 560290 326176 560350
rect 326110 557701 326170 560290
rect 326107 557700 326173 557701
rect 326107 557636 326108 557700
rect 326172 557636 326173 557700
rect 326107 557635 326173 557636
rect 326294 557565 326354 560350
rect 327030 557701 327090 560430
rect 327468 560290 327642 560350
rect 327027 557700 327093 557701
rect 327027 557636 327028 557700
rect 327092 557636 327093 557700
rect 327027 557635 327093 557636
rect 327582 557565 327642 560290
rect 328482 559330 328542 560320
rect 328482 559270 328562 559330
rect 328502 558925 328562 559270
rect 328499 558924 328565 558925
rect 328499 558860 328500 558924
rect 328564 558860 328565 558924
rect 328499 558859 328565 558860
rect 328870 557565 328930 560430
rect 330526 560430 330848 560490
rect 332140 560430 332426 560490
rect 329606 560290 329680 560350
rect 329606 558925 329666 560290
rect 329603 558924 329669 558925
rect 329603 558860 329604 558924
rect 329668 558860 329669 558924
rect 329603 558859 329669 558860
rect 329790 557565 329850 560350
rect 330526 558925 330586 560430
rect 330972 560290 331138 560350
rect 330523 558924 330589 558925
rect 330523 558860 330524 558924
rect 330588 558860 330589 558924
rect 330523 558859 330589 558860
rect 331078 557701 331138 560290
rect 331814 560290 332016 560350
rect 331814 558925 331874 560290
rect 331811 558924 331877 558925
rect 331811 558860 331812 558924
rect 331876 558860 331877 558924
rect 331811 558859 331877 558860
rect 331075 557700 331141 557701
rect 331075 557636 331076 557700
rect 331140 557636 331141 557700
rect 331075 557635 331141 557636
rect 332366 557565 332426 560430
rect 334022 560430 334352 560490
rect 335644 560430 335922 560490
rect 333102 560290 333184 560350
rect 333102 558925 333162 560290
rect 333099 558924 333165 558925
rect 333099 558860 333100 558924
rect 333164 558860 333165 558924
rect 333099 558859 333165 558860
rect 333286 557565 333346 560350
rect 334022 558925 334082 560430
rect 334476 560290 334634 560350
rect 334019 558924 334085 558925
rect 334019 558860 334020 558924
rect 334084 558860 334085 558924
rect 334019 558859 334085 558860
rect 334574 557565 334634 560290
rect 335490 560010 335550 560320
rect 335490 559950 335554 560010
rect 335494 558925 335554 559950
rect 335491 558924 335557 558925
rect 335491 558860 335492 558924
rect 335556 558860 335557 558924
rect 335491 558859 335557 558860
rect 335862 557565 335922 560430
rect 339910 560430 340192 560490
rect 341484 560430 341810 560490
rect 348492 560430 348802 560490
rect 351996 560430 352298 560490
rect 355500 560430 355794 560490
rect 359004 560430 359290 560490
rect 336414 560290 336688 560350
rect 336414 558925 336474 560290
rect 336411 558924 336477 558925
rect 336411 558860 336412 558924
rect 336476 558860 336477 558924
rect 336411 558859 336477 558860
rect 336782 557565 336842 560320
rect 337702 560290 337856 560350
rect 337702 558925 337762 560290
rect 337950 559330 338010 560320
rect 337886 559270 338010 559330
rect 337699 558924 337765 558925
rect 337699 558860 337700 558924
rect 337764 558860 337765 558924
rect 337699 558859 337765 558860
rect 337886 557701 337946 559270
rect 338990 558925 339050 560350
rect 339148 560290 339234 560350
rect 338987 558924 339053 558925
rect 338987 558860 338988 558924
rect 339052 558860 339053 558924
rect 338987 558859 339053 558860
rect 337883 557700 337949 557701
rect 337883 557636 337884 557700
rect 337948 557636 337949 557700
rect 337883 557635 337949 557636
rect 339174 557565 339234 560290
rect 339910 558925 339970 560430
rect 340316 560290 340522 560350
rect 339907 558924 339973 558925
rect 339907 558860 339908 558924
rect 339972 558860 339973 558924
rect 339907 558859 339973 558860
rect 340462 557565 340522 560290
rect 341198 560290 341360 560350
rect 341198 558925 341258 560290
rect 341195 558924 341261 558925
rect 341195 558860 341196 558924
rect 341260 558860 341261 558924
rect 341195 558859 341261 558860
rect 341750 557565 341810 560430
rect 342486 558925 342546 560350
rect 342652 560290 342730 560350
rect 342483 558924 342549 558925
rect 342483 558860 342484 558924
rect 342548 558860 342549 558924
rect 342483 558859 342549 558860
rect 342670 557565 342730 560290
rect 343666 560010 343726 560320
rect 343820 560290 344018 560350
rect 343590 559950 343726 560010
rect 343590 558925 343650 559950
rect 343587 558924 343653 558925
rect 343587 558860 343588 558924
rect 343652 558860 343653 558924
rect 343587 558859 343653 558860
rect 343958 557565 344018 560290
rect 344694 560290 344864 560350
rect 344694 558925 344754 560290
rect 344958 559330 345018 560320
rect 344878 559270 345018 559330
rect 345798 560290 346032 560350
rect 346156 560290 346226 560350
rect 344691 558924 344757 558925
rect 344691 558860 344692 558924
rect 344756 558860 344757 558924
rect 344691 558859 344757 558860
rect 344878 557701 344938 559270
rect 345798 558925 345858 560290
rect 345795 558924 345861 558925
rect 345795 558860 345796 558924
rect 345860 558860 345861 558924
rect 345795 558859 345861 558860
rect 344875 557700 344941 557701
rect 344875 557636 344876 557700
rect 344940 557636 344941 557700
rect 344875 557635 344941 557636
rect 346166 557565 346226 560290
rect 346534 560290 347200 560350
rect 347324 560290 347514 560350
rect 346534 558925 346594 560290
rect 346531 558924 346597 558925
rect 346531 558860 346532 558924
rect 346596 558860 346597 558924
rect 346531 558859 346597 558860
rect 347454 557565 347514 560290
rect 348190 560290 348368 560350
rect 348190 558925 348250 560290
rect 348187 558924 348253 558925
rect 348187 558860 348188 558924
rect 348252 558860 348253 558924
rect 348187 558859 348253 558860
rect 348742 557565 348802 560430
rect 349478 558925 349538 560350
rect 349660 560290 349722 560350
rect 349475 558924 349541 558925
rect 349475 558860 349476 558924
rect 349540 558860 349541 558924
rect 349475 558859 349541 558860
rect 349662 557565 349722 560290
rect 350674 560010 350734 560320
rect 350828 560290 351010 560350
rect 350582 559950 350734 560010
rect 350582 558925 350642 559950
rect 350579 558924 350645 558925
rect 350579 558860 350580 558924
rect 350644 558860 350645 558924
rect 350579 558859 350645 558860
rect 350950 557565 351010 560290
rect 351842 559333 351902 560320
rect 351842 559332 351933 559333
rect 351842 559270 351868 559332
rect 351867 559268 351868 559270
rect 351932 559268 351933 559332
rect 351867 559267 351933 559268
rect 322795 557564 322861 557565
rect 322795 557500 322796 557564
rect 322860 557500 322861 557564
rect 322795 557499 322861 557500
rect 324083 557564 324149 557565
rect 324083 557500 324084 557564
rect 324148 557500 324149 557564
rect 324083 557499 324149 557500
rect 325371 557564 325437 557565
rect 325371 557500 325372 557564
rect 325436 557500 325437 557564
rect 325371 557499 325437 557500
rect 326291 557564 326357 557565
rect 326291 557500 326292 557564
rect 326356 557500 326357 557564
rect 326291 557499 326357 557500
rect 327579 557564 327645 557565
rect 327579 557500 327580 557564
rect 327644 557500 327645 557564
rect 327579 557499 327645 557500
rect 328867 557564 328933 557565
rect 328867 557500 328868 557564
rect 328932 557500 328933 557564
rect 328867 557499 328933 557500
rect 329787 557564 329853 557565
rect 329787 557500 329788 557564
rect 329852 557500 329853 557564
rect 329787 557499 329853 557500
rect 332363 557564 332429 557565
rect 332363 557500 332364 557564
rect 332428 557500 332429 557564
rect 332363 557499 332429 557500
rect 333283 557564 333349 557565
rect 333283 557500 333284 557564
rect 333348 557500 333349 557564
rect 333283 557499 333349 557500
rect 334571 557564 334637 557565
rect 334571 557500 334572 557564
rect 334636 557500 334637 557564
rect 334571 557499 334637 557500
rect 335859 557564 335925 557565
rect 335859 557500 335860 557564
rect 335924 557500 335925 557564
rect 335859 557499 335925 557500
rect 336779 557564 336845 557565
rect 336779 557500 336780 557564
rect 336844 557500 336845 557564
rect 336779 557499 336845 557500
rect 339171 557564 339237 557565
rect 339171 557500 339172 557564
rect 339236 557500 339237 557564
rect 339171 557499 339237 557500
rect 340459 557564 340525 557565
rect 340459 557500 340460 557564
rect 340524 557500 340525 557564
rect 340459 557499 340525 557500
rect 341747 557564 341813 557565
rect 341747 557500 341748 557564
rect 341812 557500 341813 557564
rect 341747 557499 341813 557500
rect 342667 557564 342733 557565
rect 342667 557500 342668 557564
rect 342732 557500 342733 557564
rect 342667 557499 342733 557500
rect 343955 557564 344021 557565
rect 343955 557500 343956 557564
rect 344020 557500 344021 557564
rect 343955 557499 344021 557500
rect 346163 557564 346229 557565
rect 346163 557500 346164 557564
rect 346228 557500 346229 557564
rect 346163 557499 346229 557500
rect 347451 557564 347517 557565
rect 347451 557500 347452 557564
rect 347516 557500 347517 557564
rect 347451 557499 347517 557500
rect 348739 557564 348805 557565
rect 348739 557500 348740 557564
rect 348804 557500 348805 557564
rect 348739 557499 348805 557500
rect 349659 557564 349725 557565
rect 349659 557500 349660 557564
rect 349724 557500 349725 557564
rect 349659 557499 349725 557500
rect 350947 557564 351013 557565
rect 350947 557500 350948 557564
rect 351012 557500 351013 557564
rect 350947 557499 351013 557500
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 306804 524454 307404 557000
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 414247 307404 415898
rect 310404 528054 311004 557000
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 414247 311004 419498
rect 314004 531654 314604 557000
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 414247 314604 423098
rect 317604 535254 318204 557000
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 414247 318204 426698
rect 324804 542454 325404 557000
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 414247 325404 433898
rect 328404 546054 329004 557000
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 414247 329004 437498
rect 332004 549654 332604 557000
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 414247 332604 441098
rect 335604 553254 336204 557000
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 414247 336204 444698
rect 342804 524454 343404 557000
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 414247 343404 415898
rect 346404 528054 347004 557000
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 414247 347004 419498
rect 350004 531654 350604 557000
rect 352238 555525 352298 560430
rect 352422 560290 353040 560350
rect 352422 558925 352482 560290
rect 352419 558924 352485 558925
rect 352419 558860 352420 558924
rect 352484 558860 352485 558924
rect 352419 558859 352485 558860
rect 353158 557701 353218 560350
rect 353526 560290 354208 560350
rect 354332 560290 354506 560350
rect 353526 558925 353586 560290
rect 353523 558924 353589 558925
rect 353523 558860 353524 558924
rect 353588 558860 353589 558924
rect 353523 558859 353589 558860
rect 353155 557700 353221 557701
rect 353155 557636 353156 557700
rect 353220 557636 353221 557700
rect 353155 557635 353221 557636
rect 354446 557565 354506 560290
rect 354814 560290 355376 560350
rect 354814 558789 354874 560290
rect 354811 558788 354877 558789
rect 354811 558724 354812 558788
rect 354876 558724 354877 558788
rect 354811 558723 354877 558724
rect 355734 557565 355794 560430
rect 356102 560290 356544 560350
rect 356102 558789 356162 560290
rect 356099 558788 356165 558789
rect 356099 558724 356100 558788
rect 356164 558724 356165 558788
rect 356099 558723 356165 558724
rect 356654 557565 356714 560350
rect 357682 560010 357742 560320
rect 357836 560290 358002 560350
rect 357574 559950 357742 560010
rect 357574 558517 357634 559950
rect 357571 558516 357637 558517
rect 357571 558452 357572 558516
rect 357636 558452 357637 558516
rect 357571 558451 357637 558452
rect 357942 557565 358002 560290
rect 358850 559333 358910 560320
rect 358850 559332 358925 559333
rect 358850 559270 358860 559332
rect 358859 559268 358860 559270
rect 358924 559268 358925 559332
rect 358859 559267 358925 559268
rect 354443 557564 354509 557565
rect 354443 557500 354444 557564
rect 354508 557500 354509 557564
rect 354443 557499 354509 557500
rect 355731 557564 355797 557565
rect 355731 557500 355732 557564
rect 355796 557500 355797 557564
rect 355731 557499 355797 557500
rect 356651 557564 356717 557565
rect 356651 557500 356652 557564
rect 356716 557500 356717 557564
rect 356651 557499 356717 557500
rect 357939 557564 358005 557565
rect 357939 557500 357940 557564
rect 358004 557500 358005 557564
rect 357939 557499 358005 557500
rect 352235 555524 352301 555525
rect 352235 555460 352236 555524
rect 352300 555460 352301 555524
rect 352235 555459 352301 555460
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 414247 350604 423098
rect 353604 535254 354204 557000
rect 359230 555525 359290 560430
rect 359227 555524 359293 555525
rect 359227 555460 359228 555524
rect 359292 555460 359293 555524
rect 359227 555459 359293 555460
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 414247 354204 426698
rect 360804 542454 361404 557000
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 414247 361404 433898
rect 364404 546054 365004 557000
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 414247 365004 437498
rect 368004 549654 368604 557000
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 414247 368604 441098
rect 371604 553254 372204 557000
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 414247 372204 444698
rect 378804 524454 379404 557000
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 414247 379404 415898
rect 382404 528054 383004 557000
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 414247 383004 419498
rect 386004 531654 386604 557000
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 414247 386604 423098
rect 389604 535254 390204 557000
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 414247 390204 426698
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 383515 413268 383581 413269
rect 383515 413204 383516 413268
rect 383580 413204 383581 413268
rect 383515 413203 383581 413204
rect 383518 411770 383578 413203
rect 383433 411710 383578 411770
rect 383433 411060 383493 411710
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 310482 409254 310802 409276
rect 310482 409018 310524 409254
rect 310760 409018 310802 409254
rect 310482 408934 310802 409018
rect 310482 408698 310524 408934
rect 310760 408698 310802 408934
rect 310482 408676 310802 408698
rect 310482 405654 310802 405676
rect 310482 405418 310524 405654
rect 310760 405418 310802 405654
rect 310482 405334 310802 405418
rect 310482 405098 310524 405334
rect 310760 405098 310802 405334
rect 310482 405076 310802 405098
rect 310482 402054 310802 402076
rect 310482 401818 310524 402054
rect 310760 401818 310802 402054
rect 310482 401734 310802 401818
rect 310482 401498 310524 401734
rect 310760 401498 310802 401734
rect 310482 401476 310802 401498
rect 310482 398454 310802 398476
rect 310482 398218 310524 398454
rect 310760 398218 310802 398454
rect 310482 398134 310802 398218
rect 310482 397898 310524 398134
rect 310760 397898 310802 398134
rect 310482 397876 310802 397898
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 310034 391254 310358 391276
rect 310034 391018 310078 391254
rect 310314 391018 310358 391254
rect 310034 390934 310358 391018
rect 310034 390698 310078 390934
rect 310314 390698 310358 390934
rect 310034 390676 310358 390698
rect 310034 387654 310358 387676
rect 310034 387418 310078 387654
rect 310314 387418 310358 387654
rect 310034 387334 310358 387418
rect 310034 387098 310078 387334
rect 310314 387098 310358 387334
rect 310034 387076 310358 387098
rect 310034 384054 310358 384076
rect 310034 383818 310078 384054
rect 310314 383818 310358 384054
rect 310034 383734 310358 383818
rect 310034 383498 310078 383734
rect 310314 383498 310358 383734
rect 310034 383476 310358 383498
rect 310034 380454 310358 380476
rect 310034 380218 310078 380454
rect 310314 380218 310358 380454
rect 310034 380134 310358 380218
rect 310034 379898 310078 380134
rect 310314 379898 310358 380134
rect 310034 379876 310358 379898
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 310482 373254 310802 373276
rect 310482 373018 310524 373254
rect 310760 373018 310802 373254
rect 310482 372934 310802 373018
rect 310482 372698 310524 372934
rect 310760 372698 310802 372934
rect 310482 372676 310802 372698
rect 310482 369654 310802 369676
rect 310482 369418 310524 369654
rect 310760 369418 310802 369654
rect 310482 369334 310802 369418
rect 310482 369098 310524 369334
rect 310760 369098 310802 369334
rect 310482 369076 310802 369098
rect 310482 366054 310802 366076
rect 310482 365818 310524 366054
rect 310760 365818 310802 366054
rect 310482 365734 310802 365818
rect 310482 365498 310524 365734
rect 310760 365498 310802 365734
rect 310482 365476 310802 365498
rect 310482 362454 310802 362476
rect 310482 362218 310524 362454
rect 310760 362218 310802 362454
rect 310482 362134 310802 362218
rect 310482 361898 310524 362134
rect 310760 361898 310802 362134
rect 310482 361876 310802 361898
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 310034 355254 310358 355276
rect 310034 355018 310078 355254
rect 310314 355018 310358 355254
rect 310034 354934 310358 355018
rect 310034 354698 310078 354934
rect 310314 354698 310358 354934
rect 310034 354676 310358 354698
rect 310034 351654 310358 351676
rect 310034 351418 310078 351654
rect 310314 351418 310358 351654
rect 310034 351334 310358 351418
rect 310034 351098 310078 351334
rect 310314 351098 310358 351334
rect 310034 351076 310358 351098
rect 310034 348054 310358 348076
rect 310034 347818 310078 348054
rect 310314 347818 310358 348054
rect 310034 347734 310358 347818
rect 310034 347498 310078 347734
rect 310314 347498 310358 347734
rect 310034 347476 310358 347498
rect 310034 344454 310358 344476
rect 310034 344218 310078 344454
rect 310314 344218 310358 344454
rect 310034 344134 310358 344218
rect 310034 343898 310078 344134
rect 310314 343898 310358 344134
rect 310034 343876 310358 343898
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 310482 337254 310802 337276
rect 310482 337018 310524 337254
rect 310760 337018 310802 337254
rect 310482 336934 310802 337018
rect 310482 336698 310524 336934
rect 310760 336698 310802 336934
rect 310482 336676 310802 336698
rect 310482 333654 310802 333676
rect 310482 333418 310524 333654
rect 310760 333418 310802 333654
rect 310482 333334 310802 333418
rect 310482 333098 310524 333334
rect 310760 333098 310802 333334
rect 310482 333076 310802 333098
rect 310482 330054 310802 330076
rect 310482 329818 310524 330054
rect 310760 329818 310802 330054
rect 310482 329734 310802 329818
rect 310482 329498 310524 329734
rect 310760 329498 310802 329734
rect 310482 329476 310802 329498
rect 310482 326454 310802 326476
rect 310482 326218 310524 326454
rect 310760 326218 310802 326454
rect 310482 326134 310802 326218
rect 310482 325898 310524 326134
rect 310760 325898 310802 326134
rect 310482 325876 310802 325898
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 313414 320250 313693 320310
rect 313414 318749 313474 320250
rect 313411 318748 313477 318749
rect 313411 318684 313412 318748
rect 313476 318684 313477 318748
rect 313411 318683 313477 318684
rect 320771 318340 320837 318341
rect 320771 318276 320772 318340
rect 320836 318276 320837 318340
rect 320771 318275 320837 318276
rect 311203 318204 311269 318205
rect 311203 318140 311204 318204
rect 311268 318140 311269 318204
rect 311203 318139 311269 318140
rect 306804 308454 307404 317000
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 303000 307404 307898
rect 310404 312054 311004 317000
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 303000 311004 311498
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 56454 307404 77000
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 60054 311004 77000
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 311206 3365 311266 318139
rect 314004 315654 314604 317000
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 303000 314604 315098
rect 317604 303000 318204 317000
rect 314194 294054 314514 294076
rect 314194 293818 314236 294054
rect 314472 293818 314514 294054
rect 314194 293734 314514 293818
rect 314194 293498 314236 293734
rect 314472 293498 314514 293734
rect 314194 293476 314514 293498
rect 314194 290454 314514 290476
rect 314194 290218 314236 290454
rect 314472 290218 314514 290454
rect 314194 290134 314514 290218
rect 314194 289898 314236 290134
rect 314472 289898 314514 290134
rect 314194 289876 314514 289898
rect 314194 265254 314514 265276
rect 314194 265018 314236 265254
rect 314472 265018 314514 265254
rect 314194 264934 314514 265018
rect 314194 264698 314236 264934
rect 314472 264698 314514 264934
rect 314194 264676 314514 264698
rect 314194 261654 314514 261676
rect 314194 261418 314236 261654
rect 314472 261418 314514 261654
rect 314194 261334 314514 261418
rect 314194 261098 314236 261334
rect 314472 261098 314514 261334
rect 314194 261076 314514 261098
rect 314194 258054 314514 258076
rect 314194 257818 314236 258054
rect 314472 257818 314514 258054
rect 314194 257734 314514 257818
rect 314194 257498 314236 257734
rect 314472 257498 314514 257734
rect 314194 257476 314514 257498
rect 314194 254454 314514 254476
rect 314194 254218 314236 254454
rect 314472 254218 314514 254454
rect 314194 254134 314514 254218
rect 314194 253898 314236 254134
rect 314472 253898 314514 254134
rect 314194 253876 314514 253898
rect 314194 229254 314514 229276
rect 314194 229018 314236 229254
rect 314472 229018 314514 229254
rect 314194 228934 314514 229018
rect 314194 228698 314236 228934
rect 314472 228698 314514 228934
rect 314194 228676 314514 228698
rect 314194 225654 314514 225676
rect 314194 225418 314236 225654
rect 314472 225418 314514 225654
rect 314194 225334 314514 225418
rect 314194 225098 314236 225334
rect 314472 225098 314514 225334
rect 314194 225076 314514 225098
rect 314194 222054 314514 222076
rect 314194 221818 314236 222054
rect 314472 221818 314514 222054
rect 314194 221734 314514 221818
rect 314194 221498 314236 221734
rect 314472 221498 314514 221734
rect 314194 221476 314514 221498
rect 314194 218454 314514 218476
rect 314194 218218 314236 218454
rect 314472 218218 314514 218454
rect 314194 218134 314514 218218
rect 314194 217898 314236 218134
rect 314472 217898 314514 218134
rect 314194 217876 314514 217898
rect 314194 193254 314514 193276
rect 314194 193018 314236 193254
rect 314472 193018 314514 193254
rect 314194 192934 314514 193018
rect 314194 192698 314236 192934
rect 314472 192698 314514 192934
rect 314194 192676 314514 192698
rect 314194 189654 314514 189676
rect 314194 189418 314236 189654
rect 314472 189418 314514 189654
rect 314194 189334 314514 189418
rect 314194 189098 314236 189334
rect 314472 189098 314514 189334
rect 314194 189076 314514 189098
rect 314194 186054 314514 186076
rect 314194 185818 314236 186054
rect 314472 185818 314514 186054
rect 314194 185734 314514 185818
rect 314194 185498 314236 185734
rect 314472 185498 314514 185734
rect 314194 185476 314514 185498
rect 314194 182454 314514 182476
rect 314194 182218 314236 182454
rect 314472 182218 314514 182454
rect 314194 182134 314514 182218
rect 314194 181898 314236 182134
rect 314472 181898 314514 182134
rect 314194 181876 314514 181898
rect 314194 157254 314514 157276
rect 314194 157018 314236 157254
rect 314472 157018 314514 157254
rect 314194 156934 314514 157018
rect 314194 156698 314236 156934
rect 314472 156698 314514 156934
rect 314194 156676 314514 156698
rect 314194 153654 314514 153676
rect 314194 153418 314236 153654
rect 314472 153418 314514 153654
rect 314194 153334 314514 153418
rect 314194 153098 314236 153334
rect 314472 153098 314514 153334
rect 314194 153076 314514 153098
rect 314194 150054 314514 150076
rect 314194 149818 314236 150054
rect 314472 149818 314514 150054
rect 314194 149734 314514 149818
rect 314194 149498 314236 149734
rect 314472 149498 314514 149734
rect 314194 149476 314514 149498
rect 314194 146454 314514 146476
rect 314194 146218 314236 146454
rect 314472 146218 314514 146454
rect 314194 146134 314514 146218
rect 314194 145898 314236 146134
rect 314472 145898 314514 146134
rect 314194 145876 314514 145898
rect 314194 121254 314514 121276
rect 314194 121018 314236 121254
rect 314472 121018 314514 121254
rect 314194 120934 314514 121018
rect 314194 120698 314236 120934
rect 314472 120698 314514 120934
rect 314194 120676 314514 120698
rect 314194 117654 314514 117676
rect 314194 117418 314236 117654
rect 314472 117418 314514 117654
rect 314194 117334 314514 117418
rect 314194 117098 314236 117334
rect 314472 117098 314514 117334
rect 314194 117076 314514 117098
rect 314194 114054 314514 114076
rect 314194 113818 314236 114054
rect 314472 113818 314514 114054
rect 314194 113734 314514 113818
rect 314194 113498 314236 113734
rect 314472 113498 314514 113734
rect 314194 113476 314514 113498
rect 314194 110454 314514 110476
rect 314194 110218 314236 110454
rect 314472 110218 314514 110454
rect 314194 110134 314514 110218
rect 314194 109898 314236 110134
rect 314472 109898 314514 110134
rect 314194 109876 314514 109898
rect 314194 85254 314514 85276
rect 314194 85018 314236 85254
rect 314472 85018 314514 85254
rect 314194 84934 314514 85018
rect 314194 84698 314236 84934
rect 314472 84698 314514 84934
rect 314194 84676 314514 84698
rect 314004 63654 314604 77000
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 311203 3364 311269 3365
rect 311203 3300 311204 3364
rect 311268 3300 311269 3364
rect 311203 3299 311269 3300
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 67254 318204 77000
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 320774 3093 320834 318275
rect 321507 318068 321573 318069
rect 321507 318004 321508 318068
rect 321572 318004 321573 318068
rect 321507 318003 321573 318004
rect 321510 3365 321570 318003
rect 324804 303000 325404 317000
rect 328404 303000 329004 317000
rect 332004 303000 332604 317000
rect 335604 303000 336204 317000
rect 342804 308454 343404 317000
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 303000 343404 307898
rect 346404 312054 347004 317000
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 303000 347004 311498
rect 350004 315654 350604 317000
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 303000 350604 315098
rect 353604 303000 354204 317000
rect 360804 303000 361404 317000
rect 364404 303000 365004 317000
rect 368004 303000 368604 317000
rect 371604 303000 372204 317000
rect 378804 308454 379404 317000
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 303000 379404 307898
rect 382404 312054 383004 317000
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 303000 383004 311498
rect 386004 315654 386604 317000
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 303000 386604 315098
rect 389604 303000 390204 317000
rect 396804 303000 397404 325898
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 303000 401004 329498
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 303000 404604 333098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 303000 408204 336698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 303000 415404 307898
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 303000 419004 311498
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 303000 422604 315098
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 303000 426204 318698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654247 437004 689498
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 654247 440604 657098
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 654247 444204 660698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 654247 451404 667898
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 654247 455004 671498
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 654247 458604 675098
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 654247 462204 678698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 654247 469404 685898
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654247 473004 689498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 654247 476604 657098
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 654247 480204 660698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 654247 487404 667898
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 654247 491004 671498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 654247 494604 675098
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 654247 498204 678698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 654247 505404 685898
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654247 509004 689498
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 654247 512604 657098
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 654247 516204 660698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 508451 652900 508517 652901
rect 508451 652836 508452 652900
rect 508516 652836 508517 652900
rect 508451 652835 508517 652836
rect 513419 652900 513485 652901
rect 513419 652836 513420 652900
rect 513484 652836 513485 652900
rect 513419 652835 513485 652836
rect 508454 651130 508514 652835
rect 513422 651130 513482 652835
rect 508454 651070 508608 651130
rect 513422 651070 513603 651130
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 516938 643254 517262 643276
rect 516938 643018 516982 643254
rect 517218 643018 517262 643254
rect 516938 642934 517262 643018
rect 516938 642698 516982 642934
rect 517218 642698 517262 642934
rect 516938 642676 517262 642698
rect 516938 639654 517262 639676
rect 516938 639418 516982 639654
rect 517218 639418 517262 639654
rect 516938 639334 517262 639418
rect 516938 639098 516982 639334
rect 517218 639098 517262 639334
rect 516938 639076 517262 639098
rect 516938 636054 517262 636076
rect 516938 635818 516982 636054
rect 517218 635818 517262 636054
rect 516938 635734 517262 635818
rect 516938 635498 516982 635734
rect 517218 635498 517262 635734
rect 516938 635476 517262 635498
rect 516938 632454 517262 632476
rect 516938 632218 516982 632454
rect 517218 632218 517262 632454
rect 516938 632134 517262 632218
rect 516938 631898 516982 632134
rect 517218 631898 517262 632134
rect 516938 631876 517262 631898
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 516494 625254 516814 625276
rect 516494 625018 516536 625254
rect 516772 625018 516814 625254
rect 516494 624934 516814 625018
rect 516494 624698 516536 624934
rect 516772 624698 516814 624934
rect 516494 624676 516814 624698
rect 516494 621654 516814 621676
rect 516494 621418 516536 621654
rect 516772 621418 516814 621654
rect 516494 621334 516814 621418
rect 516494 621098 516536 621334
rect 516772 621098 516814 621334
rect 516494 621076 516814 621098
rect 516494 618054 516814 618076
rect 516494 617818 516536 618054
rect 516772 617818 516814 618054
rect 516494 617734 516814 617818
rect 516494 617498 516536 617734
rect 516772 617498 516814 617734
rect 516494 617476 516814 617498
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 516494 614454 516814 614476
rect 516494 614218 516536 614454
rect 516772 614218 516814 614454
rect 516494 614134 516814 614218
rect 516494 613898 516536 614134
rect 516772 613898 516814 614134
rect 516494 613876 516814 613898
rect 516938 607254 517262 607276
rect 516938 607018 516982 607254
rect 517218 607018 517262 607254
rect 516938 606934 517262 607018
rect 516938 606698 516982 606934
rect 517218 606698 517262 606934
rect 516938 606676 517262 606698
rect 516938 603654 517262 603676
rect 516938 603418 516982 603654
rect 517218 603418 517262 603654
rect 516938 603334 517262 603418
rect 516938 603098 516982 603334
rect 517218 603098 517262 603334
rect 516938 603076 517262 603098
rect 516938 600054 517262 600076
rect 516938 599818 516982 600054
rect 517218 599818 517262 600054
rect 516938 599734 517262 599818
rect 516938 599498 516982 599734
rect 517218 599498 517262 599734
rect 516938 599476 517262 599498
rect 516938 596454 517262 596476
rect 516938 596218 516982 596454
rect 517218 596218 517262 596454
rect 516938 596134 517262 596218
rect 516938 595898 516982 596134
rect 517218 595898 517262 596134
rect 516938 595876 517262 595898
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 516494 589254 516814 589276
rect 516494 589018 516536 589254
rect 516772 589018 516814 589254
rect 516494 588934 516814 589018
rect 516494 588698 516536 588934
rect 516772 588698 516814 588934
rect 516494 588676 516814 588698
rect 516494 585654 516814 585676
rect 516494 585418 516536 585654
rect 516772 585418 516814 585654
rect 516494 585334 516814 585418
rect 516494 585098 516536 585334
rect 516772 585098 516814 585334
rect 516494 585076 516814 585098
rect 516494 582054 516814 582076
rect 516494 581818 516536 582054
rect 516772 581818 516814 582054
rect 516494 581734 516814 581818
rect 516494 581498 516536 581734
rect 516772 581498 516814 581734
rect 516494 581476 516814 581498
rect 518939 580956 519005 580957
rect 518939 580892 518940 580956
rect 519004 580892 519005 580956
rect 518939 580891 519005 580892
rect 518942 579818 519002 580891
rect 440006 579189 440066 579582
rect 440003 579188 440069 579189
rect 440003 579124 440004 579188
rect 440068 579124 440069 579188
rect 440003 579123 440069 579124
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 516494 578454 516814 578476
rect 516494 578218 516536 578454
rect 516772 578218 516814 578454
rect 516494 578134 516814 578218
rect 516494 577898 516536 578134
rect 516772 577898 516814 578134
rect 516494 577876 516814 577898
rect 516938 571254 517262 571276
rect 516938 571018 516982 571254
rect 517218 571018 517262 571254
rect 516938 570934 517262 571018
rect 516938 570698 516982 570934
rect 517218 570698 517262 570934
rect 516938 570676 517262 570698
rect 516938 567654 517262 567676
rect 516938 567418 516982 567654
rect 517218 567418 517262 567654
rect 516938 567334 517262 567418
rect 516938 567098 516982 567334
rect 517218 567098 517262 567334
rect 516938 567076 517262 567098
rect 516938 564054 517262 564076
rect 516938 563818 516982 564054
rect 517218 563818 517262 564054
rect 516938 563734 517262 563818
rect 516938 563498 516982 563734
rect 517218 563498 517262 563734
rect 516938 563476 517262 563498
rect 454726 560430 455008 560490
rect 456300 560430 456626 560490
rect 443134 560290 443833 560350
rect 446262 560290 446832 560350
rect 447734 560290 448000 560350
rect 448470 560290 449168 560350
rect 449942 560290 450336 560350
rect 451414 560290 451504 560350
rect 443134 558925 443194 560290
rect 446262 558925 446322 560290
rect 447734 558925 447794 560290
rect 443131 558924 443197 558925
rect 443131 558860 443132 558924
rect 443196 558860 443197 558924
rect 443131 558859 443197 558860
rect 446259 558924 446325 558925
rect 446259 558860 446260 558924
rect 446324 558860 446325 558924
rect 446259 558859 446325 558860
rect 447731 558924 447797 558925
rect 447731 558860 447732 558924
rect 447796 558860 447797 558924
rect 447731 558859 447797 558860
rect 448470 558245 448530 560290
rect 449942 558517 450002 560290
rect 449939 558516 450005 558517
rect 449939 558452 449940 558516
rect 450004 558452 450005 558516
rect 449939 558451 450005 558452
rect 448467 558244 448533 558245
rect 448467 558180 448468 558244
rect 448532 558180 448533 558244
rect 448467 558179 448533 558180
rect 451414 558109 451474 560290
rect 452642 559330 452702 560320
rect 452796 560290 452946 560350
rect 452642 559270 452762 559330
rect 452702 558653 452762 559270
rect 452699 558652 452765 558653
rect 452699 558588 452700 558652
rect 452764 558588 452765 558652
rect 452699 558587 452765 558588
rect 451411 558108 451477 558109
rect 451411 558044 451412 558108
rect 451476 558044 451477 558108
rect 451411 558043 451477 558044
rect 452886 557565 452946 560290
rect 453622 560290 453840 560350
rect 453622 558925 453682 560290
rect 453934 559330 453994 560320
rect 453806 559270 453994 559330
rect 453619 558924 453685 558925
rect 453619 558860 453620 558924
rect 453684 558860 453685 558924
rect 453619 558859 453685 558860
rect 453806 558789 453866 559270
rect 454726 558925 454786 560430
rect 455132 560290 455338 560350
rect 454723 558924 454789 558925
rect 454723 558860 454724 558924
rect 454788 558860 454789 558924
rect 454723 558859 454789 558860
rect 453803 558788 453869 558789
rect 453803 558724 453804 558788
rect 453868 558724 453869 558788
rect 453803 558723 453869 558724
rect 455278 557565 455338 560290
rect 456014 560290 456176 560350
rect 456014 558925 456074 560290
rect 456011 558924 456077 558925
rect 456011 558860 456012 558924
rect 456076 558860 456077 558924
rect 456011 558859 456077 558860
rect 456566 557565 456626 560430
rect 458222 560430 458512 560490
rect 459804 560430 460122 560490
rect 463308 560430 463618 560490
rect 457302 558925 457362 560350
rect 457468 560290 457546 560350
rect 457299 558924 457365 558925
rect 457299 558860 457300 558924
rect 457364 558860 457365 558924
rect 457299 558859 457365 558860
rect 457486 557565 457546 560290
rect 458222 558925 458282 560430
rect 458636 560290 458834 560350
rect 458219 558924 458285 558925
rect 458219 558860 458220 558924
rect 458284 558860 458285 558924
rect 458219 558859 458285 558860
rect 458774 557565 458834 560290
rect 459510 560290 459680 560350
rect 459510 558653 459570 560290
rect 459507 558652 459573 558653
rect 459507 558588 459508 558652
rect 459572 558588 459573 558652
rect 459507 558587 459573 558588
rect 460062 557565 460122 560430
rect 460798 558925 460858 560350
rect 460972 560290 461042 560350
rect 460795 558924 460861 558925
rect 460795 558860 460796 558924
rect 460860 558860 460861 558924
rect 460795 558859 460861 558860
rect 460982 557565 461042 560290
rect 461718 560290 462016 560350
rect 461718 558925 461778 560290
rect 462110 559330 462170 560320
rect 462086 559270 462170 559330
rect 462638 560290 463184 560350
rect 461715 558924 461781 558925
rect 461715 558860 461716 558924
rect 461780 558860 461781 558924
rect 461715 558859 461781 558860
rect 462086 557701 462146 559270
rect 462638 558925 462698 560290
rect 462635 558924 462701 558925
rect 462635 558860 462636 558924
rect 462700 558860 462701 558924
rect 462635 558859 462701 558860
rect 462083 557700 462149 557701
rect 462083 557636 462084 557700
rect 462148 557636 462149 557700
rect 462083 557635 462149 557636
rect 463558 557565 463618 560430
rect 465214 560430 465520 560490
rect 468710 560430 469024 560490
rect 472206 560430 472528 560490
rect 473820 560430 474106 560490
rect 464294 558925 464354 560350
rect 464476 560290 464538 560350
rect 464291 558924 464357 558925
rect 464291 558860 464292 558924
rect 464356 558860 464357 558924
rect 464291 558859 464357 558860
rect 464478 557565 464538 560290
rect 465214 558925 465274 560430
rect 465644 560290 465826 560350
rect 465211 558924 465277 558925
rect 465211 558860 465212 558924
rect 465276 558860 465277 558924
rect 465211 558859 465277 558860
rect 465766 557565 465826 560290
rect 466502 560290 466688 560350
rect 466502 558789 466562 560290
rect 466782 560010 466842 560320
rect 467790 560290 467856 560350
rect 466782 559950 466930 560010
rect 466870 558925 466930 559950
rect 466867 558924 466933 558925
rect 466867 558860 466868 558924
rect 466932 558860 466933 558924
rect 466867 558859 466933 558860
rect 466499 558788 466565 558789
rect 466499 558724 466500 558788
rect 466564 558724 466565 558788
rect 466499 558723 466565 558724
rect 467790 558653 467850 560290
rect 467974 558925 468034 560350
rect 468710 558925 468770 560430
rect 469118 559330 469178 560320
rect 469078 559270 469178 559330
rect 469998 560290 470192 560350
rect 467971 558924 468037 558925
rect 467971 558860 467972 558924
rect 468036 558860 468037 558924
rect 467971 558859 468037 558860
rect 468707 558924 468773 558925
rect 468707 558860 468708 558924
rect 468772 558860 468773 558924
rect 468707 558859 468773 558860
rect 469078 558789 469138 559270
rect 469998 558789 470058 560290
rect 470286 560010 470346 560320
rect 471286 560290 471360 560350
rect 470286 559950 470426 560010
rect 470366 558925 470426 559950
rect 470363 558924 470429 558925
rect 470363 558860 470364 558924
rect 470428 558860 470429 558924
rect 470363 558859 470429 558860
rect 471286 558789 471346 560290
rect 471470 558925 471530 560350
rect 471467 558924 471533 558925
rect 471467 558860 471468 558924
rect 471532 558860 471533 558924
rect 471467 558859 471533 558860
rect 472206 558789 472266 560430
rect 472652 560290 472818 560350
rect 472758 558925 472818 560290
rect 473494 560290 473696 560350
rect 472755 558924 472821 558925
rect 472755 558860 472756 558924
rect 472820 558860 472821 558924
rect 472755 558859 472821 558860
rect 469075 558788 469141 558789
rect 469075 558724 469076 558788
rect 469140 558724 469141 558788
rect 469075 558723 469141 558724
rect 469995 558788 470061 558789
rect 469995 558724 469996 558788
rect 470060 558724 470061 558788
rect 469995 558723 470061 558724
rect 471283 558788 471349 558789
rect 471283 558724 471284 558788
rect 471348 558724 471349 558788
rect 471283 558723 471349 558724
rect 472203 558788 472269 558789
rect 472203 558724 472204 558788
rect 472268 558724 472269 558788
rect 472203 558723 472269 558724
rect 473494 558653 473554 560290
rect 474046 558925 474106 560430
rect 481590 560430 481872 560490
rect 483164 560430 483490 560490
rect 486668 560430 486986 560490
rect 474782 560290 474864 560350
rect 474782 558925 474842 560290
rect 474043 558924 474109 558925
rect 474043 558860 474044 558924
rect 474108 558860 474109 558924
rect 474043 558859 474109 558860
rect 474779 558924 474845 558925
rect 474779 558860 474780 558924
rect 474844 558860 474845 558924
rect 474779 558859 474845 558860
rect 467787 558652 467853 558653
rect 467787 558588 467788 558652
rect 467852 558588 467853 558652
rect 467787 558587 467853 558588
rect 473491 558652 473557 558653
rect 473491 558588 473492 558652
rect 473556 558588 473557 558652
rect 473491 558587 473557 558588
rect 474966 558381 475026 560350
rect 475518 560290 476032 560350
rect 476156 560290 476314 560350
rect 475518 558925 475578 560290
rect 475515 558924 475581 558925
rect 475515 558860 475516 558924
rect 475580 558860 475581 558924
rect 475515 558859 475581 558860
rect 476254 558381 476314 560290
rect 477170 560010 477230 560320
rect 477294 560010 477354 560320
rect 478278 560290 478368 560350
rect 477170 559950 477234 560010
rect 477294 559950 477418 560010
rect 477174 558925 477234 559950
rect 477171 558924 477237 558925
rect 477171 558860 477172 558924
rect 477236 558860 477237 558924
rect 477171 558859 477237 558860
rect 477358 558517 477418 559950
rect 478278 558925 478338 560290
rect 478275 558924 478341 558925
rect 478275 558860 478276 558924
rect 478340 558860 478341 558924
rect 478275 558859 478341 558860
rect 477355 558516 477421 558517
rect 477355 558452 477356 558516
rect 477420 558452 477421 558516
rect 477355 558451 477421 558452
rect 478462 558381 478522 560320
rect 479014 560290 479536 560350
rect 479660 560290 479810 560350
rect 479014 558925 479074 560290
rect 479011 558924 479077 558925
rect 479011 558860 479012 558924
rect 479076 558860 479077 558924
rect 479011 558859 479077 558860
rect 474963 558380 475029 558381
rect 474963 558316 474964 558380
rect 475028 558316 475029 558380
rect 474963 558315 475029 558316
rect 476251 558380 476317 558381
rect 476251 558316 476252 558380
rect 476316 558316 476317 558380
rect 476251 558315 476317 558316
rect 478459 558380 478525 558381
rect 478459 558316 478460 558380
rect 478524 558316 478525 558380
rect 478459 558315 478525 558316
rect 479750 558245 479810 560290
rect 480486 560290 480704 560350
rect 480828 560290 480914 560350
rect 480486 558789 480546 560290
rect 480854 558925 480914 560290
rect 480851 558924 480917 558925
rect 480851 558860 480852 558924
rect 480916 558860 480917 558924
rect 480851 558859 480917 558860
rect 481590 558789 481650 560430
rect 481996 560290 482202 560350
rect 480483 558788 480549 558789
rect 480483 558724 480484 558788
rect 480548 558724 480549 558788
rect 480483 558723 480549 558724
rect 481587 558788 481653 558789
rect 481587 558724 481588 558788
rect 481652 558724 481653 558788
rect 481587 558723 481653 558724
rect 482142 558517 482202 560290
rect 483010 559330 483070 560320
rect 483010 559270 483122 559330
rect 482139 558516 482205 558517
rect 482139 558452 482140 558516
rect 482204 558452 482205 558516
rect 482139 558451 482205 558452
rect 479747 558244 479813 558245
rect 479747 558180 479748 558244
rect 479812 558180 479813 558244
rect 479747 558179 479813 558180
rect 483062 557701 483122 559270
rect 483430 558245 483490 560430
rect 483614 560290 484208 560350
rect 483614 558925 483674 560290
rect 484302 559330 484362 560320
rect 484166 559270 484362 559330
rect 484718 560290 485376 560350
rect 485500 560290 485698 560350
rect 483611 558924 483677 558925
rect 483611 558860 483612 558924
rect 483676 558860 483677 558924
rect 483611 558859 483677 558860
rect 483427 558244 483493 558245
rect 483427 558180 483428 558244
rect 483492 558180 483493 558244
rect 483427 558179 483493 558180
rect 484166 558109 484226 559270
rect 484718 558653 484778 560290
rect 484715 558652 484781 558653
rect 484715 558588 484716 558652
rect 484780 558588 484781 558652
rect 484715 558587 484781 558588
rect 485638 558245 485698 560290
rect 486006 560290 486544 560350
rect 486006 558517 486066 560290
rect 486003 558516 486069 558517
rect 486003 558452 486004 558516
rect 486068 558452 486069 558516
rect 486003 558451 486069 558452
rect 486926 558245 486986 560430
rect 522804 560454 523404 595898
rect 487294 560290 487712 560350
rect 487836 560290 487906 560350
rect 487294 558517 487354 560290
rect 487291 558516 487357 558517
rect 487291 558452 487292 558516
rect 487356 558452 487357 558516
rect 487291 558451 487357 558452
rect 485635 558244 485701 558245
rect 485635 558180 485636 558244
rect 485700 558180 485701 558244
rect 485635 558179 485701 558180
rect 486923 558244 486989 558245
rect 486923 558180 486924 558244
rect 486988 558180 486989 558244
rect 486923 558179 486989 558180
rect 484163 558108 484229 558109
rect 484163 558044 484164 558108
rect 484228 558044 484229 558108
rect 484163 558043 484229 558044
rect 487846 557973 487906 560290
rect 488582 560290 488880 560350
rect 489004 560290 489194 560350
rect 488582 558653 488642 560290
rect 488579 558652 488645 558653
rect 488579 558588 488580 558652
rect 488644 558588 488645 558652
rect 488579 558587 488645 558588
rect 489134 558109 489194 560290
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 489131 558108 489197 558109
rect 489131 558044 489132 558108
rect 489196 558044 489197 558108
rect 489131 558043 489197 558044
rect 487843 557972 487909 557973
rect 487843 557908 487844 557972
rect 487908 557908 487909 557972
rect 487843 557907 487909 557908
rect 483059 557700 483125 557701
rect 483059 557636 483060 557700
rect 483124 557636 483125 557700
rect 483059 557635 483125 557636
rect 452883 557564 452949 557565
rect 452883 557500 452884 557564
rect 452948 557500 452949 557564
rect 452883 557499 452949 557500
rect 455275 557564 455341 557565
rect 455275 557500 455276 557564
rect 455340 557500 455341 557564
rect 455275 557499 455341 557500
rect 456563 557564 456629 557565
rect 456563 557500 456564 557564
rect 456628 557500 456629 557564
rect 456563 557499 456629 557500
rect 457483 557564 457549 557565
rect 457483 557500 457484 557564
rect 457548 557500 457549 557564
rect 457483 557499 457549 557500
rect 458771 557564 458837 557565
rect 458771 557500 458772 557564
rect 458836 557500 458837 557564
rect 458771 557499 458837 557500
rect 460059 557564 460125 557565
rect 460059 557500 460060 557564
rect 460124 557500 460125 557564
rect 460059 557499 460125 557500
rect 460979 557564 461045 557565
rect 460979 557500 460980 557564
rect 461044 557500 461045 557564
rect 460979 557499 461045 557500
rect 463555 557564 463621 557565
rect 463555 557500 463556 557564
rect 463620 557500 463621 557564
rect 463555 557499 463621 557500
rect 464475 557564 464541 557565
rect 464475 557500 464476 557564
rect 464540 557500 464541 557564
rect 464475 557499 464541 557500
rect 465763 557564 465829 557565
rect 465763 557500 465764 557564
rect 465828 557500 465829 557564
rect 465763 557499 465829 557500
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 436404 546054 437004 557000
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 414247 437004 437498
rect 440004 549654 440604 557000
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 414247 440604 441098
rect 443604 553254 444204 557000
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 414247 444204 444698
rect 450804 524454 451404 557000
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 414247 451404 415898
rect 454404 528054 455004 557000
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 414247 455004 419498
rect 458004 531654 458604 557000
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 414247 458604 423098
rect 461604 535254 462204 557000
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 414247 462204 426698
rect 468804 542454 469404 557000
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 414247 469404 433898
rect 472404 546054 473004 557000
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 414247 473004 437498
rect 476004 549654 476604 557000
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 414247 476604 441098
rect 479604 553254 480204 557000
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 414247 480204 444698
rect 486804 524454 487404 557000
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 414247 487404 415898
rect 490404 528054 491004 557000
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 414247 491004 419498
rect 494004 531654 494604 557000
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 414247 494604 423098
rect 497604 535254 498204 557000
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 414247 498204 426698
rect 504804 542454 505404 557000
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 414247 505404 433898
rect 508404 546054 509004 557000
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 414247 509004 437498
rect 512004 549654 512604 557000
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 414247 512604 441098
rect 515604 553254 516204 557000
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 414247 516204 444698
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 513419 412724 513485 412725
rect 513419 412660 513420 412724
rect 513484 412660 513485 412724
rect 513419 412659 513485 412660
rect 513422 411090 513482 412659
rect 513422 411030 513603 411090
rect 516494 405654 516814 405676
rect 516494 405418 516536 405654
rect 516772 405418 516814 405654
rect 516494 405334 516814 405418
rect 516494 405098 516536 405334
rect 516772 405098 516814 405334
rect 516494 405076 516814 405098
rect 516494 402054 516814 402076
rect 516494 401818 516536 402054
rect 516772 401818 516814 402054
rect 516494 401734 516814 401818
rect 516494 401498 516536 401734
rect 516772 401498 516814 401734
rect 516494 401476 516814 401498
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 516494 398454 516814 398476
rect 516494 398218 516536 398454
rect 516772 398218 516814 398454
rect 516494 398134 516814 398218
rect 516494 397898 516536 398134
rect 516772 397898 516814 398134
rect 516494 397876 516814 397898
rect 516938 391254 517262 391276
rect 516938 391018 516982 391254
rect 517218 391018 517262 391254
rect 516938 390934 517262 391018
rect 516938 390698 516982 390934
rect 517218 390698 517262 390934
rect 516938 390676 517262 390698
rect 516938 387654 517262 387676
rect 516938 387418 516982 387654
rect 517218 387418 517262 387654
rect 516938 387334 517262 387418
rect 516938 387098 516982 387334
rect 517218 387098 517262 387334
rect 516938 387076 517262 387098
rect 516938 384054 517262 384076
rect 516938 383818 516982 384054
rect 517218 383818 517262 384054
rect 516938 383734 517262 383818
rect 516938 383498 516982 383734
rect 517218 383498 517262 383734
rect 516938 383476 517262 383498
rect 516938 380454 517262 380476
rect 516938 380218 516982 380454
rect 517218 380218 517262 380454
rect 516938 380134 517262 380218
rect 516938 379898 516982 380134
rect 517218 379898 517262 380134
rect 516938 379876 517262 379898
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 516494 373254 516814 373276
rect 516494 373018 516536 373254
rect 516772 373018 516814 373254
rect 516494 372934 516814 373018
rect 516494 372698 516536 372934
rect 516772 372698 516814 372934
rect 516494 372676 516814 372698
rect 516494 369654 516814 369676
rect 516494 369418 516536 369654
rect 516772 369418 516814 369654
rect 516494 369334 516814 369418
rect 516494 369098 516536 369334
rect 516772 369098 516814 369334
rect 516494 369076 516814 369098
rect 516494 366054 516814 366076
rect 516494 365818 516536 366054
rect 516772 365818 516814 366054
rect 516494 365734 516814 365818
rect 516494 365498 516536 365734
rect 516772 365498 516814 365734
rect 516494 365476 516814 365498
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 516494 362454 516814 362476
rect 516494 362218 516536 362454
rect 516772 362218 516814 362454
rect 516494 362134 516814 362218
rect 516494 361898 516536 362134
rect 516772 361898 516814 362134
rect 516494 361876 516814 361898
rect 516938 355254 517262 355276
rect 516938 355018 516982 355254
rect 517218 355018 517262 355254
rect 516938 354934 517262 355018
rect 516938 354698 516982 354934
rect 517218 354698 517262 354934
rect 516938 354676 517262 354698
rect 516938 351654 517262 351676
rect 516938 351418 516982 351654
rect 517218 351418 517262 351654
rect 516938 351334 517262 351418
rect 516938 351098 516982 351334
rect 517218 351098 517262 351334
rect 516938 351076 517262 351098
rect 516938 348054 517262 348076
rect 516938 347818 516982 348054
rect 517218 347818 517262 348054
rect 516938 347734 517262 347818
rect 516938 347498 516982 347734
rect 517218 347498 517262 347734
rect 516938 347476 517262 347498
rect 516938 344454 517262 344476
rect 516938 344218 516982 344454
rect 517218 344218 517262 344454
rect 516938 344134 517262 344218
rect 516938 343898 516982 344134
rect 517218 343898 517262 344134
rect 516938 343876 517262 343898
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 516494 337254 516814 337276
rect 516494 337018 516536 337254
rect 516772 337018 516814 337254
rect 516494 336934 516814 337018
rect 516494 336698 516536 336934
rect 516772 336698 516814 336934
rect 516494 336676 516814 336698
rect 516494 333654 516814 333676
rect 516494 333418 516536 333654
rect 516772 333418 516814 333654
rect 516494 333334 516814 333418
rect 516494 333098 516536 333334
rect 516772 333098 516814 333334
rect 516494 333076 516814 333098
rect 516494 330054 516814 330076
rect 516494 329818 516536 330054
rect 516772 329818 516814 330054
rect 516494 329734 516814 329818
rect 516494 329498 516536 329734
rect 516772 329498 516814 329734
rect 516494 329476 516814 329498
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 303000 433404 325898
rect 516494 326454 516814 326476
rect 516494 326218 516536 326454
rect 516772 326218 516814 326454
rect 516494 326134 516814 326218
rect 516494 325898 516536 326134
rect 516772 325898 516814 326134
rect 516494 325876 516814 325898
rect 443134 320250 443833 320310
rect 443134 318749 443194 320250
rect 443131 318748 443197 318749
rect 443131 318684 443132 318748
rect 443196 318684 443197 318748
rect 443131 318683 443197 318684
rect 436404 303000 437004 317000
rect 440004 303000 440604 317000
rect 443604 303000 444204 317000
rect 450804 308454 451404 317000
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 303000 451404 307898
rect 454404 312054 455004 317000
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 303000 455004 311498
rect 458004 315654 458604 317000
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 303000 458604 315098
rect 461604 303000 462204 317000
rect 468804 303000 469404 317000
rect 472404 303000 473004 317000
rect 476004 303000 476604 317000
rect 479604 303000 480204 317000
rect 486804 308454 487404 317000
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 303000 487404 307898
rect 490404 312054 491004 317000
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 303000 491004 311498
rect 494004 315654 494604 317000
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 303000 494604 315098
rect 497604 303000 498204 317000
rect 504804 303000 505404 317000
rect 508404 303000 509004 317000
rect 512004 303000 512604 317000
rect 515604 303000 516204 317000
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 303000 523404 307898
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 303000 527004 311498
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 303000 530604 315098
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 329554 283254 329874 283276
rect 329554 283018 329596 283254
rect 329832 283018 329874 283254
rect 329554 282934 329874 283018
rect 329554 282698 329596 282934
rect 329832 282698 329874 282934
rect 329554 282676 329874 282698
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 329554 279654 329874 279676
rect 329554 279418 329596 279654
rect 329832 279418 329874 279654
rect 329554 279334 329874 279418
rect 329554 279098 329596 279334
rect 329832 279098 329874 279334
rect 329554 279076 329874 279098
rect 329554 276054 329874 276076
rect 329554 275818 329596 276054
rect 329832 275818 329874 276054
rect 329554 275734 329874 275818
rect 329554 275498 329596 275734
rect 329832 275498 329874 275734
rect 329554 275476 329874 275498
rect 329554 272454 329874 272476
rect 329554 272218 329596 272454
rect 329832 272218 329874 272454
rect 329554 272134 329874 272218
rect 329554 271898 329596 272134
rect 329832 271898 329874 272134
rect 329554 271876 329874 271898
rect 329554 247254 329874 247276
rect 329554 247018 329596 247254
rect 329832 247018 329874 247254
rect 329554 246934 329874 247018
rect 329554 246698 329596 246934
rect 329832 246698 329874 246934
rect 329554 246676 329874 246698
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 329554 243654 329874 243676
rect 329554 243418 329596 243654
rect 329832 243418 329874 243654
rect 329554 243334 329874 243418
rect 329554 243098 329596 243334
rect 329832 243098 329874 243334
rect 329554 243076 329874 243098
rect 329554 240054 329874 240076
rect 329554 239818 329596 240054
rect 329832 239818 329874 240054
rect 329554 239734 329874 239818
rect 329554 239498 329596 239734
rect 329832 239498 329874 239734
rect 329554 239476 329874 239498
rect 329554 236454 329874 236476
rect 329554 236218 329596 236454
rect 329832 236218 329874 236454
rect 329554 236134 329874 236218
rect 329554 235898 329596 236134
rect 329832 235898 329874 236134
rect 329554 235876 329874 235898
rect 329554 211254 329874 211276
rect 329554 211018 329596 211254
rect 329832 211018 329874 211254
rect 329554 210934 329874 211018
rect 329554 210698 329596 210934
rect 329832 210698 329874 210934
rect 329554 210676 329874 210698
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 329554 207654 329874 207676
rect 329554 207418 329596 207654
rect 329832 207418 329874 207654
rect 329554 207334 329874 207418
rect 329554 207098 329596 207334
rect 329832 207098 329874 207334
rect 329554 207076 329874 207098
rect 329554 204054 329874 204076
rect 329554 203818 329596 204054
rect 329832 203818 329874 204054
rect 329554 203734 329874 203818
rect 329554 203498 329596 203734
rect 329832 203498 329874 203734
rect 329554 203476 329874 203498
rect 329554 200454 329874 200476
rect 329554 200218 329596 200454
rect 329832 200218 329874 200454
rect 329554 200134 329874 200218
rect 329554 199898 329596 200134
rect 329832 199898 329874 200134
rect 329554 199876 329874 199898
rect 329554 175254 329874 175276
rect 329554 175018 329596 175254
rect 329832 175018 329874 175254
rect 329554 174934 329874 175018
rect 329554 174698 329596 174934
rect 329832 174698 329874 174934
rect 329554 174676 329874 174698
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 329554 171654 329874 171676
rect 329554 171418 329596 171654
rect 329832 171418 329874 171654
rect 329554 171334 329874 171418
rect 329554 171098 329596 171334
rect 329832 171098 329874 171334
rect 329554 171076 329874 171098
rect 329554 168054 329874 168076
rect 329554 167818 329596 168054
rect 329832 167818 329874 168054
rect 329554 167734 329874 167818
rect 329554 167498 329596 167734
rect 329832 167498 329874 167734
rect 329554 167476 329874 167498
rect 329554 164454 329874 164476
rect 329554 164218 329596 164454
rect 329832 164218 329874 164454
rect 329554 164134 329874 164218
rect 329554 163898 329596 164134
rect 329832 163898 329874 164134
rect 329554 163876 329874 163898
rect 329554 139254 329874 139276
rect 329554 139018 329596 139254
rect 329832 139018 329874 139254
rect 329554 138934 329874 139018
rect 329554 138698 329596 138934
rect 329832 138698 329874 138934
rect 329554 138676 329874 138698
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 329554 135654 329874 135676
rect 329554 135418 329596 135654
rect 329832 135418 329874 135654
rect 329554 135334 329874 135418
rect 329554 135098 329596 135334
rect 329832 135098 329874 135334
rect 329554 135076 329874 135098
rect 329554 132054 329874 132076
rect 329554 131818 329596 132054
rect 329832 131818 329874 132054
rect 329554 131734 329874 131818
rect 329554 131498 329596 131734
rect 329832 131498 329874 131734
rect 329554 131476 329874 131498
rect 329554 128454 329874 128476
rect 329554 128218 329596 128454
rect 329832 128218 329874 128454
rect 329554 128134 329874 128218
rect 329554 127898 329596 128134
rect 329832 127898 329874 128134
rect 329554 127876 329874 127898
rect 329554 103254 329874 103276
rect 329554 103018 329596 103254
rect 329832 103018 329874 103254
rect 329554 102934 329874 103018
rect 329554 102698 329596 102934
rect 329832 102698 329874 102934
rect 329554 102676 329874 102698
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 329554 99654 329874 99676
rect 329554 99418 329596 99654
rect 329832 99418 329874 99654
rect 329554 99334 329874 99418
rect 329554 99098 329596 99334
rect 329832 99098 329874 99334
rect 329554 99076 329874 99098
rect 329554 96054 329874 96076
rect 329554 95818 329596 96054
rect 329832 95818 329874 96054
rect 329554 95734 329874 95818
rect 329554 95498 329596 95734
rect 329832 95498 329874 95734
rect 329554 95476 329874 95498
rect 329554 92454 329874 92476
rect 329554 92218 329596 92454
rect 329832 92218 329874 92454
rect 329554 92134 329874 92218
rect 329554 91898 329596 92134
rect 329832 91898 329874 92134
rect 329554 91876 329874 91898
rect 324804 74454 325404 77000
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 321507 3364 321573 3365
rect 321507 3300 321508 3364
rect 321572 3300 321573 3364
rect 321507 3299 321573 3300
rect 320771 3092 320837 3093
rect 320771 3028 320772 3092
rect 320836 3028 320837 3092
rect 320771 3027 320837 3028
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 42054 329004 77000
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 45654 332604 77000
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 49254 336204 77000
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 56454 343404 77000
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 60054 347004 77000
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 63654 350604 77000
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 67254 354204 77000
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 74454 361404 77000
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 42054 365004 77000
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 45654 368604 77000
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 49254 372204 77000
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 56454 379404 77000
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 60054 383004 77000
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 63654 386604 77000
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 67254 390204 77000
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 74454 397404 77000
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 42054 401004 77000
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 45654 404604 77000
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 49254 408204 77000
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 56454 415404 77000
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 60054 419004 77000
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 63654 422604 77000
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 67254 426204 77000
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 74454 433404 77000
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 42054 437004 77000
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 45654 440604 77000
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 49254 444204 77000
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 56454 451404 77000
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 60054 455004 77000
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 63654 458604 77000
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 67254 462204 77000
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 74454 469404 77000
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 42054 473004 77000
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 45654 476604 77000
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 49254 480204 77000
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 56454 487404 77000
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 60054 491004 77000
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 63654 494604 77000
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 67254 498204 77000
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 74454 505404 77000
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 42054 509004 77000
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 45654 512604 77000
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 49254 516204 77000
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 56454 523404 77000
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 60054 527004 77000
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 63654 530604 77000
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 136982 643018 137218 643254
rect 136982 642698 137218 642934
rect 136982 639418 137218 639654
rect 136982 639098 137218 639334
rect 136982 635818 137218 636054
rect 136982 635498 137218 635734
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 136982 632218 137218 632454
rect 136982 631898 137218 632134
rect 136536 625018 136772 625254
rect 136536 624698 136772 624934
rect 136536 621418 136772 621654
rect 136536 621098 136772 621334
rect 136536 617818 136772 618054
rect 136536 617498 136772 617734
rect 136536 614218 136772 614454
rect 136536 613898 136772 614134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 136982 607018 137218 607254
rect 136982 606698 137218 606934
rect 136982 603418 137218 603654
rect 136982 603098 137218 603334
rect 136982 599818 137218 600054
rect 136982 599498 137218 599734
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 136982 596218 137218 596454
rect 136982 595898 137218 596134
rect 136536 589018 136772 589254
rect 136536 588698 136772 588934
rect 136536 585418 136772 585654
rect 136536 585098 136772 585334
rect 136536 581818 136772 582054
rect 136536 581498 136772 581734
rect 60510 579052 60746 579138
rect 60510 578988 60596 579052
rect 60596 578988 60660 579052
rect 60660 578988 60746 579052
rect 60510 578902 60746 578988
rect 137422 578902 137658 579138
rect 136536 578218 136772 578454
rect 136536 577898 136772 578134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 136982 571018 137218 571254
rect 136982 570698 137218 570934
rect 136982 567418 137218 567654
rect 136982 567098 137218 567334
rect 136982 563818 137218 564054
rect 136982 563498 137218 563734
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 266982 643018 267218 643254
rect 266982 642698 267218 642934
rect 266982 639418 267218 639654
rect 266982 639098 267218 639334
rect 266982 635818 267218 636054
rect 266982 635498 267218 635734
rect 266982 632218 267218 632454
rect 266982 631898 267218 632134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 266536 625018 266772 625254
rect 266536 624698 266772 624934
rect 266536 621418 266772 621654
rect 266536 621098 266772 621334
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 266536 617818 266772 618054
rect 266536 617498 266772 617734
rect 266536 614218 266772 614454
rect 266536 613898 266772 614134
rect 266982 607018 267218 607254
rect 266982 606698 267218 606934
rect 266982 603418 267218 603654
rect 266982 603098 267218 603334
rect 266982 599818 267218 600054
rect 266982 599498 267218 599734
rect 266982 596218 267218 596454
rect 266982 595898 267218 596134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 266536 589018 266772 589254
rect 266536 588698 266772 588934
rect 266536 585418 266772 585654
rect 266536 585098 266772 585334
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 266536 581818 266772 582054
rect 266536 581498 266772 581734
rect 190046 579052 190282 579138
rect 190046 578988 190132 579052
rect 190132 578988 190196 579052
rect 190196 578988 190282 579052
rect 190046 578902 190282 578988
rect 268982 578902 269218 579138
rect 266536 578218 266772 578454
rect 266536 577898 266772 578134
rect 266982 571018 267218 571254
rect 266982 570698 267218 570934
rect 266982 567418 267218 567654
rect 266982 567098 267218 567334
rect 266982 563818 267218 564054
rect 266982 563498 267218 563734
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 79596 535018 79832 535254
rect 79596 534698 79832 534934
rect 79596 531418 79832 531654
rect 79596 531098 79832 531334
rect 79596 527818 79832 528054
rect 79596 527498 79832 527734
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 79596 524218 79832 524454
rect 79596 523898 79832 524134
rect 64236 517018 64472 517254
rect 64236 516698 64472 516934
rect 64236 513418 64472 513654
rect 64236 513098 64472 513334
rect 64236 509818 64472 510054
rect 64236 509498 64472 509734
rect 64236 506218 64472 506454
rect 64236 505898 64472 506134
rect 79596 499018 79832 499254
rect 79596 498698 79832 498934
rect 79596 495418 79832 495654
rect 79596 495098 79832 495334
rect 79596 491818 79832 492054
rect 79596 491498 79832 491734
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 79596 488218 79832 488454
rect 79596 487898 79832 488134
rect 64236 481018 64472 481254
rect 64236 480698 64472 480934
rect 64236 477418 64472 477654
rect 64236 477098 64472 477334
rect 64236 473818 64472 474054
rect 64236 473498 64472 473734
rect 64236 470218 64472 470454
rect 64236 469898 64472 470134
rect 79596 463018 79832 463254
rect 79596 462698 79832 462934
rect 79596 459418 79832 459654
rect 79596 459098 79832 459334
rect 79596 455818 79832 456054
rect 79596 455498 79832 455734
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 79596 452218 79832 452454
rect 79596 451898 79832 452134
rect 64236 445018 64472 445254
rect 64236 444698 64472 444934
rect 64236 441418 64472 441654
rect 64236 441098 64472 441334
rect 64236 437818 64472 438054
rect 64236 437498 64472 437734
rect 64236 434218 64472 434454
rect 64236 433898 64472 434134
rect 79596 427018 79832 427254
rect 79596 426698 79832 426934
rect 79596 423418 79832 423654
rect 79596 423098 79832 423334
rect 79596 419818 79832 420054
rect 79596 419498 79832 419734
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 79596 416218 79832 416454
rect 79596 415898 79832 416134
rect 64236 409018 64472 409254
rect 64236 408698 64472 408934
rect 64236 405418 64472 405654
rect 64236 405098 64472 405334
rect 64236 401818 64472 402054
rect 64236 401498 64472 401734
rect 64236 398218 64472 398454
rect 64236 397898 64472 398134
rect 79596 391018 79832 391254
rect 79596 390698 79832 390934
rect 79596 387418 79832 387654
rect 79596 387098 79832 387334
rect 79596 383818 79832 384054
rect 79596 383498 79832 383734
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 79596 380218 79832 380454
rect 79596 379898 79832 380134
rect 64236 373018 64472 373254
rect 64236 372698 64472 372934
rect 64236 369418 64472 369654
rect 64236 369098 64472 369334
rect 64236 365818 64472 366054
rect 64236 365498 64472 365734
rect 64236 362218 64472 362454
rect 64236 361898 64472 362134
rect 79596 355018 79832 355254
rect 79596 354698 79832 354934
rect 79596 351418 79832 351654
rect 79596 351098 79832 351334
rect 79596 347818 79832 348054
rect 79596 347498 79832 347734
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 79596 344218 79832 344454
rect 79596 343898 79832 344134
rect 64236 337018 64472 337254
rect 64236 336698 64472 336934
rect 64236 333418 64472 333654
rect 64236 333098 64472 333334
rect 64236 329818 64472 330054
rect 64236 329498 64472 329734
rect 64236 326218 64472 326454
rect 64236 325898 64472 326134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 282598 587212 282834 587298
rect 282598 587148 282684 587212
rect 282684 587148 282748 587212
rect 282748 587148 282834 587212
rect 282598 587062 282834 587148
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 386982 643018 387218 643254
rect 386982 642698 387218 642934
rect 386982 639418 387218 639654
rect 386982 639098 387218 639334
rect 386982 635818 387218 636054
rect 386982 635498 387218 635734
rect 386982 632218 387218 632454
rect 386982 631898 387218 632134
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 386536 625018 386772 625254
rect 386536 624698 386772 624934
rect 386536 621418 386772 621654
rect 386536 621098 386772 621334
rect 386536 617818 386772 618054
rect 386536 617498 386772 617734
rect 386536 614218 386772 614454
rect 386536 613898 386772 614134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 386982 607018 387218 607254
rect 386982 606698 387218 606934
rect 386982 603418 387218 603654
rect 386982 603098 387218 603334
rect 386982 599818 387218 600054
rect 386982 599498 387218 599734
rect 386982 596218 387218 596454
rect 386982 595898 387218 596134
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 386536 589018 386772 589254
rect 386536 588698 386772 588934
rect 387478 587212 387714 587298
rect 387478 587148 387564 587212
rect 387564 587148 387628 587212
rect 387628 587148 387714 587212
rect 387478 587062 387714 587148
rect 386536 585418 386772 585654
rect 386536 585098 386772 585334
rect 386536 581818 386772 582054
rect 386536 581498 386772 581734
rect 386536 578218 386772 578454
rect 386536 577898 386772 578134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 386982 571018 387218 571254
rect 386982 570698 387218 570934
rect 386982 567418 387218 567654
rect 386982 567098 387218 567334
rect 386982 563818 387218 564054
rect 386982 563498 387218 563734
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 310524 409018 310760 409254
rect 310524 408698 310760 408934
rect 310524 405418 310760 405654
rect 310524 405098 310760 405334
rect 310524 401818 310760 402054
rect 310524 401498 310760 401734
rect 310524 398218 310760 398454
rect 310524 397898 310760 398134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 310078 391018 310314 391254
rect 310078 390698 310314 390934
rect 310078 387418 310314 387654
rect 310078 387098 310314 387334
rect 310078 383818 310314 384054
rect 310078 383498 310314 383734
rect 310078 380218 310314 380454
rect 310078 379898 310314 380134
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 310524 373018 310760 373254
rect 310524 372698 310760 372934
rect 310524 369418 310760 369654
rect 310524 369098 310760 369334
rect 310524 365818 310760 366054
rect 310524 365498 310760 365734
rect 310524 362218 310760 362454
rect 310524 361898 310760 362134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 310078 355018 310314 355254
rect 310078 354698 310314 354934
rect 310078 351418 310314 351654
rect 310078 351098 310314 351334
rect 310078 347818 310314 348054
rect 310078 347498 310314 347734
rect 310078 344218 310314 344454
rect 310078 343898 310314 344134
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 310524 337018 310760 337254
rect 310524 336698 310760 336934
rect 310524 333418 310760 333654
rect 310524 333098 310760 333334
rect 310524 329818 310760 330054
rect 310524 329498 310760 329734
rect 310524 326218 310760 326454
rect 310524 325898 310760 326134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314236 293818 314472 294054
rect 314236 293498 314472 293734
rect 314236 290218 314472 290454
rect 314236 289898 314472 290134
rect 314236 265018 314472 265254
rect 314236 264698 314472 264934
rect 314236 261418 314472 261654
rect 314236 261098 314472 261334
rect 314236 257818 314472 258054
rect 314236 257498 314472 257734
rect 314236 254218 314472 254454
rect 314236 253898 314472 254134
rect 314236 229018 314472 229254
rect 314236 228698 314472 228934
rect 314236 225418 314472 225654
rect 314236 225098 314472 225334
rect 314236 221818 314472 222054
rect 314236 221498 314472 221734
rect 314236 218218 314472 218454
rect 314236 217898 314472 218134
rect 314236 193018 314472 193254
rect 314236 192698 314472 192934
rect 314236 189418 314472 189654
rect 314236 189098 314472 189334
rect 314236 185818 314472 186054
rect 314236 185498 314472 185734
rect 314236 182218 314472 182454
rect 314236 181898 314472 182134
rect 314236 157018 314472 157254
rect 314236 156698 314472 156934
rect 314236 153418 314472 153654
rect 314236 153098 314472 153334
rect 314236 149818 314472 150054
rect 314236 149498 314472 149734
rect 314236 146218 314472 146454
rect 314236 145898 314472 146134
rect 314236 121018 314472 121254
rect 314236 120698 314472 120934
rect 314236 117418 314472 117654
rect 314236 117098 314472 117334
rect 314236 113818 314472 114054
rect 314236 113498 314472 113734
rect 314236 110218 314472 110454
rect 314236 109898 314472 110134
rect 314236 85018 314472 85254
rect 314236 84698 314472 84934
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 516982 643018 517218 643254
rect 516982 642698 517218 642934
rect 516982 639418 517218 639654
rect 516982 639098 517218 639334
rect 516982 635818 517218 636054
rect 516982 635498 517218 635734
rect 516982 632218 517218 632454
rect 516982 631898 517218 632134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 516536 625018 516772 625254
rect 516536 624698 516772 624934
rect 516536 621418 516772 621654
rect 516536 621098 516772 621334
rect 516536 617818 516772 618054
rect 516536 617498 516772 617734
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 516536 614218 516772 614454
rect 516536 613898 516772 614134
rect 516982 607018 517218 607254
rect 516982 606698 517218 606934
rect 516982 603418 517218 603654
rect 516982 603098 517218 603334
rect 516982 599818 517218 600054
rect 516982 599498 517218 599734
rect 516982 596218 517218 596454
rect 516982 595898 517218 596134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 516536 589018 516772 589254
rect 516536 588698 516772 588934
rect 516536 585418 516772 585654
rect 516536 585098 516772 585334
rect 516536 581818 516772 582054
rect 516536 581498 516772 581734
rect 439918 579582 440154 579818
rect 518854 579582 519090 579818
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 516536 578218 516772 578454
rect 516536 577898 516772 578134
rect 516982 571018 517218 571254
rect 516982 570698 517218 570934
rect 516982 567418 517218 567654
rect 516982 567098 517218 567334
rect 516982 563818 517218 564054
rect 516982 563498 517218 563734
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 516536 405418 516772 405654
rect 516536 405098 516772 405334
rect 516536 401818 516772 402054
rect 516536 401498 516772 401734
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 516536 398218 516772 398454
rect 516536 397898 516772 398134
rect 516982 391018 517218 391254
rect 516982 390698 517218 390934
rect 516982 387418 517218 387654
rect 516982 387098 517218 387334
rect 516982 383818 517218 384054
rect 516982 383498 517218 383734
rect 516982 380218 517218 380454
rect 516982 379898 517218 380134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 516536 373018 516772 373254
rect 516536 372698 516772 372934
rect 516536 369418 516772 369654
rect 516536 369098 516772 369334
rect 516536 365818 516772 366054
rect 516536 365498 516772 365734
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 516536 362218 516772 362454
rect 516536 361898 516772 362134
rect 516982 355018 517218 355254
rect 516982 354698 517218 354934
rect 516982 351418 517218 351654
rect 516982 351098 517218 351334
rect 516982 347818 517218 348054
rect 516982 347498 517218 347734
rect 516982 344218 517218 344454
rect 516982 343898 517218 344134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 516536 337018 516772 337254
rect 516536 336698 516772 336934
rect 516536 333418 516772 333654
rect 516536 333098 516772 333334
rect 516536 329818 516772 330054
rect 516536 329498 516772 329734
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 516536 326218 516772 326454
rect 516536 325898 516772 326134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 329596 283018 329832 283254
rect 329596 282698 329832 282934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 329596 279418 329832 279654
rect 329596 279098 329832 279334
rect 329596 275818 329832 276054
rect 329596 275498 329832 275734
rect 329596 272218 329832 272454
rect 329596 271898 329832 272134
rect 329596 247018 329832 247254
rect 329596 246698 329832 246934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 329596 243418 329832 243654
rect 329596 243098 329832 243334
rect 329596 239818 329832 240054
rect 329596 239498 329832 239734
rect 329596 236218 329832 236454
rect 329596 235898 329832 236134
rect 329596 211018 329832 211254
rect 329596 210698 329832 210934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 329596 207418 329832 207654
rect 329596 207098 329832 207334
rect 329596 203818 329832 204054
rect 329596 203498 329832 203734
rect 329596 200218 329832 200454
rect 329596 199898 329832 200134
rect 329596 175018 329832 175254
rect 329596 174698 329832 174934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 329596 171418 329832 171654
rect 329596 171098 329832 171334
rect 329596 167818 329832 168054
rect 329596 167498 329832 167734
rect 329596 164218 329832 164454
rect 329596 163898 329832 164134
rect 329596 139018 329832 139254
rect 329596 138698 329832 138934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 329596 135418 329832 135654
rect 329596 135098 329832 135334
rect 329596 131818 329832 132054
rect 329596 131498 329832 131734
rect 329596 128218 329832 128454
rect 329596 127898 329832 128134
rect 329596 103018 329832 103254
rect 329596 102698 329832 102934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 329596 99418 329832 99654
rect 329596 99098 329832 99334
rect 329596 95818 329832 96054
rect 329596 95498 329832 95734
rect 329596 92218 329832 92454
rect 329596 91898 329832 92134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 292404 654076 293004 654078
rect 400404 654076 401004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 292586 654054
rect 292822 653818 400586 654054
rect 400822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 292586 653734
rect 292822 653498 400586 653734
rect 400822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 292404 653474 293004 653476
rect 400404 653474 401004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 288804 650476 289404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 288986 650454
rect 289222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 288986 650134
rect 289222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 288804 649874 289404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 136938 643276 137262 643278
rect 173604 643276 174204 643278
rect 266938 643276 267262 643278
rect 281604 643276 282204 643278
rect 386938 643276 387262 643278
rect 425604 643276 426204 643278
rect 516938 643276 517262 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 136982 643254
rect 137218 643018 173786 643254
rect 174022 643018 266982 643254
rect 267218 643018 281786 643254
rect 282022 643018 386982 643254
rect 387218 643018 425786 643254
rect 426022 643018 516982 643254
rect 517218 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 136982 642934
rect 137218 642698 173786 642934
rect 174022 642698 266982 642934
rect 267218 642698 281786 642934
rect 282022 642698 386982 642934
rect 387218 642698 425786 642934
rect 426022 642698 516982 642934
rect 517218 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 136938 642674 137262 642676
rect 173604 642674 174204 642676
rect 266938 642674 267262 642676
rect 281604 642674 282204 642676
rect 386938 642674 387262 642676
rect 425604 642674 426204 642676
rect 516938 642674 517262 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 136938 639676 137262 639678
rect 170004 639676 170604 639678
rect 266938 639676 267262 639678
rect 278004 639676 278604 639678
rect 386938 639676 387262 639678
rect 422004 639676 422604 639678
rect 516938 639676 517262 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 136982 639654
rect 137218 639418 170186 639654
rect 170422 639418 266982 639654
rect 267218 639418 278186 639654
rect 278422 639418 386982 639654
rect 387218 639418 422186 639654
rect 422422 639418 516982 639654
rect 517218 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 136982 639334
rect 137218 639098 170186 639334
rect 170422 639098 266982 639334
rect 267218 639098 278186 639334
rect 278422 639098 386982 639334
rect 387218 639098 422186 639334
rect 422422 639098 516982 639334
rect 517218 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 136938 639074 137262 639076
rect 170004 639074 170604 639076
rect 266938 639074 267262 639076
rect 278004 639074 278604 639076
rect 386938 639074 387262 639076
rect 422004 639074 422604 639076
rect 516938 639074 517262 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 136938 636076 137262 636078
rect 166404 636076 167004 636078
rect 266938 636076 267262 636078
rect 274404 636076 275004 636078
rect 386938 636076 387262 636078
rect 418404 636076 419004 636078
rect 516938 636076 517262 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 136982 636054
rect 137218 635818 166586 636054
rect 166822 635818 266982 636054
rect 267218 635818 274586 636054
rect 274822 635818 386982 636054
rect 387218 635818 418586 636054
rect 418822 635818 516982 636054
rect 517218 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 136982 635734
rect 137218 635498 166586 635734
rect 166822 635498 266982 635734
rect 267218 635498 274586 635734
rect 274822 635498 386982 635734
rect 387218 635498 418586 635734
rect 418822 635498 516982 635734
rect 517218 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 136938 635474 137262 635476
rect 166404 635474 167004 635476
rect 266938 635474 267262 635476
rect 274404 635474 275004 635476
rect 386938 635474 387262 635476
rect 418404 635474 419004 635476
rect 516938 635474 517262 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 136938 632476 137262 632478
rect 162804 632476 163404 632478
rect 266938 632476 267262 632478
rect 270804 632476 271404 632478
rect 386938 632476 387262 632478
rect 414804 632476 415404 632478
rect 516938 632476 517262 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 136982 632454
rect 137218 632218 162986 632454
rect 163222 632218 266982 632454
rect 267218 632218 270986 632454
rect 271222 632218 386982 632454
rect 387218 632218 414986 632454
rect 415222 632218 516982 632454
rect 517218 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 136982 632134
rect 137218 631898 162986 632134
rect 163222 631898 266982 632134
rect 267218 631898 270986 632134
rect 271222 631898 386982 632134
rect 387218 631898 414986 632134
rect 415222 631898 516982 632134
rect 517218 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 136938 631874 137262 631876
rect 162804 631874 163404 631876
rect 266938 631874 267262 631876
rect 270804 631874 271404 631876
rect 386938 631874 387262 631876
rect 414804 631874 415404 631876
rect 516938 631874 517262 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 136494 625276 136814 625278
rect 155604 625276 156204 625278
rect 266494 625276 266814 625278
rect 299604 625276 300204 625278
rect 386494 625276 386814 625278
rect 407604 625276 408204 625278
rect 516494 625276 516814 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 136536 625254
rect 136772 625018 155786 625254
rect 156022 625018 266536 625254
rect 266772 625018 299786 625254
rect 300022 625018 386536 625254
rect 386772 625018 407786 625254
rect 408022 625018 516536 625254
rect 516772 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 136536 624934
rect 136772 624698 155786 624934
rect 156022 624698 266536 624934
rect 266772 624698 299786 624934
rect 300022 624698 386536 624934
rect 386772 624698 407786 624934
rect 408022 624698 516536 624934
rect 516772 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 136494 624674 136814 624676
rect 155604 624674 156204 624676
rect 266494 624674 266814 624676
rect 299604 624674 300204 624676
rect 386494 624674 386814 624676
rect 407604 624674 408204 624676
rect 516494 624674 516814 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 136494 621676 136814 621678
rect 152004 621676 152604 621678
rect 266494 621676 266814 621678
rect 296004 621676 296604 621678
rect 386494 621676 386814 621678
rect 404004 621676 404604 621678
rect 516494 621676 516814 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 136536 621654
rect 136772 621418 152186 621654
rect 152422 621418 266536 621654
rect 266772 621418 296186 621654
rect 296422 621418 386536 621654
rect 386772 621418 404186 621654
rect 404422 621418 516536 621654
rect 516772 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 136536 621334
rect 136772 621098 152186 621334
rect 152422 621098 266536 621334
rect 266772 621098 296186 621334
rect 296422 621098 386536 621334
rect 386772 621098 404186 621334
rect 404422 621098 516536 621334
rect 516772 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 136494 621074 136814 621076
rect 152004 621074 152604 621076
rect 266494 621074 266814 621076
rect 296004 621074 296604 621076
rect 386494 621074 386814 621076
rect 404004 621074 404604 621076
rect 516494 621074 516814 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 136494 618076 136814 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 266494 618076 266814 618078
rect 292404 618076 293004 618078
rect 386494 618076 386814 618078
rect 400404 618076 401004 618078
rect 516494 618076 516814 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 136536 618054
rect 136772 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 266536 618054
rect 266772 617818 292586 618054
rect 292822 617818 386536 618054
rect 386772 617818 400586 618054
rect 400822 617818 516536 618054
rect 516772 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 136536 617734
rect 136772 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 266536 617734
rect 266772 617498 292586 617734
rect 292822 617498 386536 617734
rect 386772 617498 400586 617734
rect 400822 617498 516536 617734
rect 516772 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 136494 617474 136814 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 266494 617474 266814 617476
rect 292404 617474 293004 617476
rect 386494 617474 386814 617476
rect 400404 617474 401004 617476
rect 516494 617474 516814 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 136494 614476 136814 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 266494 614476 266814 614478
rect 288804 614476 289404 614478
rect 386494 614476 386814 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 516494 614476 516814 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 136536 614454
rect 136772 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 266536 614454
rect 266772 614218 288986 614454
rect 289222 614218 386536 614454
rect 386772 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 516536 614454
rect 516772 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 136536 614134
rect 136772 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 266536 614134
rect 266772 613898 288986 614134
rect 289222 613898 386536 614134
rect 386772 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 516536 614134
rect 516772 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 136494 613874 136814 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 266494 613874 266814 613876
rect 288804 613874 289404 613876
rect 386494 613874 386814 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 516494 613874 516814 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 136938 607276 137262 607278
rect 173604 607276 174204 607278
rect 266938 607276 267262 607278
rect 281604 607276 282204 607278
rect 386938 607276 387262 607278
rect 425604 607276 426204 607278
rect 516938 607276 517262 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 136982 607254
rect 137218 607018 173786 607254
rect 174022 607018 266982 607254
rect 267218 607018 281786 607254
rect 282022 607018 386982 607254
rect 387218 607018 425786 607254
rect 426022 607018 516982 607254
rect 517218 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 136982 606934
rect 137218 606698 173786 606934
rect 174022 606698 266982 606934
rect 267218 606698 281786 606934
rect 282022 606698 386982 606934
rect 387218 606698 425786 606934
rect 426022 606698 516982 606934
rect 517218 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 136938 606674 137262 606676
rect 173604 606674 174204 606676
rect 266938 606674 267262 606676
rect 281604 606674 282204 606676
rect 386938 606674 387262 606676
rect 425604 606674 426204 606676
rect 516938 606674 517262 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 136938 603676 137262 603678
rect 170004 603676 170604 603678
rect 266938 603676 267262 603678
rect 278004 603676 278604 603678
rect 386938 603676 387262 603678
rect 422004 603676 422604 603678
rect 516938 603676 517262 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 136982 603654
rect 137218 603418 170186 603654
rect 170422 603418 266982 603654
rect 267218 603418 278186 603654
rect 278422 603418 386982 603654
rect 387218 603418 422186 603654
rect 422422 603418 516982 603654
rect 517218 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 136982 603334
rect 137218 603098 170186 603334
rect 170422 603098 266982 603334
rect 267218 603098 278186 603334
rect 278422 603098 386982 603334
rect 387218 603098 422186 603334
rect 422422 603098 516982 603334
rect 517218 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 136938 603074 137262 603076
rect 170004 603074 170604 603076
rect 266938 603074 267262 603076
rect 278004 603074 278604 603076
rect 386938 603074 387262 603076
rect 422004 603074 422604 603076
rect 516938 603074 517262 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 136938 600076 137262 600078
rect 166404 600076 167004 600078
rect 266938 600076 267262 600078
rect 274404 600076 275004 600078
rect 386938 600076 387262 600078
rect 418404 600076 419004 600078
rect 516938 600076 517262 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 136982 600054
rect 137218 599818 166586 600054
rect 166822 599818 266982 600054
rect 267218 599818 274586 600054
rect 274822 599818 386982 600054
rect 387218 599818 418586 600054
rect 418822 599818 516982 600054
rect 517218 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 136982 599734
rect 137218 599498 166586 599734
rect 166822 599498 266982 599734
rect 267218 599498 274586 599734
rect 274822 599498 386982 599734
rect 387218 599498 418586 599734
rect 418822 599498 516982 599734
rect 517218 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 136938 599474 137262 599476
rect 166404 599474 167004 599476
rect 266938 599474 267262 599476
rect 274404 599474 275004 599476
rect 386938 599474 387262 599476
rect 418404 599474 419004 599476
rect 516938 599474 517262 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 136938 596476 137262 596478
rect 162804 596476 163404 596478
rect 266938 596476 267262 596478
rect 270804 596476 271404 596478
rect 386938 596476 387262 596478
rect 414804 596476 415404 596478
rect 516938 596476 517262 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 136982 596454
rect 137218 596218 162986 596454
rect 163222 596218 266982 596454
rect 267218 596218 270986 596454
rect 271222 596218 386982 596454
rect 387218 596218 414986 596454
rect 415222 596218 516982 596454
rect 517218 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 136982 596134
rect 137218 595898 162986 596134
rect 163222 595898 266982 596134
rect 267218 595898 270986 596134
rect 271222 595898 386982 596134
rect 387218 595898 414986 596134
rect 415222 595898 516982 596134
rect 517218 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 136938 595874 137262 595876
rect 162804 595874 163404 595876
rect 266938 595874 267262 595876
rect 270804 595874 271404 595876
rect 386938 595874 387262 595876
rect 414804 595874 415404 595876
rect 516938 595874 517262 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 136494 589276 136814 589278
rect 155604 589276 156204 589278
rect 266494 589276 266814 589278
rect 299604 589276 300204 589278
rect 386494 589276 386814 589278
rect 407604 589276 408204 589278
rect 516494 589276 516814 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 136536 589254
rect 136772 589018 155786 589254
rect 156022 589018 266536 589254
rect 266772 589018 299786 589254
rect 300022 589018 386536 589254
rect 386772 589018 407786 589254
rect 408022 589018 516536 589254
rect 516772 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 136536 588934
rect 136772 588698 155786 588934
rect 156022 588698 266536 588934
rect 266772 588698 299786 588934
rect 300022 588698 386536 588934
rect 386772 588698 407786 588934
rect 408022 588698 516536 588934
rect 516772 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 136494 588674 136814 588676
rect 155604 588674 156204 588676
rect 266494 588674 266814 588676
rect 299604 588674 300204 588676
rect 386494 588674 386814 588676
rect 407604 588674 408204 588676
rect 516494 588674 516814 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect 282556 587298 387756 587340
rect 282556 587062 282598 587298
rect 282834 587062 387478 587298
rect 387714 587062 387756 587298
rect 282556 587020 387756 587062
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 136494 585676 136814 585678
rect 152004 585676 152604 585678
rect 266494 585676 266814 585678
rect 296004 585676 296604 585678
rect 386494 585676 386814 585678
rect 404004 585676 404604 585678
rect 516494 585676 516814 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 136536 585654
rect 136772 585418 152186 585654
rect 152422 585418 266536 585654
rect 266772 585418 296186 585654
rect 296422 585418 386536 585654
rect 386772 585418 404186 585654
rect 404422 585418 516536 585654
rect 516772 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 136536 585334
rect 136772 585098 152186 585334
rect 152422 585098 266536 585334
rect 266772 585098 296186 585334
rect 296422 585098 386536 585334
rect 386772 585098 404186 585334
rect 404422 585098 516536 585334
rect 516772 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 136494 585074 136814 585076
rect 152004 585074 152604 585076
rect 266494 585074 266814 585076
rect 296004 585074 296604 585076
rect 386494 585074 386814 585076
rect 404004 585074 404604 585076
rect 516494 585074 516814 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 136494 582076 136814 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 266494 582076 266814 582078
rect 292404 582076 293004 582078
rect 386494 582076 386814 582078
rect 400404 582076 401004 582078
rect 516494 582076 516814 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 136536 582054
rect 136772 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 266536 582054
rect 266772 581818 292586 582054
rect 292822 581818 386536 582054
rect 386772 581818 400586 582054
rect 400822 581818 516536 582054
rect 516772 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 136536 581734
rect 136772 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 266536 581734
rect 266772 581498 292586 581734
rect 292822 581498 386536 581734
rect 386772 581498 400586 581734
rect 400822 581498 516536 581734
rect 516772 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 136494 581474 136814 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 266494 581474 266814 581476
rect 292404 581474 293004 581476
rect 386494 581474 386814 581476
rect 400404 581474 401004 581476
rect 516494 581474 516814 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect 439876 579818 519132 579860
rect 439876 579582 439918 579818
rect 440154 579582 518854 579818
rect 519090 579582 519132 579818
rect 439876 579540 519132 579582
rect 60468 579138 137700 579180
rect 60468 578902 60510 579138
rect 60746 578902 137422 579138
rect 137658 578902 137700 579138
rect 60468 578860 137700 578902
rect 190004 579138 269260 579180
rect 190004 578902 190046 579138
rect 190282 578902 268982 579138
rect 269218 578902 269260 579138
rect 190004 578860 269260 578902
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 136494 578476 136814 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 266494 578476 266814 578478
rect 288804 578476 289404 578478
rect 386494 578476 386814 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 516494 578476 516814 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 136536 578454
rect 136772 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 266536 578454
rect 266772 578218 288986 578454
rect 289222 578218 386536 578454
rect 386772 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 516536 578454
rect 516772 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 136536 578134
rect 136772 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 266536 578134
rect 266772 577898 288986 578134
rect 289222 577898 386536 578134
rect 386772 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 516536 578134
rect 516772 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 136494 577874 136814 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 266494 577874 266814 577876
rect 288804 577874 289404 577876
rect 386494 577874 386814 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 516494 577874 516814 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 136938 571276 137262 571278
rect 173604 571276 174204 571278
rect 266938 571276 267262 571278
rect 281604 571276 282204 571278
rect 386938 571276 387262 571278
rect 425604 571276 426204 571278
rect 516938 571276 517262 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 136982 571254
rect 137218 571018 173786 571254
rect 174022 571018 266982 571254
rect 267218 571018 281786 571254
rect 282022 571018 386982 571254
rect 387218 571018 425786 571254
rect 426022 571018 516982 571254
rect 517218 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 136982 570934
rect 137218 570698 173786 570934
rect 174022 570698 266982 570934
rect 267218 570698 281786 570934
rect 282022 570698 386982 570934
rect 387218 570698 425786 570934
rect 426022 570698 516982 570934
rect 517218 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 136938 570674 137262 570676
rect 173604 570674 174204 570676
rect 266938 570674 267262 570676
rect 281604 570674 282204 570676
rect 386938 570674 387262 570676
rect 425604 570674 426204 570676
rect 516938 570674 517262 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 136938 567676 137262 567678
rect 170004 567676 170604 567678
rect 266938 567676 267262 567678
rect 278004 567676 278604 567678
rect 386938 567676 387262 567678
rect 422004 567676 422604 567678
rect 516938 567676 517262 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 136982 567654
rect 137218 567418 170186 567654
rect 170422 567418 266982 567654
rect 267218 567418 278186 567654
rect 278422 567418 386982 567654
rect 387218 567418 422186 567654
rect 422422 567418 516982 567654
rect 517218 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 136982 567334
rect 137218 567098 170186 567334
rect 170422 567098 266982 567334
rect 267218 567098 278186 567334
rect 278422 567098 386982 567334
rect 387218 567098 422186 567334
rect 422422 567098 516982 567334
rect 517218 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 136938 567074 137262 567076
rect 170004 567074 170604 567076
rect 266938 567074 267262 567076
rect 278004 567074 278604 567076
rect 386938 567074 387262 567076
rect 422004 567074 422604 567076
rect 516938 567074 517262 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 136938 564076 137262 564078
rect 166404 564076 167004 564078
rect 266938 564076 267262 564078
rect 274404 564076 275004 564078
rect 386938 564076 387262 564078
rect 418404 564076 419004 564078
rect 516938 564076 517262 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 136982 564054
rect 137218 563818 166586 564054
rect 166822 563818 266982 564054
rect 267218 563818 274586 564054
rect 274822 563818 386982 564054
rect 387218 563818 418586 564054
rect 418822 563818 516982 564054
rect 517218 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 136982 563734
rect 137218 563498 166586 563734
rect 166822 563498 266982 563734
rect 267218 563498 274586 563734
rect 274822 563498 386982 563734
rect 387218 563498 418586 563734
rect 418822 563498 516982 563734
rect 517218 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 136938 563474 137262 563476
rect 166404 563474 167004 563476
rect 266938 563474 267262 563476
rect 274404 563474 275004 563476
rect 386938 563474 387262 563476
rect 418404 563474 419004 563476
rect 516938 563474 517262 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 162804 560476 163404 560478
rect 270804 560476 271404 560478
rect 414804 560476 415404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 162986 560454
rect 163222 560218 270986 560454
rect 271222 560218 414986 560454
rect 415222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 162986 560134
rect 163222 559898 270986 560134
rect 271222 559898 414986 560134
rect 415222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 162804 559874 163404 559876
rect 270804 559874 271404 559876
rect 414804 559874 415404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 79554 535276 79874 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 79596 535254
rect 79832 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 79596 534934
rect 79832 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 79554 534674 79874 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 79554 531676 79874 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 79596 531654
rect 79832 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 79596 531334
rect 79832 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 79554 531074 79874 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 79554 528076 79874 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 79596 528054
rect 79832 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 79596 527734
rect 79832 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 79554 527474 79874 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 79554 524476 79874 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 79596 524454
rect 79832 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 79596 524134
rect 79832 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 79554 523874 79874 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 64194 517276 64514 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 64236 517254
rect 64472 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 64236 516934
rect 64472 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 64194 516674 64514 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 64194 513676 64514 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 64236 513654
rect 64472 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 64236 513334
rect 64472 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 64194 513074 64514 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 64194 510076 64514 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 64236 510054
rect 64472 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 64236 509734
rect 64472 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 64194 509474 64514 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 64194 506476 64514 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 64236 506454
rect 64472 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 64236 506134
rect 64472 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 64194 505874 64514 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 79554 499276 79874 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 79596 499254
rect 79832 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 79596 498934
rect 79832 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 79554 498674 79874 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 79554 495676 79874 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 79596 495654
rect 79832 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 79596 495334
rect 79832 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 79554 495074 79874 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 79554 492076 79874 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 79596 492054
rect 79832 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 79596 491734
rect 79832 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 79554 491474 79874 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 79554 488476 79874 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 79596 488454
rect 79832 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 79596 488134
rect 79832 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 79554 487874 79874 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 64194 481276 64514 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 64236 481254
rect 64472 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 64236 480934
rect 64472 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 64194 480674 64514 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 64194 477676 64514 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 64236 477654
rect 64472 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 64236 477334
rect 64472 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 64194 477074 64514 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 64194 474076 64514 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 64236 474054
rect 64472 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 64236 473734
rect 64472 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 64194 473474 64514 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 64194 470476 64514 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 64236 470454
rect 64472 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 64236 470134
rect 64472 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 64194 469874 64514 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 79554 463276 79874 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 79596 463254
rect 79832 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 79596 462934
rect 79832 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 79554 462674 79874 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 79554 459676 79874 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 79596 459654
rect 79832 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 79596 459334
rect 79832 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 79554 459074 79874 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 79554 456076 79874 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 79596 456054
rect 79832 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 79596 455734
rect 79832 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 79554 455474 79874 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 79554 452476 79874 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 79596 452454
rect 79832 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 79596 452134
rect 79832 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 79554 451874 79874 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 64194 445276 64514 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 64236 445254
rect 64472 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 64236 444934
rect 64472 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 64194 444674 64514 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 64194 441676 64514 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 64236 441654
rect 64472 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 64236 441334
rect 64472 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 64194 441074 64514 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 64194 438076 64514 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 64236 438054
rect 64472 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 64236 437734
rect 64472 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 64194 437474 64514 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 64194 434476 64514 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 64236 434454
rect 64472 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 64236 434134
rect 64472 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 64194 433874 64514 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 79554 427276 79874 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 79596 427254
rect 79832 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 79596 426934
rect 79832 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 79554 426674 79874 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 79554 423676 79874 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 79596 423654
rect 79832 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 79596 423334
rect 79832 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 79554 423074 79874 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 79554 420076 79874 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 79596 420054
rect 79832 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 79596 419734
rect 79832 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 79554 419474 79874 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 79554 416476 79874 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 79596 416454
rect 79832 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 79596 416134
rect 79832 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 79554 415874 79874 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 64194 409276 64514 409278
rect 299604 409276 300204 409278
rect 310482 409276 310802 409278
rect 407604 409276 408204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 64236 409254
rect 64472 409018 299786 409254
rect 300022 409018 310524 409254
rect 310760 409018 407786 409254
rect 408022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 64236 408934
rect 64472 408698 299786 408934
rect 300022 408698 310524 408934
rect 310760 408698 407786 408934
rect 408022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 64194 408674 64514 408676
rect 299604 408674 300204 408676
rect 310482 408674 310802 408676
rect 407604 408674 408204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 64194 405676 64514 405678
rect 296004 405676 296604 405678
rect 310482 405676 310802 405678
rect 404004 405676 404604 405678
rect 516494 405676 516814 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 64236 405654
rect 64472 405418 296186 405654
rect 296422 405418 310524 405654
rect 310760 405418 404186 405654
rect 404422 405418 516536 405654
rect 516772 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 64236 405334
rect 64472 405098 296186 405334
rect 296422 405098 310524 405334
rect 310760 405098 404186 405334
rect 404422 405098 516536 405334
rect 516772 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 64194 405074 64514 405076
rect 296004 405074 296604 405076
rect 310482 405074 310802 405076
rect 404004 405074 404604 405076
rect 516494 405074 516814 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 64194 402076 64514 402078
rect 292404 402076 293004 402078
rect 310482 402076 310802 402078
rect 400404 402076 401004 402078
rect 516494 402076 516814 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 64236 402054
rect 64472 401818 292586 402054
rect 292822 401818 310524 402054
rect 310760 401818 400586 402054
rect 400822 401818 516536 402054
rect 516772 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 64236 401734
rect 64472 401498 292586 401734
rect 292822 401498 310524 401734
rect 310760 401498 400586 401734
rect 400822 401498 516536 401734
rect 516772 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 64194 401474 64514 401476
rect 292404 401474 293004 401476
rect 310482 401474 310802 401476
rect 400404 401474 401004 401476
rect 516494 401474 516814 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 64194 398476 64514 398478
rect 288804 398476 289404 398478
rect 310482 398476 310802 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 516494 398476 516814 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 64236 398454
rect 64472 398218 288986 398454
rect 289222 398218 310524 398454
rect 310760 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 516536 398454
rect 516772 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 64236 398134
rect 64472 397898 288986 398134
rect 289222 397898 310524 398134
rect 310760 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 516536 398134
rect 516772 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 64194 397874 64514 397876
rect 288804 397874 289404 397876
rect 310482 397874 310802 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 516494 397874 516814 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 79554 391276 79874 391278
rect 310034 391276 310358 391278
rect 425604 391276 426204 391278
rect 516938 391276 517262 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 79596 391254
rect 79832 391018 310078 391254
rect 310314 391018 425786 391254
rect 426022 391018 516982 391254
rect 517218 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 79596 390934
rect 79832 390698 310078 390934
rect 310314 390698 425786 390934
rect 426022 390698 516982 390934
rect 517218 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 79554 390674 79874 390676
rect 310034 390674 310358 390676
rect 425604 390674 426204 390676
rect 516938 390674 517262 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 79554 387676 79874 387678
rect 310034 387676 310358 387678
rect 422004 387676 422604 387678
rect 516938 387676 517262 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 79596 387654
rect 79832 387418 310078 387654
rect 310314 387418 422186 387654
rect 422422 387418 516982 387654
rect 517218 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 79596 387334
rect 79832 387098 310078 387334
rect 310314 387098 422186 387334
rect 422422 387098 516982 387334
rect 517218 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 79554 387074 79874 387076
rect 310034 387074 310358 387076
rect 422004 387074 422604 387076
rect 516938 387074 517262 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 79554 384076 79874 384078
rect 310034 384076 310358 384078
rect 418404 384076 419004 384078
rect 516938 384076 517262 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 79596 384054
rect 79832 383818 310078 384054
rect 310314 383818 418586 384054
rect 418822 383818 516982 384054
rect 517218 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 79596 383734
rect 79832 383498 310078 383734
rect 310314 383498 418586 383734
rect 418822 383498 516982 383734
rect 517218 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 79554 383474 79874 383476
rect 310034 383474 310358 383476
rect 418404 383474 419004 383476
rect 516938 383474 517262 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 79554 380476 79874 380478
rect 310034 380476 310358 380478
rect 414804 380476 415404 380478
rect 516938 380476 517262 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 79596 380454
rect 79832 380218 310078 380454
rect 310314 380218 414986 380454
rect 415222 380218 516982 380454
rect 517218 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 79596 380134
rect 79832 379898 310078 380134
rect 310314 379898 414986 380134
rect 415222 379898 516982 380134
rect 517218 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 79554 379874 79874 379876
rect 310034 379874 310358 379876
rect 414804 379874 415404 379876
rect 516938 379874 517262 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 64194 373276 64514 373278
rect 299604 373276 300204 373278
rect 310482 373276 310802 373278
rect 407604 373276 408204 373278
rect 516494 373276 516814 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 64236 373254
rect 64472 373018 299786 373254
rect 300022 373018 310524 373254
rect 310760 373018 407786 373254
rect 408022 373018 516536 373254
rect 516772 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 64236 372934
rect 64472 372698 299786 372934
rect 300022 372698 310524 372934
rect 310760 372698 407786 372934
rect 408022 372698 516536 372934
rect 516772 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 64194 372674 64514 372676
rect 299604 372674 300204 372676
rect 310482 372674 310802 372676
rect 407604 372674 408204 372676
rect 516494 372674 516814 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 64194 369676 64514 369678
rect 296004 369676 296604 369678
rect 310482 369676 310802 369678
rect 404004 369676 404604 369678
rect 516494 369676 516814 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 64236 369654
rect 64472 369418 296186 369654
rect 296422 369418 310524 369654
rect 310760 369418 404186 369654
rect 404422 369418 516536 369654
rect 516772 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 64236 369334
rect 64472 369098 296186 369334
rect 296422 369098 310524 369334
rect 310760 369098 404186 369334
rect 404422 369098 516536 369334
rect 516772 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 64194 369074 64514 369076
rect 296004 369074 296604 369076
rect 310482 369074 310802 369076
rect 404004 369074 404604 369076
rect 516494 369074 516814 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 64194 366076 64514 366078
rect 292404 366076 293004 366078
rect 310482 366076 310802 366078
rect 400404 366076 401004 366078
rect 516494 366076 516814 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 64236 366054
rect 64472 365818 292586 366054
rect 292822 365818 310524 366054
rect 310760 365818 400586 366054
rect 400822 365818 516536 366054
rect 516772 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 64236 365734
rect 64472 365498 292586 365734
rect 292822 365498 310524 365734
rect 310760 365498 400586 365734
rect 400822 365498 516536 365734
rect 516772 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 64194 365474 64514 365476
rect 292404 365474 293004 365476
rect 310482 365474 310802 365476
rect 400404 365474 401004 365476
rect 516494 365474 516814 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 64194 362476 64514 362478
rect 288804 362476 289404 362478
rect 310482 362476 310802 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 516494 362476 516814 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 64236 362454
rect 64472 362218 288986 362454
rect 289222 362218 310524 362454
rect 310760 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 516536 362454
rect 516772 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 64236 362134
rect 64472 361898 288986 362134
rect 289222 361898 310524 362134
rect 310760 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 516536 362134
rect 516772 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 64194 361874 64514 361876
rect 288804 361874 289404 361876
rect 310482 361874 310802 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 516494 361874 516814 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 79554 355276 79874 355278
rect 310034 355276 310358 355278
rect 425604 355276 426204 355278
rect 516938 355276 517262 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 79596 355254
rect 79832 355018 310078 355254
rect 310314 355018 425786 355254
rect 426022 355018 516982 355254
rect 517218 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 79596 354934
rect 79832 354698 310078 354934
rect 310314 354698 425786 354934
rect 426022 354698 516982 354934
rect 517218 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 79554 354674 79874 354676
rect 310034 354674 310358 354676
rect 425604 354674 426204 354676
rect 516938 354674 517262 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 79554 351676 79874 351678
rect 310034 351676 310358 351678
rect 422004 351676 422604 351678
rect 516938 351676 517262 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 79596 351654
rect 79832 351418 310078 351654
rect 310314 351418 422186 351654
rect 422422 351418 516982 351654
rect 517218 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 79596 351334
rect 79832 351098 310078 351334
rect 310314 351098 422186 351334
rect 422422 351098 516982 351334
rect 517218 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 79554 351074 79874 351076
rect 310034 351074 310358 351076
rect 422004 351074 422604 351076
rect 516938 351074 517262 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 79554 348076 79874 348078
rect 310034 348076 310358 348078
rect 418404 348076 419004 348078
rect 516938 348076 517262 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 79596 348054
rect 79832 347818 310078 348054
rect 310314 347818 418586 348054
rect 418822 347818 516982 348054
rect 517218 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 79596 347734
rect 79832 347498 310078 347734
rect 310314 347498 418586 347734
rect 418822 347498 516982 347734
rect 517218 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 79554 347474 79874 347476
rect 310034 347474 310358 347476
rect 418404 347474 419004 347476
rect 516938 347474 517262 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 79554 344476 79874 344478
rect 310034 344476 310358 344478
rect 414804 344476 415404 344478
rect 516938 344476 517262 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 79596 344454
rect 79832 344218 310078 344454
rect 310314 344218 414986 344454
rect 415222 344218 516982 344454
rect 517218 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 79596 344134
rect 79832 343898 310078 344134
rect 310314 343898 414986 344134
rect 415222 343898 516982 344134
rect 517218 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 79554 343874 79874 343876
rect 310034 343874 310358 343876
rect 414804 343874 415404 343876
rect 516938 343874 517262 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 64194 337276 64514 337278
rect 299604 337276 300204 337278
rect 310482 337276 310802 337278
rect 407604 337276 408204 337278
rect 516494 337276 516814 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 64236 337254
rect 64472 337018 299786 337254
rect 300022 337018 310524 337254
rect 310760 337018 407786 337254
rect 408022 337018 516536 337254
rect 516772 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 64236 336934
rect 64472 336698 299786 336934
rect 300022 336698 310524 336934
rect 310760 336698 407786 336934
rect 408022 336698 516536 336934
rect 516772 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 64194 336674 64514 336676
rect 299604 336674 300204 336676
rect 310482 336674 310802 336676
rect 407604 336674 408204 336676
rect 516494 336674 516814 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 64194 333676 64514 333678
rect 296004 333676 296604 333678
rect 310482 333676 310802 333678
rect 404004 333676 404604 333678
rect 516494 333676 516814 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 64236 333654
rect 64472 333418 296186 333654
rect 296422 333418 310524 333654
rect 310760 333418 404186 333654
rect 404422 333418 516536 333654
rect 516772 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 64236 333334
rect 64472 333098 296186 333334
rect 296422 333098 310524 333334
rect 310760 333098 404186 333334
rect 404422 333098 516536 333334
rect 516772 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 64194 333074 64514 333076
rect 296004 333074 296604 333076
rect 310482 333074 310802 333076
rect 404004 333074 404604 333076
rect 516494 333074 516814 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 64194 330076 64514 330078
rect 292404 330076 293004 330078
rect 310482 330076 310802 330078
rect 400404 330076 401004 330078
rect 516494 330076 516814 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 64236 330054
rect 64472 329818 292586 330054
rect 292822 329818 310524 330054
rect 310760 329818 400586 330054
rect 400822 329818 516536 330054
rect 516772 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 64236 329734
rect 64472 329498 292586 329734
rect 292822 329498 310524 329734
rect 310760 329498 400586 329734
rect 400822 329498 516536 329734
rect 516772 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 64194 329474 64514 329476
rect 292404 329474 293004 329476
rect 310482 329474 310802 329476
rect 400404 329474 401004 329476
rect 516494 329474 516814 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 64194 326476 64514 326478
rect 288804 326476 289404 326478
rect 310482 326476 310802 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 516494 326476 516814 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 64236 326454
rect 64472 326218 288986 326454
rect 289222 326218 310524 326454
rect 310760 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 516536 326454
rect 516772 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 64236 326134
rect 64472 325898 288986 326134
rect 289222 325898 310524 326134
rect 310760 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 516536 326134
rect 516772 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 64194 325874 64514 325876
rect 288804 325874 289404 325876
rect 310482 325874 310802 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 516494 325874 516814 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 425604 319276 426204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 425786 319254
rect 426022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 425786 318934
rect 426022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 425604 318674 426204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 314194 294076 314514 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 314236 294054
rect 314472 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 314236 293734
rect 314472 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 314194 293474 314514 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 314194 290476 314514 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 314236 290454
rect 314472 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 314236 290134
rect 314472 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 314194 289874 314514 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 329554 283276 329874 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 329596 283254
rect 329832 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 329596 282934
rect 329832 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 329554 282674 329874 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 329554 279676 329874 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 329596 279654
rect 329832 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 329596 279334
rect 329832 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 329554 279074 329874 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 329554 276076 329874 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 329596 276054
rect 329832 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 329596 275734
rect 329832 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 329554 275474 329874 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 329554 272476 329874 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 329596 272454
rect 329832 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 329596 272134
rect 329832 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 329554 271874 329874 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 314194 265276 314514 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 314236 265254
rect 314472 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 314236 264934
rect 314472 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 314194 264674 314514 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 314194 261676 314514 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 314236 261654
rect 314472 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 314236 261334
rect 314472 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 314194 261074 314514 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 314194 258076 314514 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 314236 258054
rect 314472 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 314236 257734
rect 314472 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 314194 257474 314514 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 314194 254476 314514 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 314236 254454
rect 314472 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 314236 254134
rect 314472 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 314194 253874 314514 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 329554 247276 329874 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 329596 247254
rect 329832 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 329596 246934
rect 329832 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 329554 246674 329874 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 329554 243676 329874 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 329596 243654
rect 329832 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 329596 243334
rect 329832 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 329554 243074 329874 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 329554 240076 329874 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 329596 240054
rect 329832 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 329596 239734
rect 329832 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 329554 239474 329874 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 329554 236476 329874 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 329596 236454
rect 329832 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 329596 236134
rect 329832 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 329554 235874 329874 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 314194 229276 314514 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 314236 229254
rect 314472 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 314236 228934
rect 314472 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 314194 228674 314514 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 314194 225676 314514 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 314236 225654
rect 314472 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 314236 225334
rect 314472 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 314194 225074 314514 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 314194 222076 314514 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 314236 222054
rect 314472 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 314236 221734
rect 314472 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 314194 221474 314514 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 314194 218476 314514 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 314236 218454
rect 314472 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 314236 218134
rect 314472 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 314194 217874 314514 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 329554 211276 329874 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 329596 211254
rect 329832 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 329596 210934
rect 329832 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 329554 210674 329874 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 329554 207676 329874 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 329596 207654
rect 329832 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 329596 207334
rect 329832 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 329554 207074 329874 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 329554 204076 329874 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 329596 204054
rect 329832 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 329596 203734
rect 329832 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 329554 203474 329874 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 329554 200476 329874 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 329596 200454
rect 329832 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 329596 200134
rect 329832 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 329554 199874 329874 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 314194 193276 314514 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 314236 193254
rect 314472 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 314236 192934
rect 314472 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 314194 192674 314514 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 314194 189676 314514 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 314236 189654
rect 314472 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 314236 189334
rect 314472 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 314194 189074 314514 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 314194 186076 314514 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 314236 186054
rect 314472 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 314236 185734
rect 314472 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 314194 185474 314514 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 314194 182476 314514 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 314236 182454
rect 314472 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 314236 182134
rect 314472 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 314194 181874 314514 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 329554 175276 329874 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 329596 175254
rect 329832 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 329596 174934
rect 329832 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 329554 174674 329874 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 329554 171676 329874 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 329596 171654
rect 329832 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 329596 171334
rect 329832 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 329554 171074 329874 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 329554 168076 329874 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 329596 168054
rect 329832 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 329596 167734
rect 329832 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 329554 167474 329874 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 329554 164476 329874 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 329596 164454
rect 329832 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 329596 164134
rect 329832 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 329554 163874 329874 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 314194 157276 314514 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 314236 157254
rect 314472 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 314236 156934
rect 314472 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 314194 156674 314514 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 314194 153676 314514 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 314236 153654
rect 314472 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 314236 153334
rect 314472 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 314194 153074 314514 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 314194 150076 314514 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 314236 150054
rect 314472 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 314236 149734
rect 314472 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 314194 149474 314514 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 314194 146476 314514 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 314236 146454
rect 314472 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 314236 146134
rect 314472 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 314194 145874 314514 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 329554 139276 329874 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 329596 139254
rect 329832 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 329596 138934
rect 329832 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 329554 138674 329874 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 329554 135676 329874 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 329596 135654
rect 329832 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 329596 135334
rect 329832 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 329554 135074 329874 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 329554 132076 329874 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 329596 132054
rect 329832 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 329596 131734
rect 329832 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 329554 131474 329874 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 329554 128476 329874 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 329596 128454
rect 329832 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 329596 128134
rect 329832 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 329554 127874 329874 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 314194 121276 314514 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 314236 121254
rect 314472 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 314236 120934
rect 314472 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 314194 120674 314514 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 314194 117676 314514 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 314236 117654
rect 314472 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 314236 117334
rect 314472 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 314194 117074 314514 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 314194 114076 314514 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 314236 114054
rect 314472 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 314236 113734
rect 314472 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 314194 113474 314514 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 314194 110476 314514 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 314236 110454
rect 314472 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 314236 110134
rect 314472 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 314194 109874 314514 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 329554 103276 329874 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 329596 103254
rect 329832 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 329596 102934
rect 329832 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 329554 102674 329874 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 329554 99676 329874 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 329596 99654
rect 329832 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 329596 99334
rect 329832 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 329554 99074 329874 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 329554 96076 329874 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 329596 96054
rect 329832 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 329596 95734
rect 329832 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 329554 95474 329874 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 329554 92476 329874 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 329596 92454
rect 329832 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 329596 92134
rect 329832 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 329554 91874 329874 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 314194 85276 314514 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 314236 85254
rect 314472 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 314236 84934
rect 314472 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 314194 84674 314514 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use sram_1rw1r_32_256_8_sky130  sram5
timestamp 1607837775
transform 1 0 440000 0 1 320000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram4
timestamp 1607837775
transform -1 0 387296 0 -1 411247
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram3
timestamp 1607837775
transform 1 0 440000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram2
timestamp 1607837775
transform 1 0 310000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram1
timestamp 1607837775
transform 1 0 190000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram0
timestamp 1607837775
transform 1 0 60000 0 1 560000
box 0 0 77296 91247
use hs32_core1  core1
timestamp 1607837775
transform 1 0 60000 0 1 320000
box 0 0 219986 220000
use hs32_core1  core0
timestamp 1607837775
transform 1 0 310000 0 1 80000
box 0 0 219986 220000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
