VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 2.400 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 2.400 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 2.400 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 2.400 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 2.400 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 2.400 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 2.400 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 2.400 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 2.400 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 2.400 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 2.400 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 2.400 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 2.400 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 2.400 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 2.400 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 17.920 633.350 17.980 ;
        RECT 676.270 17.920 676.590 17.980 ;
        RECT 633.030 17.780 676.590 17.920 ;
        RECT 633.030 17.720 633.350 17.780 ;
        RECT 676.270 17.720 676.590 17.780 ;
        RECT 678.110 17.920 678.430 17.980 ;
        RECT 814.730 17.920 815.050 17.980 ;
        RECT 678.110 17.780 815.050 17.920 ;
        RECT 678.110 17.720 678.430 17.780 ;
        RECT 814.730 17.720 815.050 17.780 ;
      LAYER via ;
        RECT 633.060 17.720 633.320 17.980 ;
        RECT 676.300 17.720 676.560 17.980 ;
        RECT 678.140 17.720 678.400 17.980 ;
        RECT 814.760 17.720 815.020 17.980 ;
      LAYER met2 ;
        RECT 815.680 1600.450 815.960 1604.000 ;
        RECT 814.820 1600.310 815.960 1600.450 ;
        RECT 633.060 17.690 633.320 18.010 ;
        RECT 676.290 17.835 676.570 18.205 ;
        RECT 678.130 17.835 678.410 18.205 ;
        RECT 814.820 18.010 814.960 1600.310 ;
        RECT 815.680 1600.000 815.960 1600.310 ;
        RECT 676.300 17.690 676.560 17.835 ;
        RECT 678.140 17.690 678.400 17.835 ;
        RECT 814.760 17.690 815.020 18.010 ;
        RECT 633.120 2.400 633.260 17.690 ;
        RECT 632.910 -4.800 633.470 2.400 ;
      LAYER via2 ;
        RECT 676.290 17.880 676.570 18.160 ;
        RECT 678.130 17.880 678.410 18.160 ;
      LAYER met3 ;
        RECT 676.265 18.170 676.595 18.185 ;
        RECT 678.105 18.170 678.435 18.185 ;
        RECT 676.265 17.870 678.435 18.170 ;
        RECT 676.265 17.855 676.595 17.870 ;
        RECT 678.105 17.855 678.435 17.870 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 796.790 1590.760 797.110 1590.820 ;
        RECT 830.370 1590.760 830.690 1590.820 ;
        RECT 796.790 1590.620 830.690 1590.760 ;
        RECT 796.790 1590.560 797.110 1590.620 ;
        RECT 830.370 1590.560 830.690 1590.620 ;
        RECT 650.970 15.540 651.290 15.600 ;
        RECT 796.790 15.540 797.110 15.600 ;
        RECT 650.970 15.400 797.110 15.540 ;
        RECT 650.970 15.340 651.290 15.400 ;
        RECT 796.790 15.340 797.110 15.400 ;
      LAYER via ;
        RECT 796.820 1590.560 797.080 1590.820 ;
        RECT 830.400 1590.560 830.660 1590.820 ;
        RECT 651.000 15.340 651.260 15.600 ;
        RECT 796.820 15.340 797.080 15.600 ;
      LAYER met2 ;
        RECT 830.400 1600.000 830.680 1604.000 ;
        RECT 830.460 1590.850 830.600 1600.000 ;
        RECT 796.820 1590.530 797.080 1590.850 ;
        RECT 830.400 1590.530 830.660 1590.850 ;
        RECT 796.880 15.630 797.020 1590.530 ;
        RECT 651.000 15.310 651.260 15.630 ;
        RECT 796.820 15.310 797.080 15.630 ;
        RECT 651.060 2.400 651.200 15.310 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 748.490 1591.780 748.810 1591.840 ;
        RECT 820.710 1591.780 821.030 1591.840 ;
        RECT 748.490 1591.640 821.030 1591.780 ;
        RECT 748.490 1591.580 748.810 1591.640 ;
        RECT 820.710 1591.580 821.030 1591.640 ;
        RECT 639.010 15.200 639.330 15.260 ;
        RECT 748.490 15.200 748.810 15.260 ;
        RECT 639.010 15.060 748.810 15.200 ;
        RECT 639.010 15.000 639.330 15.060 ;
        RECT 748.490 15.000 748.810 15.060 ;
      LAYER via ;
        RECT 748.520 1591.580 748.780 1591.840 ;
        RECT 820.740 1591.580 821.000 1591.840 ;
        RECT 639.040 15.000 639.300 15.260 ;
        RECT 748.520 15.000 748.780 15.260 ;
      LAYER met2 ;
        RECT 820.740 1600.000 821.020 1604.000 ;
        RECT 820.800 1591.870 820.940 1600.000 ;
        RECT 748.520 1591.550 748.780 1591.870 ;
        RECT 820.740 1591.550 821.000 1591.870 ;
        RECT 748.580 15.290 748.720 1591.550 ;
        RECT 639.040 14.970 639.300 15.290 ;
        RECT 748.520 14.970 748.780 15.290 ;
        RECT 639.100 2.400 639.240 14.970 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 17.240 657.270 17.300 ;
        RECT 676.270 17.240 676.590 17.300 ;
        RECT 656.950 17.100 676.590 17.240 ;
        RECT 656.950 17.040 657.270 17.100 ;
        RECT 676.270 17.040 676.590 17.100 ;
        RECT 678.110 17.240 678.430 17.300 ;
        RECT 835.430 17.240 835.750 17.300 ;
        RECT 678.110 17.100 835.750 17.240 ;
        RECT 678.110 17.040 678.430 17.100 ;
        RECT 835.430 17.040 835.750 17.100 ;
      LAYER via ;
        RECT 656.980 17.040 657.240 17.300 ;
        RECT 676.300 17.040 676.560 17.300 ;
        RECT 678.140 17.040 678.400 17.300 ;
        RECT 835.460 17.040 835.720 17.300 ;
      LAYER met2 ;
        RECT 835.000 1600.450 835.280 1604.000 ;
        RECT 835.000 1600.310 835.660 1600.450 ;
        RECT 835.000 1600.000 835.280 1600.310 ;
        RECT 835.520 17.330 835.660 1600.310 ;
        RECT 656.980 17.010 657.240 17.330 ;
        RECT 676.300 17.010 676.560 17.330 ;
        RECT 678.140 17.010 678.400 17.330 ;
        RECT 835.460 17.010 835.720 17.330 ;
        RECT 657.040 2.400 657.180 17.010 ;
        RECT 676.360 16.220 676.500 17.010 ;
        RECT 678.200 16.220 678.340 17.010 ;
        RECT 676.360 16.080 678.340 16.220 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 674.430 20.300 674.750 20.360 ;
        RECT 841.870 20.300 842.190 20.360 ;
        RECT 674.430 20.160 842.190 20.300 ;
        RECT 674.430 20.100 674.750 20.160 ;
        RECT 841.870 20.100 842.190 20.160 ;
      LAYER via ;
        RECT 674.460 20.100 674.720 20.360 ;
        RECT 841.900 20.100 842.160 20.360 ;
      LAYER met2 ;
        RECT 844.660 1600.450 844.940 1604.000 ;
        RECT 841.960 1600.310 844.940 1600.450 ;
        RECT 841.960 20.390 842.100 1600.310 ;
        RECT 844.660 1600.000 844.940 1600.310 ;
        RECT 674.460 20.070 674.720 20.390 ;
        RECT 841.900 20.070 842.160 20.390 ;
        RECT 674.520 2.400 674.660 20.070 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 676.805 18.785 677.895 18.955 ;
      LAYER mcon ;
        RECT 677.725 18.785 677.895 18.955 ;
      LAYER met1 ;
        RECT 644.990 18.940 645.310 19.000 ;
        RECT 676.745 18.940 677.035 18.985 ;
        RECT 644.990 18.800 677.035 18.940 ;
        RECT 644.990 18.740 645.310 18.800 ;
        RECT 676.745 18.755 677.035 18.800 ;
        RECT 677.665 18.940 677.955 18.985 ;
        RECT 821.170 18.940 821.490 19.000 ;
        RECT 677.665 18.800 821.490 18.940 ;
        RECT 677.665 18.755 677.955 18.800 ;
        RECT 821.170 18.740 821.490 18.800 ;
      LAYER via ;
        RECT 645.020 18.740 645.280 19.000 ;
        RECT 821.200 18.740 821.460 19.000 ;
      LAYER met2 ;
        RECT 825.340 1600.450 825.620 1604.000 ;
        RECT 821.260 1600.310 825.620 1600.450 ;
        RECT 821.260 19.030 821.400 1600.310 ;
        RECT 825.340 1600.000 825.620 1600.310 ;
        RECT 645.020 18.710 645.280 19.030 ;
        RECT 821.200 18.710 821.460 19.030 ;
        RECT 645.080 2.400 645.220 18.710 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.970 1590.080 835.290 1590.140 ;
        RECT 838.190 1590.080 838.510 1590.140 ;
        RECT 834.970 1589.940 838.510 1590.080 ;
        RECT 834.970 1589.880 835.290 1589.940 ;
        RECT 838.190 1589.880 838.510 1589.940 ;
        RECT 662.930 19.960 663.250 20.020 ;
        RECT 834.970 19.960 835.290 20.020 ;
        RECT 662.930 19.820 835.290 19.960 ;
        RECT 662.930 19.760 663.250 19.820 ;
        RECT 834.970 19.760 835.290 19.820 ;
      LAYER via ;
        RECT 835.000 1589.880 835.260 1590.140 ;
        RECT 838.220 1589.880 838.480 1590.140 ;
        RECT 662.960 19.760 663.220 20.020 ;
        RECT 835.000 19.760 835.260 20.020 ;
      LAYER met2 ;
        RECT 840.060 1600.450 840.340 1604.000 ;
        RECT 838.280 1600.310 840.340 1600.450 ;
        RECT 838.280 1590.170 838.420 1600.310 ;
        RECT 840.060 1600.000 840.340 1600.310 ;
        RECT 835.000 1589.850 835.260 1590.170 ;
        RECT 838.220 1589.850 838.480 1590.170 ;
        RECT 835.060 20.050 835.200 1589.850 ;
        RECT 662.960 19.730 663.220 20.050 ;
        RECT 835.000 19.730 835.260 20.050 ;
        RECT 663.020 2.400 663.160 19.730 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 327.205 1587.545 327.375 1590.435 ;
      LAYER mcon ;
        RECT 327.205 1590.265 327.375 1590.435 ;
      LAYER met1 ;
        RECT 321.610 2794.700 321.930 2794.760 ;
        RECT 972.050 2794.700 972.370 2794.760 ;
        RECT 1569.130 2794.700 1569.450 2794.760 ;
        RECT 1917.810 2794.700 1918.130 2794.760 ;
        RECT 321.610 2794.560 1918.130 2794.700 ;
        RECT 321.610 2794.500 321.930 2794.560 ;
        RECT 972.050 2794.500 972.370 2794.560 ;
        RECT 1569.130 2794.500 1569.450 2794.560 ;
        RECT 1917.810 2794.500 1918.130 2794.560 ;
        RECT 1917.810 2791.300 1918.130 2791.360 ;
        RECT 2215.430 2791.300 2215.750 2791.360 ;
        RECT 1917.810 2791.160 2215.750 2791.300 ;
        RECT 1917.810 2791.100 1918.130 2791.160 ;
        RECT 2215.430 2791.100 2215.750 2791.160 ;
        RECT 1917.810 2066.420 1918.130 2066.480 ;
        RECT 2024.990 2066.420 2025.310 2066.480 ;
        RECT 1917.810 2066.280 2025.310 2066.420 ;
        RECT 1917.810 2066.220 1918.130 2066.280 ;
        RECT 2024.990 2066.220 2025.310 2066.280 ;
        RECT 2024.990 2063.360 2025.310 2063.420 ;
        RECT 2566.870 2063.360 2567.190 2063.420 ;
        RECT 2024.990 2063.220 2567.190 2063.360 ;
        RECT 2024.990 2063.160 2025.310 2063.220 ;
        RECT 2566.870 2063.160 2567.190 2063.220 ;
        RECT 1566.370 1593.820 1566.690 1593.880 ;
        RECT 2024.990 1593.820 2025.310 1593.880 ;
        RECT 2215.430 1593.820 2215.750 1593.880 ;
        RECT 1566.370 1593.680 2215.750 1593.820 ;
        RECT 1566.370 1593.620 1566.690 1593.680 ;
        RECT 2024.990 1593.620 2025.310 1593.680 ;
        RECT 2215.430 1593.620 2215.750 1593.680 ;
        RECT 327.145 1590.420 327.435 1590.465 ;
        RECT 1566.370 1590.420 1566.690 1590.480 ;
        RECT 327.145 1590.280 1566.690 1590.420 ;
        RECT 327.145 1590.235 327.435 1590.280 ;
        RECT 1566.370 1590.220 1566.690 1590.280 ;
        RECT 327.145 1587.700 327.435 1587.745 ;
        RECT 313.880 1587.560 327.435 1587.700 ;
        RECT 299.990 1587.360 300.310 1587.420 ;
        RECT 313.880 1587.360 314.020 1587.560 ;
        RECT 327.145 1587.515 327.435 1587.560 ;
        RECT 299.990 1587.220 314.020 1587.360 ;
        RECT 299.990 1587.160 300.310 1587.220 ;
        RECT 2.830 24.040 3.150 24.100 ;
        RECT 299.990 24.040 300.310 24.100 ;
        RECT 2.830 23.900 300.310 24.040 ;
        RECT 2.830 23.840 3.150 23.900 ;
        RECT 299.990 23.840 300.310 23.900 ;
      LAYER via ;
        RECT 321.640 2794.500 321.900 2794.760 ;
        RECT 972.080 2794.500 972.340 2794.760 ;
        RECT 1569.160 2794.500 1569.420 2794.760 ;
        RECT 1917.840 2794.500 1918.100 2794.760 ;
        RECT 1917.840 2791.100 1918.100 2791.360 ;
        RECT 2215.460 2791.100 2215.720 2791.360 ;
        RECT 1917.840 2066.220 1918.100 2066.480 ;
        RECT 2025.020 2066.220 2025.280 2066.480 ;
        RECT 2025.020 2063.160 2025.280 2063.420 ;
        RECT 2566.900 2063.160 2567.160 2063.420 ;
        RECT 1566.400 1593.620 1566.660 1593.880 ;
        RECT 2025.020 1593.620 2025.280 1593.880 ;
        RECT 2215.460 1593.620 2215.720 1593.880 ;
        RECT 1566.400 1590.220 1566.660 1590.480 ;
        RECT 300.020 1587.160 300.280 1587.420 ;
        RECT 2.860 23.840 3.120 24.100 ;
        RECT 300.020 23.840 300.280 24.100 ;
      LAYER met2 ;
        RECT 321.640 2794.645 321.900 2794.790 ;
        RECT 972.080 2794.645 972.340 2794.790 ;
        RECT 1569.160 2794.645 1569.420 2794.790 ;
        RECT 321.630 2794.275 321.910 2794.645 ;
        RECT 972.070 2794.275 972.350 2794.645 ;
        RECT 1569.150 2794.275 1569.430 2794.645 ;
        RECT 1917.840 2794.470 1918.100 2794.790 ;
        RECT 1917.900 2791.390 1918.040 2794.470 ;
        RECT 2215.450 2794.275 2215.730 2794.645 ;
        RECT 2215.520 2791.390 2215.660 2794.275 ;
        RECT 1917.840 2791.070 1918.100 2791.390 ;
        RECT 2215.460 2791.070 2215.720 2791.390 ;
        RECT 1917.900 2066.510 1918.040 2791.070 ;
        RECT 1917.840 2066.365 1918.100 2066.510 ;
        RECT 1917.830 2065.995 1918.110 2066.365 ;
        RECT 2025.020 2066.190 2025.280 2066.510 ;
        RECT 2025.080 2063.450 2025.220 2066.190 ;
        RECT 2025.020 2063.130 2025.280 2063.450 ;
        RECT 2566.890 2063.275 2567.170 2063.645 ;
        RECT 2566.900 2063.130 2567.160 2063.275 ;
        RECT 302.320 1600.450 302.600 1604.000 ;
        RECT 300.080 1600.310 302.600 1600.450 ;
        RECT 300.080 1587.450 300.220 1600.310 ;
        RECT 302.320 1600.000 302.600 1600.310 ;
        RECT 2025.080 1593.910 2025.220 2063.130 ;
        RECT 1566.400 1593.765 1566.660 1593.910 ;
        RECT 1566.390 1593.395 1566.670 1593.765 ;
        RECT 2025.020 1593.590 2025.280 1593.910 ;
        RECT 2215.460 1593.765 2215.720 1593.910 ;
        RECT 2215.450 1593.395 2215.730 1593.765 ;
        RECT 1566.460 1590.510 1566.600 1593.395 ;
        RECT 1566.400 1590.190 1566.660 1590.510 ;
        RECT 300.020 1587.130 300.280 1587.450 ;
        RECT 300.080 24.130 300.220 1587.130 ;
        RECT 2.860 23.810 3.120 24.130 ;
        RECT 300.020 23.810 300.280 24.130 ;
        RECT 2.920 2.400 3.060 23.810 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 321.630 2794.320 321.910 2794.600 ;
        RECT 972.070 2794.320 972.350 2794.600 ;
        RECT 1569.150 2794.320 1569.430 2794.600 ;
        RECT 2215.450 2794.320 2215.730 2794.600 ;
        RECT 1917.830 2066.040 1918.110 2066.320 ;
        RECT 2566.890 2063.320 2567.170 2063.600 ;
        RECT 1566.390 1593.440 1566.670 1593.720 ;
        RECT 2215.450 1593.440 2215.730 1593.720 ;
      LAYER met3 ;
        RECT 321.605 2794.620 321.935 2794.625 ;
        RECT 972.045 2794.620 972.375 2794.625 ;
        RECT 1569.125 2794.620 1569.455 2794.625 ;
        RECT 321.350 2794.610 321.935 2794.620 ;
        RECT 971.790 2794.610 972.375 2794.620 ;
        RECT 1568.870 2794.610 1569.455 2794.620 ;
        RECT 321.150 2794.310 321.935 2794.610 ;
        RECT 971.590 2794.310 972.375 2794.610 ;
        RECT 1568.670 2794.310 1569.455 2794.610 ;
        RECT 321.350 2794.300 321.935 2794.310 ;
        RECT 971.790 2794.300 972.375 2794.310 ;
        RECT 1568.870 2794.300 1569.455 2794.310 ;
        RECT 321.605 2794.295 321.935 2794.300 ;
        RECT 972.045 2794.295 972.375 2794.300 ;
        RECT 1569.125 2794.295 1569.455 2794.300 ;
        RECT 2215.425 2794.620 2215.755 2794.625 ;
        RECT 2215.425 2794.610 2216.010 2794.620 ;
        RECT 2215.425 2794.310 2216.210 2794.610 ;
        RECT 2215.425 2794.300 2216.010 2794.310 ;
        RECT 2215.425 2794.295 2215.755 2794.300 ;
        RECT 1917.805 2066.340 1918.135 2066.345 ;
        RECT 1917.550 2066.330 1918.135 2066.340 ;
        RECT 1917.350 2066.030 1918.135 2066.330 ;
        RECT 1917.550 2066.020 1918.135 2066.030 ;
        RECT 1917.805 2066.015 1918.135 2066.020 ;
        RECT 2566.865 2063.620 2567.195 2063.625 ;
        RECT 2566.865 2063.610 2567.450 2063.620 ;
        RECT 2566.640 2063.310 2567.450 2063.610 ;
        RECT 2566.865 2063.300 2567.450 2063.310 ;
        RECT 2566.865 2063.295 2567.195 2063.300 ;
        RECT 1566.365 1593.730 1566.695 1593.745 ;
        RECT 2215.425 1593.740 2215.755 1593.745 ;
        RECT 1567.030 1593.730 1567.410 1593.740 ;
        RECT 1566.365 1593.430 1567.410 1593.730 ;
        RECT 1566.365 1593.415 1566.695 1593.430 ;
        RECT 1567.030 1593.420 1567.410 1593.430 ;
        RECT 2215.425 1593.730 2216.010 1593.740 ;
        RECT 2215.425 1593.430 2216.210 1593.730 ;
        RECT 2215.425 1593.420 2216.010 1593.430 ;
        RECT 2215.425 1593.415 2215.755 1593.420 ;
      LAYER via3 ;
        RECT 321.380 2794.300 321.700 2794.620 ;
        RECT 971.820 2794.300 972.140 2794.620 ;
        RECT 1568.900 2794.300 1569.220 2794.620 ;
        RECT 2215.660 2794.300 2215.980 2794.620 ;
        RECT 1917.580 2066.020 1917.900 2066.340 ;
        RECT 2567.100 2063.300 2567.420 2063.620 ;
        RECT 1567.060 1593.420 1567.380 1593.740 ;
        RECT 2215.660 1593.420 2215.980 1593.740 ;
      LAYER met4 ;
        RECT 319.015 2801.750 319.315 2804.600 ;
        RECT 969.015 2801.750 969.315 2804.600 ;
        RECT 1569.015 2801.750 1569.315 2804.600 ;
        RECT 2219.015 2801.750 2219.315 2804.600 ;
        RECT 319.015 2801.450 321.690 2801.750 ;
        RECT 319.015 2800.000 319.315 2801.450 ;
        RECT 321.390 2794.625 321.690 2801.450 ;
        RECT 969.015 2801.450 972.130 2801.750 ;
        RECT 969.015 2800.000 969.315 2801.450 ;
        RECT 971.830 2794.625 972.130 2801.450 ;
        RECT 1568.910 2800.000 1569.315 2801.750 ;
        RECT 2215.670 2801.450 2219.315 2801.750 ;
        RECT 1568.910 2794.625 1569.210 2800.000 ;
        RECT 2215.670 2794.625 2215.970 2801.450 ;
        RECT 2219.015 2800.000 2219.315 2801.450 ;
        RECT 321.375 2794.295 321.705 2794.625 ;
        RECT 971.815 2794.295 972.145 2794.625 ;
        RECT 1568.895 2794.295 1569.225 2794.625 ;
        RECT 2215.655 2794.295 2215.985 2794.625 ;
        RECT 1917.575 2066.015 1917.905 2066.345 ;
        RECT 1917.590 2058.850 1917.890 2066.015 ;
        RECT 2567.095 2063.295 2567.425 2063.625 ;
        RECT 1917.165 2058.550 1917.890 2058.850 ;
        RECT 1917.165 2051.635 1917.465 2058.550 ;
        RECT 2567.110 2055.450 2567.410 2063.295 ;
        RECT 2567.865 2055.450 2568.165 2056.235 ;
        RECT 2567.110 2055.150 2568.165 2055.450 ;
        RECT 2567.865 2051.635 2568.165 2055.150 ;
        RECT 1568.315 1601.550 1568.615 1604.600 ;
        RECT 2219.015 1601.550 2219.315 1604.600 ;
        RECT 1567.070 1601.250 1568.615 1601.550 ;
        RECT 1567.070 1593.745 1567.370 1601.250 ;
        RECT 1568.315 1600.000 1568.615 1601.250 ;
        RECT 2215.670 1601.250 2219.315 1601.550 ;
        RECT 2215.670 1593.745 2215.970 1601.250 ;
        RECT 2219.015 1600.000 2219.315 1601.250 ;
        RECT 1567.055 1593.415 1567.385 1593.745 ;
        RECT 2215.655 1593.415 2215.985 1593.745 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 24.720 8.670 24.780 ;
        RECT 303.670 24.720 303.990 24.780 ;
        RECT 8.350 24.580 303.990 24.720 ;
        RECT 8.350 24.520 8.670 24.580 ;
        RECT 303.670 24.520 303.990 24.580 ;
      LAYER via ;
        RECT 8.380 24.520 8.640 24.780 ;
        RECT 303.700 24.520 303.960 24.780 ;
      LAYER met2 ;
        RECT 306.920 1600.450 307.200 1604.000 ;
        RECT 303.760 1600.310 307.200 1600.450 ;
        RECT 303.760 24.810 303.900 1600.310 ;
        RECT 306.920 1600.000 307.200 1600.310 ;
        RECT 8.380 24.490 8.640 24.810 ;
        RECT 303.700 24.490 303.960 24.810 ;
        RECT 8.440 2.400 8.580 24.490 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 24.380 14.650 24.440 ;
        RECT 311.030 24.380 311.350 24.440 ;
        RECT 14.330 24.240 311.350 24.380 ;
        RECT 14.330 24.180 14.650 24.240 ;
        RECT 311.030 24.180 311.350 24.240 ;
      LAYER via ;
        RECT 14.360 24.180 14.620 24.440 ;
        RECT 311.060 24.180 311.320 24.440 ;
      LAYER met2 ;
        RECT 311.980 1600.450 312.260 1604.000 ;
        RECT 311.120 1600.310 312.260 1600.450 ;
        RECT 311.120 24.470 311.260 1600.310 ;
        RECT 311.980 1600.000 312.260 1600.310 ;
        RECT 14.360 24.150 14.620 24.470 ;
        RECT 311.060 24.150 311.320 24.470 ;
        RECT 14.420 2.400 14.560 24.150 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 331.730 25.060 332.050 25.120 ;
        RECT 38.250 24.920 332.050 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 331.730 24.860 332.050 24.920 ;
      LAYER via ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 331.760 24.860 332.020 25.120 ;
      LAYER met2 ;
        RECT 331.300 1600.450 331.580 1604.000 ;
        RECT 331.300 1600.310 331.960 1600.450 ;
        RECT 331.300 1600.000 331.580 1600.310 ;
        RECT 331.820 25.150 331.960 1600.310 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 331.760 24.830 332.020 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 490.965 1256.045 491.135 1304.155 ;
        RECT 490.045 386.325 490.215 434.775 ;
        RECT 490.965 241.485 491.135 289.595 ;
        RECT 490.965 144.925 491.135 193.035 ;
        RECT 491.425 48.365 491.595 96.475 ;
      LAYER mcon ;
        RECT 490.965 1303.985 491.135 1304.155 ;
        RECT 490.045 434.605 490.215 434.775 ;
        RECT 490.965 289.425 491.135 289.595 ;
        RECT 490.965 192.865 491.135 193.035 ;
        RECT 491.425 96.305 491.595 96.475 ;
      LAYER met1 ;
        RECT 490.430 1511.200 490.750 1511.260 ;
        RECT 491.350 1511.200 491.670 1511.260 ;
        RECT 490.430 1511.060 491.670 1511.200 ;
        RECT 490.430 1511.000 490.750 1511.060 ;
        RECT 491.350 1511.000 491.670 1511.060 ;
        RECT 490.890 1442.180 491.210 1442.240 ;
        RECT 491.810 1442.180 492.130 1442.240 ;
        RECT 490.890 1442.040 492.130 1442.180 ;
        RECT 490.890 1441.980 491.210 1442.040 ;
        RECT 491.810 1441.980 492.130 1442.040 ;
        RECT 491.810 1345.620 492.130 1345.680 ;
        RECT 492.270 1345.620 492.590 1345.680 ;
        RECT 491.810 1345.480 492.590 1345.620 ;
        RECT 491.810 1345.420 492.130 1345.480 ;
        RECT 492.270 1345.420 492.590 1345.480 ;
        RECT 490.890 1304.140 491.210 1304.200 ;
        RECT 490.695 1304.000 491.210 1304.140 ;
        RECT 490.890 1303.940 491.210 1304.000 ;
        RECT 490.905 1256.200 491.195 1256.245 ;
        RECT 491.350 1256.200 491.670 1256.260 ;
        RECT 490.905 1256.060 491.670 1256.200 ;
        RECT 490.905 1256.015 491.195 1256.060 ;
        RECT 491.350 1256.000 491.670 1256.060 ;
        RECT 489.970 1159.300 490.290 1159.360 ;
        RECT 491.350 1159.300 491.670 1159.360 ;
        RECT 489.970 1159.160 491.670 1159.300 ;
        RECT 489.970 1159.100 490.290 1159.160 ;
        RECT 491.350 1159.100 491.670 1159.160 ;
        RECT 489.970 1062.740 490.290 1062.800 ;
        RECT 491.350 1062.740 491.670 1062.800 ;
        RECT 489.970 1062.600 491.670 1062.740 ;
        RECT 489.970 1062.540 490.290 1062.600 ;
        RECT 491.350 1062.540 491.670 1062.600 ;
        RECT 489.970 966.180 490.290 966.240 ;
        RECT 491.350 966.180 491.670 966.240 ;
        RECT 489.970 966.040 491.670 966.180 ;
        RECT 489.970 965.980 490.290 966.040 ;
        RECT 491.350 965.980 491.670 966.040 ;
        RECT 489.970 869.620 490.290 869.680 ;
        RECT 491.350 869.620 491.670 869.680 ;
        RECT 489.970 869.480 491.670 869.620 ;
        RECT 489.970 869.420 490.290 869.480 ;
        RECT 491.350 869.420 491.670 869.480 ;
        RECT 489.970 821.000 490.290 821.060 ;
        RECT 490.890 821.000 491.210 821.060 ;
        RECT 489.970 820.860 491.210 821.000 ;
        RECT 489.970 820.800 490.290 820.860 ;
        RECT 490.890 820.800 491.210 820.860 ;
        RECT 489.985 434.760 490.275 434.805 ;
        RECT 490.430 434.760 490.750 434.820 ;
        RECT 489.985 434.620 490.750 434.760 ;
        RECT 489.985 434.575 490.275 434.620 ;
        RECT 490.430 434.560 490.750 434.620 ;
        RECT 489.970 386.480 490.290 386.540 ;
        RECT 489.775 386.340 490.290 386.480 ;
        RECT 489.970 386.280 490.290 386.340 ;
        RECT 489.970 338.340 490.290 338.600 ;
        RECT 490.060 338.200 490.200 338.340 ;
        RECT 490.430 338.200 490.750 338.260 ;
        RECT 490.060 338.060 490.750 338.200 ;
        RECT 490.430 338.000 490.750 338.060 ;
        RECT 490.430 303.520 490.750 303.580 ;
        RECT 491.350 303.520 491.670 303.580 ;
        RECT 490.430 303.380 491.670 303.520 ;
        RECT 490.430 303.320 490.750 303.380 ;
        RECT 491.350 303.320 491.670 303.380 ;
        RECT 490.905 289.580 491.195 289.625 ;
        RECT 491.350 289.580 491.670 289.640 ;
        RECT 490.905 289.440 491.670 289.580 ;
        RECT 490.905 289.395 491.195 289.440 ;
        RECT 491.350 289.380 491.670 289.440 ;
        RECT 490.890 241.640 491.210 241.700 ;
        RECT 490.695 241.500 491.210 241.640 ;
        RECT 490.890 241.440 491.210 241.500 ;
        RECT 490.430 206.960 490.750 207.020 ;
        RECT 491.350 206.960 491.670 207.020 ;
        RECT 490.430 206.820 491.670 206.960 ;
        RECT 490.430 206.760 490.750 206.820 ;
        RECT 491.350 206.760 491.670 206.820 ;
        RECT 490.905 193.020 491.195 193.065 ;
        RECT 491.350 193.020 491.670 193.080 ;
        RECT 490.905 192.880 491.670 193.020 ;
        RECT 490.905 192.835 491.195 192.880 ;
        RECT 491.350 192.820 491.670 192.880 ;
        RECT 490.890 145.080 491.210 145.140 ;
        RECT 490.695 144.940 491.210 145.080 ;
        RECT 490.890 144.880 491.210 144.940 ;
        RECT 490.430 110.400 490.750 110.460 ;
        RECT 491.350 110.400 491.670 110.460 ;
        RECT 490.430 110.260 491.670 110.400 ;
        RECT 490.430 110.200 490.750 110.260 ;
        RECT 491.350 110.200 491.670 110.260 ;
        RECT 491.350 96.460 491.670 96.520 ;
        RECT 491.155 96.320 491.670 96.460 ;
        RECT 491.350 96.260 491.670 96.320 ;
        RECT 491.350 48.520 491.670 48.580 ;
        RECT 491.155 48.380 491.670 48.520 ;
        RECT 491.350 48.320 491.670 48.380 ;
        RECT 240.650 23.700 240.970 23.760 ;
        RECT 491.350 23.700 491.670 23.760 ;
        RECT 240.650 23.560 491.670 23.700 ;
        RECT 240.650 23.500 240.970 23.560 ;
        RECT 491.350 23.500 491.670 23.560 ;
      LAYER via ;
        RECT 490.460 1511.000 490.720 1511.260 ;
        RECT 491.380 1511.000 491.640 1511.260 ;
        RECT 490.920 1441.980 491.180 1442.240 ;
        RECT 491.840 1441.980 492.100 1442.240 ;
        RECT 491.840 1345.420 492.100 1345.680 ;
        RECT 492.300 1345.420 492.560 1345.680 ;
        RECT 490.920 1303.940 491.180 1304.200 ;
        RECT 491.380 1256.000 491.640 1256.260 ;
        RECT 490.000 1159.100 490.260 1159.360 ;
        RECT 491.380 1159.100 491.640 1159.360 ;
        RECT 490.000 1062.540 490.260 1062.800 ;
        RECT 491.380 1062.540 491.640 1062.800 ;
        RECT 490.000 965.980 490.260 966.240 ;
        RECT 491.380 965.980 491.640 966.240 ;
        RECT 490.000 869.420 490.260 869.680 ;
        RECT 491.380 869.420 491.640 869.680 ;
        RECT 490.000 820.800 490.260 821.060 ;
        RECT 490.920 820.800 491.180 821.060 ;
        RECT 490.460 434.560 490.720 434.820 ;
        RECT 490.000 386.280 490.260 386.540 ;
        RECT 490.000 338.340 490.260 338.600 ;
        RECT 490.460 338.000 490.720 338.260 ;
        RECT 490.460 303.320 490.720 303.580 ;
        RECT 491.380 303.320 491.640 303.580 ;
        RECT 491.380 289.380 491.640 289.640 ;
        RECT 490.920 241.440 491.180 241.700 ;
        RECT 490.460 206.760 490.720 207.020 ;
        RECT 491.380 206.760 491.640 207.020 ;
        RECT 491.380 192.820 491.640 193.080 ;
        RECT 490.920 144.880 491.180 145.140 ;
        RECT 490.460 110.200 490.720 110.460 ;
        RECT 491.380 110.200 491.640 110.460 ;
        RECT 491.380 96.260 491.640 96.520 ;
        RECT 491.380 48.320 491.640 48.580 ;
        RECT 240.680 23.500 240.940 23.760 ;
        RECT 491.380 23.500 491.640 23.760 ;
      LAYER met2 ;
        RECT 495.980 1600.450 496.260 1604.000 ;
        RECT 491.440 1600.310 496.260 1600.450 ;
        RECT 491.440 1511.290 491.580 1600.310 ;
        RECT 495.980 1600.000 496.260 1600.310 ;
        RECT 490.460 1510.970 490.720 1511.290 ;
        RECT 491.380 1510.970 491.640 1511.290 ;
        RECT 490.520 1510.690 490.660 1510.970 ;
        RECT 490.520 1510.550 491.120 1510.690 ;
        RECT 490.980 1442.270 491.120 1510.550 ;
        RECT 490.920 1441.950 491.180 1442.270 ;
        RECT 491.840 1442.125 492.100 1442.270 ;
        RECT 491.830 1441.755 492.110 1442.125 ;
        RECT 492.750 1441.755 493.030 1442.125 ;
        RECT 492.820 1393.730 492.960 1441.755 ;
        RECT 492.360 1393.590 492.960 1393.730 ;
        RECT 492.360 1345.710 492.500 1393.590 ;
        RECT 491.840 1345.390 492.100 1345.710 ;
        RECT 492.300 1345.390 492.560 1345.710 ;
        RECT 491.900 1316.890 492.040 1345.390 ;
        RECT 490.980 1316.750 492.040 1316.890 ;
        RECT 490.980 1304.230 491.120 1316.750 ;
        RECT 490.920 1303.910 491.180 1304.230 ;
        RECT 491.380 1255.970 491.640 1256.290 ;
        RECT 491.440 1221.010 491.580 1255.970 ;
        RECT 490.980 1220.870 491.580 1221.010 ;
        RECT 490.980 1207.525 491.120 1220.870 ;
        RECT 489.990 1207.155 490.270 1207.525 ;
        RECT 490.910 1207.155 491.190 1207.525 ;
        RECT 490.060 1159.390 490.200 1207.155 ;
        RECT 490.000 1159.070 490.260 1159.390 ;
        RECT 491.380 1159.070 491.640 1159.390 ;
        RECT 491.440 1124.450 491.580 1159.070 ;
        RECT 490.980 1124.310 491.580 1124.450 ;
        RECT 490.980 1110.965 491.120 1124.310 ;
        RECT 489.990 1110.595 490.270 1110.965 ;
        RECT 490.910 1110.595 491.190 1110.965 ;
        RECT 490.060 1062.830 490.200 1110.595 ;
        RECT 490.000 1062.510 490.260 1062.830 ;
        RECT 491.380 1062.510 491.640 1062.830 ;
        RECT 491.440 1027.890 491.580 1062.510 ;
        RECT 490.980 1027.750 491.580 1027.890 ;
        RECT 490.980 1014.405 491.120 1027.750 ;
        RECT 489.990 1014.035 490.270 1014.405 ;
        RECT 490.910 1014.035 491.190 1014.405 ;
        RECT 490.060 966.270 490.200 1014.035 ;
        RECT 490.000 965.950 490.260 966.270 ;
        RECT 491.380 965.950 491.640 966.270 ;
        RECT 491.440 931.330 491.580 965.950 ;
        RECT 490.980 931.190 491.580 931.330 ;
        RECT 490.980 917.845 491.120 931.190 ;
        RECT 489.990 917.475 490.270 917.845 ;
        RECT 490.910 917.475 491.190 917.845 ;
        RECT 490.060 869.710 490.200 917.475 ;
        RECT 490.000 869.390 490.260 869.710 ;
        RECT 491.380 869.390 491.640 869.710 ;
        RECT 491.440 834.770 491.580 869.390 ;
        RECT 490.980 834.630 491.580 834.770 ;
        RECT 490.980 821.090 491.120 834.630 ;
        RECT 490.000 820.770 490.260 821.090 ;
        RECT 490.920 820.770 491.180 821.090 ;
        RECT 490.060 773.005 490.200 820.770 ;
        RECT 489.990 772.635 490.270 773.005 ;
        RECT 491.370 772.635 491.650 773.005 ;
        RECT 491.440 738.210 491.580 772.635 ;
        RECT 490.980 738.070 491.580 738.210 ;
        RECT 490.980 700.130 491.120 738.070 ;
        RECT 490.060 699.990 491.120 700.130 ;
        RECT 490.060 676.445 490.200 699.990 ;
        RECT 489.990 676.075 490.270 676.445 ;
        RECT 491.370 676.075 491.650 676.445 ;
        RECT 491.440 641.650 491.580 676.075 ;
        RECT 490.980 641.510 491.580 641.650 ;
        RECT 490.980 603.570 491.120 641.510 ;
        RECT 490.060 603.430 491.120 603.570 ;
        RECT 490.060 579.885 490.200 603.430 ;
        RECT 489.990 579.515 490.270 579.885 ;
        RECT 491.370 579.515 491.650 579.885 ;
        RECT 491.440 545.090 491.580 579.515 ;
        RECT 490.980 544.950 491.580 545.090 ;
        RECT 490.980 507.010 491.120 544.950 ;
        RECT 490.060 506.870 491.120 507.010 ;
        RECT 490.060 483.325 490.200 506.870 ;
        RECT 489.990 482.955 490.270 483.325 ;
        RECT 491.370 482.955 491.650 483.325 ;
        RECT 491.440 448.530 491.580 482.955 ;
        RECT 490.520 448.390 491.580 448.530 ;
        RECT 490.520 434.850 490.660 448.390 ;
        RECT 490.460 434.530 490.720 434.850 ;
        RECT 490.000 386.250 490.260 386.570 ;
        RECT 490.060 338.630 490.200 386.250 ;
        RECT 490.000 338.310 490.260 338.630 ;
        RECT 490.460 337.970 490.720 338.290 ;
        RECT 490.520 303.610 490.660 337.970 ;
        RECT 490.460 303.290 490.720 303.610 ;
        RECT 491.380 303.290 491.640 303.610 ;
        RECT 491.440 289.670 491.580 303.290 ;
        RECT 491.380 289.350 491.640 289.670 ;
        RECT 490.920 241.410 491.180 241.730 ;
        RECT 490.980 207.130 491.120 241.410 ;
        RECT 490.520 207.050 491.120 207.130 ;
        RECT 490.460 206.990 491.120 207.050 ;
        RECT 490.460 206.730 490.720 206.990 ;
        RECT 491.380 206.730 491.640 207.050 ;
        RECT 491.440 193.110 491.580 206.730 ;
        RECT 491.380 192.790 491.640 193.110 ;
        RECT 490.920 144.850 491.180 145.170 ;
        RECT 490.980 110.570 491.120 144.850 ;
        RECT 490.520 110.490 491.120 110.570 ;
        RECT 490.460 110.430 491.120 110.490 ;
        RECT 490.460 110.170 490.720 110.430 ;
        RECT 491.380 110.170 491.640 110.490 ;
        RECT 491.440 96.550 491.580 110.170 ;
        RECT 491.380 96.230 491.640 96.550 ;
        RECT 491.380 48.290 491.640 48.610 ;
        RECT 491.440 23.790 491.580 48.290 ;
        RECT 240.680 23.470 240.940 23.790 ;
        RECT 491.380 23.470 491.640 23.790 ;
        RECT 240.740 2.400 240.880 23.470 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 491.830 1441.800 492.110 1442.080 ;
        RECT 492.750 1441.800 493.030 1442.080 ;
        RECT 489.990 1207.200 490.270 1207.480 ;
        RECT 490.910 1207.200 491.190 1207.480 ;
        RECT 489.990 1110.640 490.270 1110.920 ;
        RECT 490.910 1110.640 491.190 1110.920 ;
        RECT 489.990 1014.080 490.270 1014.360 ;
        RECT 490.910 1014.080 491.190 1014.360 ;
        RECT 489.990 917.520 490.270 917.800 ;
        RECT 490.910 917.520 491.190 917.800 ;
        RECT 489.990 772.680 490.270 772.960 ;
        RECT 491.370 772.680 491.650 772.960 ;
        RECT 489.990 676.120 490.270 676.400 ;
        RECT 491.370 676.120 491.650 676.400 ;
        RECT 489.990 579.560 490.270 579.840 ;
        RECT 491.370 579.560 491.650 579.840 ;
        RECT 489.990 483.000 490.270 483.280 ;
        RECT 491.370 483.000 491.650 483.280 ;
      LAYER met3 ;
        RECT 491.805 1442.090 492.135 1442.105 ;
        RECT 492.725 1442.090 493.055 1442.105 ;
        RECT 491.805 1441.790 493.055 1442.090 ;
        RECT 491.805 1441.775 492.135 1441.790 ;
        RECT 492.725 1441.775 493.055 1441.790 ;
        RECT 489.965 1207.490 490.295 1207.505 ;
        RECT 490.885 1207.490 491.215 1207.505 ;
        RECT 489.965 1207.190 491.215 1207.490 ;
        RECT 489.965 1207.175 490.295 1207.190 ;
        RECT 490.885 1207.175 491.215 1207.190 ;
        RECT 489.965 1110.930 490.295 1110.945 ;
        RECT 490.885 1110.930 491.215 1110.945 ;
        RECT 489.965 1110.630 491.215 1110.930 ;
        RECT 489.965 1110.615 490.295 1110.630 ;
        RECT 490.885 1110.615 491.215 1110.630 ;
        RECT 489.965 1014.370 490.295 1014.385 ;
        RECT 490.885 1014.370 491.215 1014.385 ;
        RECT 489.965 1014.070 491.215 1014.370 ;
        RECT 489.965 1014.055 490.295 1014.070 ;
        RECT 490.885 1014.055 491.215 1014.070 ;
        RECT 489.965 917.810 490.295 917.825 ;
        RECT 490.885 917.810 491.215 917.825 ;
        RECT 489.965 917.510 491.215 917.810 ;
        RECT 489.965 917.495 490.295 917.510 ;
        RECT 490.885 917.495 491.215 917.510 ;
        RECT 489.965 772.970 490.295 772.985 ;
        RECT 491.345 772.970 491.675 772.985 ;
        RECT 489.965 772.670 491.675 772.970 ;
        RECT 489.965 772.655 490.295 772.670 ;
        RECT 491.345 772.655 491.675 772.670 ;
        RECT 489.965 676.410 490.295 676.425 ;
        RECT 491.345 676.410 491.675 676.425 ;
        RECT 489.965 676.110 491.675 676.410 ;
        RECT 489.965 676.095 490.295 676.110 ;
        RECT 491.345 676.095 491.675 676.110 ;
        RECT 489.965 579.850 490.295 579.865 ;
        RECT 491.345 579.850 491.675 579.865 ;
        RECT 489.965 579.550 491.675 579.850 ;
        RECT 489.965 579.535 490.295 579.550 ;
        RECT 491.345 579.535 491.675 579.550 ;
        RECT 489.965 483.290 490.295 483.305 ;
        RECT 491.345 483.290 491.675 483.305 ;
        RECT 489.965 482.990 491.675 483.290 ;
        RECT 489.965 482.975 490.295 482.990 ;
        RECT 491.345 482.975 491.675 482.990 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 504.765 1256.045 504.935 1304.155 ;
        RECT 503.845 386.325 504.015 434.775 ;
        RECT 504.765 241.485 504.935 289.595 ;
        RECT 504.765 144.925 504.935 193.035 ;
        RECT 505.225 61.285 505.395 96.475 ;
      LAYER mcon ;
        RECT 504.765 1303.985 504.935 1304.155 ;
        RECT 503.845 434.605 504.015 434.775 ;
        RECT 504.765 289.425 504.935 289.595 ;
        RECT 504.765 192.865 504.935 193.035 ;
        RECT 505.225 96.305 505.395 96.475 ;
      LAYER met1 ;
        RECT 504.230 1511.200 504.550 1511.260 ;
        RECT 505.150 1511.200 505.470 1511.260 ;
        RECT 504.230 1511.060 505.470 1511.200 ;
        RECT 504.230 1511.000 504.550 1511.060 ;
        RECT 505.150 1511.000 505.470 1511.060 ;
        RECT 504.230 1442.180 504.550 1442.240 ;
        RECT 505.610 1442.180 505.930 1442.240 ;
        RECT 504.230 1442.040 505.930 1442.180 ;
        RECT 504.230 1441.980 504.550 1442.040 ;
        RECT 505.610 1441.980 505.930 1442.040 ;
        RECT 506.070 1393.900 506.390 1393.960 ;
        RECT 506.530 1393.900 506.850 1393.960 ;
        RECT 506.070 1393.760 506.850 1393.900 ;
        RECT 506.070 1393.700 506.390 1393.760 ;
        RECT 506.530 1393.700 506.850 1393.760 ;
        RECT 504.690 1304.140 505.010 1304.200 ;
        RECT 504.495 1304.000 505.010 1304.140 ;
        RECT 504.690 1303.940 505.010 1304.000 ;
        RECT 504.705 1256.200 504.995 1256.245 ;
        RECT 505.150 1256.200 505.470 1256.260 ;
        RECT 504.705 1256.060 505.470 1256.200 ;
        RECT 504.705 1256.015 504.995 1256.060 ;
        RECT 505.150 1256.000 505.470 1256.060 ;
        RECT 504.690 1207.240 505.010 1207.300 ;
        RECT 505.150 1207.240 505.470 1207.300 ;
        RECT 504.690 1207.100 505.470 1207.240 ;
        RECT 504.690 1207.040 505.010 1207.100 ;
        RECT 505.150 1207.040 505.470 1207.100 ;
        RECT 504.690 1110.680 505.010 1110.740 ;
        RECT 505.150 1110.680 505.470 1110.740 ;
        RECT 504.690 1110.540 505.470 1110.680 ;
        RECT 504.690 1110.480 505.010 1110.540 ;
        RECT 505.150 1110.480 505.470 1110.540 ;
        RECT 504.690 1014.120 505.010 1014.180 ;
        RECT 505.150 1014.120 505.470 1014.180 ;
        RECT 504.690 1013.980 505.470 1014.120 ;
        RECT 504.690 1013.920 505.010 1013.980 ;
        RECT 505.150 1013.920 505.470 1013.980 ;
        RECT 504.690 917.560 505.010 917.620 ;
        RECT 505.150 917.560 505.470 917.620 ;
        RECT 504.690 917.420 505.470 917.560 ;
        RECT 504.690 917.360 505.010 917.420 ;
        RECT 505.150 917.360 505.470 917.420 ;
        RECT 504.690 821.000 505.010 821.060 ;
        RECT 505.150 821.000 505.470 821.060 ;
        RECT 504.690 820.860 505.470 821.000 ;
        RECT 504.690 820.800 505.010 820.860 ;
        RECT 505.150 820.800 505.470 820.860 ;
        RECT 503.785 434.760 504.075 434.805 ;
        RECT 504.230 434.760 504.550 434.820 ;
        RECT 503.785 434.620 504.550 434.760 ;
        RECT 503.785 434.575 504.075 434.620 ;
        RECT 504.230 434.560 504.550 434.620 ;
        RECT 503.770 386.480 504.090 386.540 ;
        RECT 503.575 386.340 504.090 386.480 ;
        RECT 503.770 386.280 504.090 386.340 ;
        RECT 504.230 303.520 504.550 303.580 ;
        RECT 505.150 303.520 505.470 303.580 ;
        RECT 504.230 303.380 505.470 303.520 ;
        RECT 504.230 303.320 504.550 303.380 ;
        RECT 505.150 303.320 505.470 303.380 ;
        RECT 504.705 289.580 504.995 289.625 ;
        RECT 505.150 289.580 505.470 289.640 ;
        RECT 504.705 289.440 505.470 289.580 ;
        RECT 504.705 289.395 504.995 289.440 ;
        RECT 505.150 289.380 505.470 289.440 ;
        RECT 504.690 241.640 505.010 241.700 ;
        RECT 504.495 241.500 505.010 241.640 ;
        RECT 504.690 241.440 505.010 241.500 ;
        RECT 504.230 206.960 504.550 207.020 ;
        RECT 505.150 206.960 505.470 207.020 ;
        RECT 504.230 206.820 505.470 206.960 ;
        RECT 504.230 206.760 504.550 206.820 ;
        RECT 505.150 206.760 505.470 206.820 ;
        RECT 504.705 193.020 504.995 193.065 ;
        RECT 505.150 193.020 505.470 193.080 ;
        RECT 504.705 192.880 505.470 193.020 ;
        RECT 504.705 192.835 504.995 192.880 ;
        RECT 505.150 192.820 505.470 192.880 ;
        RECT 504.690 145.080 505.010 145.140 ;
        RECT 504.495 144.940 505.010 145.080 ;
        RECT 504.690 144.880 505.010 144.940 ;
        RECT 504.230 110.400 504.550 110.460 ;
        RECT 505.150 110.400 505.470 110.460 ;
        RECT 504.230 110.260 505.470 110.400 ;
        RECT 504.230 110.200 504.550 110.260 ;
        RECT 505.150 110.200 505.470 110.260 ;
        RECT 505.150 96.460 505.470 96.520 ;
        RECT 504.955 96.320 505.470 96.460 ;
        RECT 505.150 96.260 505.470 96.320 ;
        RECT 505.150 61.440 505.470 61.500 ;
        RECT 504.955 61.300 505.470 61.440 ;
        RECT 505.150 61.240 505.470 61.300 ;
        RECT 258.130 23.020 258.450 23.080 ;
        RECT 505.150 23.020 505.470 23.080 ;
        RECT 258.130 22.880 505.470 23.020 ;
        RECT 258.130 22.820 258.450 22.880 ;
        RECT 505.150 22.820 505.470 22.880 ;
      LAYER via ;
        RECT 504.260 1511.000 504.520 1511.260 ;
        RECT 505.180 1511.000 505.440 1511.260 ;
        RECT 504.260 1441.980 504.520 1442.240 ;
        RECT 505.640 1441.980 505.900 1442.240 ;
        RECT 506.100 1393.700 506.360 1393.960 ;
        RECT 506.560 1393.700 506.820 1393.960 ;
        RECT 504.720 1303.940 504.980 1304.200 ;
        RECT 505.180 1256.000 505.440 1256.260 ;
        RECT 504.720 1207.040 504.980 1207.300 ;
        RECT 505.180 1207.040 505.440 1207.300 ;
        RECT 504.720 1110.480 504.980 1110.740 ;
        RECT 505.180 1110.480 505.440 1110.740 ;
        RECT 504.720 1013.920 504.980 1014.180 ;
        RECT 505.180 1013.920 505.440 1014.180 ;
        RECT 504.720 917.360 504.980 917.620 ;
        RECT 505.180 917.360 505.440 917.620 ;
        RECT 504.720 820.800 504.980 821.060 ;
        RECT 505.180 820.800 505.440 821.060 ;
        RECT 504.260 434.560 504.520 434.820 ;
        RECT 503.800 386.280 504.060 386.540 ;
        RECT 504.260 303.320 504.520 303.580 ;
        RECT 505.180 303.320 505.440 303.580 ;
        RECT 505.180 289.380 505.440 289.640 ;
        RECT 504.720 241.440 504.980 241.700 ;
        RECT 504.260 206.760 504.520 207.020 ;
        RECT 505.180 206.760 505.440 207.020 ;
        RECT 505.180 192.820 505.440 193.080 ;
        RECT 504.720 144.880 504.980 145.140 ;
        RECT 504.260 110.200 504.520 110.460 ;
        RECT 505.180 110.200 505.440 110.460 ;
        RECT 505.180 96.260 505.440 96.520 ;
        RECT 505.180 61.240 505.440 61.500 ;
        RECT 258.160 22.820 258.420 23.080 ;
        RECT 505.180 22.820 505.440 23.080 ;
      LAYER met2 ;
        RECT 510.240 1600.450 510.520 1604.000 ;
        RECT 506.620 1600.310 510.520 1600.450 ;
        RECT 506.620 1580.050 506.760 1600.310 ;
        RECT 510.240 1600.000 510.520 1600.310 ;
        RECT 505.240 1579.910 506.760 1580.050 ;
        RECT 505.240 1511.290 505.380 1579.910 ;
        RECT 504.260 1510.970 504.520 1511.290 ;
        RECT 505.180 1510.970 505.440 1511.290 ;
        RECT 504.320 1510.690 504.460 1510.970 ;
        RECT 504.320 1510.550 504.920 1510.690 ;
        RECT 504.780 1467.170 504.920 1510.550 ;
        RECT 504.320 1467.030 504.920 1467.170 ;
        RECT 504.320 1442.270 504.460 1467.030 ;
        RECT 504.260 1441.950 504.520 1442.270 ;
        RECT 505.640 1442.125 505.900 1442.270 ;
        RECT 505.630 1441.755 505.910 1442.125 ;
        RECT 506.550 1441.755 506.830 1442.125 ;
        RECT 506.160 1393.990 506.300 1394.145 ;
        RECT 506.620 1393.990 506.760 1441.755 ;
        RECT 506.100 1393.730 506.360 1393.990 ;
        RECT 506.560 1393.845 506.820 1393.990 ;
        RECT 506.550 1393.730 506.830 1393.845 ;
        RECT 506.100 1393.670 506.830 1393.730 ;
        RECT 506.160 1393.590 506.830 1393.670 ;
        RECT 506.550 1393.475 506.830 1393.590 ;
        RECT 504.710 1392.795 504.990 1393.165 ;
        RECT 504.780 1304.230 504.920 1392.795 ;
        RECT 504.720 1303.910 504.980 1304.230 ;
        RECT 505.180 1255.970 505.440 1256.290 ;
        RECT 505.240 1221.010 505.380 1255.970 ;
        RECT 504.780 1220.870 505.380 1221.010 ;
        RECT 504.780 1207.330 504.920 1220.870 ;
        RECT 504.720 1207.010 504.980 1207.330 ;
        RECT 505.180 1207.010 505.440 1207.330 ;
        RECT 505.240 1124.450 505.380 1207.010 ;
        RECT 504.780 1124.310 505.380 1124.450 ;
        RECT 504.780 1110.770 504.920 1124.310 ;
        RECT 504.720 1110.450 504.980 1110.770 ;
        RECT 505.180 1110.450 505.440 1110.770 ;
        RECT 505.240 1027.890 505.380 1110.450 ;
        RECT 504.780 1027.750 505.380 1027.890 ;
        RECT 504.780 1014.210 504.920 1027.750 ;
        RECT 504.720 1013.890 504.980 1014.210 ;
        RECT 505.180 1013.890 505.440 1014.210 ;
        RECT 505.240 931.330 505.380 1013.890 ;
        RECT 504.780 931.190 505.380 931.330 ;
        RECT 504.780 917.650 504.920 931.190 ;
        RECT 504.720 917.330 504.980 917.650 ;
        RECT 505.180 917.330 505.440 917.650 ;
        RECT 505.240 834.770 505.380 917.330 ;
        RECT 504.780 834.630 505.380 834.770 ;
        RECT 504.780 821.090 504.920 834.630 ;
        RECT 504.720 820.770 504.980 821.090 ;
        RECT 505.180 820.770 505.440 821.090 ;
        RECT 505.240 738.210 505.380 820.770 ;
        RECT 504.780 738.070 505.380 738.210 ;
        RECT 504.780 700.130 504.920 738.070 ;
        RECT 503.860 699.990 504.920 700.130 ;
        RECT 503.860 676.445 504.000 699.990 ;
        RECT 503.790 676.075 504.070 676.445 ;
        RECT 505.170 676.075 505.450 676.445 ;
        RECT 505.240 641.650 505.380 676.075 ;
        RECT 504.780 641.510 505.380 641.650 ;
        RECT 504.780 603.570 504.920 641.510 ;
        RECT 503.860 603.430 504.920 603.570 ;
        RECT 503.860 579.885 504.000 603.430 ;
        RECT 503.790 579.515 504.070 579.885 ;
        RECT 505.170 579.515 505.450 579.885 ;
        RECT 505.240 545.090 505.380 579.515 ;
        RECT 504.780 544.950 505.380 545.090 ;
        RECT 504.780 507.010 504.920 544.950 ;
        RECT 503.860 506.870 504.920 507.010 ;
        RECT 503.860 483.325 504.000 506.870 ;
        RECT 503.790 482.955 504.070 483.325 ;
        RECT 505.170 482.955 505.450 483.325 ;
        RECT 505.240 448.530 505.380 482.955 ;
        RECT 504.320 448.390 505.380 448.530 ;
        RECT 504.320 434.850 504.460 448.390 ;
        RECT 504.260 434.530 504.520 434.850 ;
        RECT 503.800 386.250 504.060 386.570 ;
        RECT 503.860 351.290 504.000 386.250 ;
        RECT 503.860 351.150 504.460 351.290 ;
        RECT 504.320 303.610 504.460 351.150 ;
        RECT 504.260 303.290 504.520 303.610 ;
        RECT 505.180 303.290 505.440 303.610 ;
        RECT 505.240 289.670 505.380 303.290 ;
        RECT 505.180 289.350 505.440 289.670 ;
        RECT 504.720 241.410 504.980 241.730 ;
        RECT 504.780 207.130 504.920 241.410 ;
        RECT 504.320 207.050 504.920 207.130 ;
        RECT 504.260 206.990 504.920 207.050 ;
        RECT 504.260 206.730 504.520 206.990 ;
        RECT 505.180 206.730 505.440 207.050 ;
        RECT 505.240 193.110 505.380 206.730 ;
        RECT 505.180 192.790 505.440 193.110 ;
        RECT 504.720 144.850 504.980 145.170 ;
        RECT 504.780 110.570 504.920 144.850 ;
        RECT 504.320 110.490 504.920 110.570 ;
        RECT 504.260 110.430 504.920 110.490 ;
        RECT 504.260 110.170 504.520 110.430 ;
        RECT 505.180 110.170 505.440 110.490 ;
        RECT 505.240 96.550 505.380 110.170 ;
        RECT 505.180 96.230 505.440 96.550 ;
        RECT 505.180 61.210 505.440 61.530 ;
        RECT 505.240 23.110 505.380 61.210 ;
        RECT 258.160 22.790 258.420 23.110 ;
        RECT 505.180 22.790 505.440 23.110 ;
        RECT 258.220 2.400 258.360 22.790 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 505.630 1441.800 505.910 1442.080 ;
        RECT 506.550 1441.800 506.830 1442.080 ;
        RECT 506.550 1393.520 506.830 1393.800 ;
        RECT 504.710 1392.840 504.990 1393.120 ;
        RECT 503.790 676.120 504.070 676.400 ;
        RECT 505.170 676.120 505.450 676.400 ;
        RECT 503.790 579.560 504.070 579.840 ;
        RECT 505.170 579.560 505.450 579.840 ;
        RECT 503.790 483.000 504.070 483.280 ;
        RECT 505.170 483.000 505.450 483.280 ;
      LAYER met3 ;
        RECT 505.605 1442.090 505.935 1442.105 ;
        RECT 506.525 1442.090 506.855 1442.105 ;
        RECT 505.605 1441.790 506.855 1442.090 ;
        RECT 505.605 1441.775 505.935 1441.790 ;
        RECT 506.525 1441.775 506.855 1441.790 ;
        RECT 506.525 1393.810 506.855 1393.825 ;
        RECT 506.525 1393.510 507.530 1393.810 ;
        RECT 506.525 1393.495 506.855 1393.510 ;
        RECT 504.685 1393.130 505.015 1393.145 ;
        RECT 507.230 1393.130 507.530 1393.510 ;
        RECT 504.685 1392.830 507.530 1393.130 ;
        RECT 504.685 1392.815 505.015 1392.830 ;
        RECT 503.765 676.410 504.095 676.425 ;
        RECT 505.145 676.410 505.475 676.425 ;
        RECT 503.765 676.110 505.475 676.410 ;
        RECT 503.765 676.095 504.095 676.110 ;
        RECT 505.145 676.095 505.475 676.110 ;
        RECT 503.765 579.850 504.095 579.865 ;
        RECT 505.145 579.850 505.475 579.865 ;
        RECT 503.765 579.550 505.475 579.850 ;
        RECT 503.765 579.535 504.095 579.550 ;
        RECT 505.145 579.535 505.475 579.550 ;
        RECT 503.765 483.290 504.095 483.305 ;
        RECT 505.145 483.290 505.475 483.305 ;
        RECT 503.765 482.990 505.475 483.290 ;
        RECT 503.765 482.975 504.095 482.990 ;
        RECT 505.145 482.975 505.475 482.990 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 23.360 276.390 23.420 ;
        RECT 524.930 23.360 525.250 23.420 ;
        RECT 276.070 23.220 525.250 23.360 ;
        RECT 276.070 23.160 276.390 23.220 ;
        RECT 524.930 23.160 525.250 23.220 ;
      LAYER via ;
        RECT 276.100 23.160 276.360 23.420 ;
        RECT 524.960 23.160 525.220 23.420 ;
      LAYER met2 ;
        RECT 524.960 1600.000 525.240 1604.000 ;
        RECT 525.020 23.450 525.160 1600.000 ;
        RECT 276.100 23.130 276.360 23.450 ;
        RECT 524.960 23.130 525.220 23.450 ;
        RECT 276.160 2.400 276.300 23.130 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 22.680 294.330 22.740 ;
        RECT 538.730 22.680 539.050 22.740 ;
        RECT 294.010 22.540 539.050 22.680 ;
        RECT 294.010 22.480 294.330 22.540 ;
        RECT 538.730 22.480 539.050 22.540 ;
      LAYER via ;
        RECT 294.040 22.480 294.300 22.740 ;
        RECT 538.760 22.480 539.020 22.740 ;
      LAYER met2 ;
        RECT 539.680 1600.450 539.960 1604.000 ;
        RECT 538.820 1600.310 539.960 1600.450 ;
        RECT 538.820 22.770 538.960 1600.310 ;
        RECT 539.680 1600.000 539.960 1600.310 ;
        RECT 294.040 22.450 294.300 22.770 ;
        RECT 538.760 22.450 539.020 22.770 ;
        RECT 294.100 2.400 294.240 22.450 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 24.380 312.270 24.440 ;
        RECT 552.070 24.380 552.390 24.440 ;
        RECT 311.950 24.240 552.390 24.380 ;
        RECT 311.950 24.180 312.270 24.240 ;
        RECT 552.070 24.180 552.390 24.240 ;
      LAYER via ;
        RECT 311.980 24.180 312.240 24.440 ;
        RECT 552.100 24.180 552.360 24.440 ;
      LAYER met2 ;
        RECT 553.940 1600.450 554.220 1604.000 ;
        RECT 552.160 1600.310 554.220 1600.450 ;
        RECT 552.160 24.470 552.300 1600.310 ;
        RECT 553.940 1600.000 554.220 1600.310 ;
        RECT 311.980 24.150 312.240 24.470 ;
        RECT 552.100 24.150 552.360 24.470 ;
        RECT 312.040 2.400 312.180 24.150 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 24.040 330.210 24.100 ;
        RECT 565.870 24.040 566.190 24.100 ;
        RECT 329.890 23.900 566.190 24.040 ;
        RECT 329.890 23.840 330.210 23.900 ;
        RECT 565.870 23.840 566.190 23.900 ;
      LAYER via ;
        RECT 329.920 23.840 330.180 24.100 ;
        RECT 565.900 23.840 566.160 24.100 ;
      LAYER met2 ;
        RECT 568.660 1600.450 568.940 1604.000 ;
        RECT 565.960 1600.310 568.940 1600.450 ;
        RECT 565.960 24.130 566.100 1600.310 ;
        RECT 568.660 1600.000 568.940 1600.310 ;
        RECT 329.920 23.810 330.180 24.130 ;
        RECT 565.900 23.810 566.160 24.130 ;
        RECT 329.980 2.400 330.120 23.810 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 25.060 347.690 25.120 ;
        RECT 579.670 25.060 579.990 25.120 ;
        RECT 347.370 24.920 579.990 25.060 ;
        RECT 347.370 24.860 347.690 24.920 ;
        RECT 579.670 24.860 579.990 24.920 ;
      LAYER via ;
        RECT 347.400 24.860 347.660 25.120 ;
        RECT 579.700 24.860 579.960 25.120 ;
      LAYER met2 ;
        RECT 582.920 1600.450 583.200 1604.000 ;
        RECT 579.760 1600.310 583.200 1600.450 ;
        RECT 579.760 25.150 579.900 1600.310 ;
        RECT 582.920 1600.000 583.200 1600.310 ;
        RECT 347.400 24.830 347.660 25.150 ;
        RECT 579.700 24.830 579.960 25.150 ;
        RECT 347.460 2.400 347.600 24.830 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 24.720 365.630 24.780 ;
        RECT 593.470 24.720 593.790 24.780 ;
        RECT 365.310 24.580 593.790 24.720 ;
        RECT 365.310 24.520 365.630 24.580 ;
        RECT 593.470 24.520 593.790 24.580 ;
      LAYER via ;
        RECT 365.340 24.520 365.600 24.780 ;
        RECT 593.500 24.520 593.760 24.780 ;
      LAYER met2 ;
        RECT 597.640 1600.450 597.920 1604.000 ;
        RECT 593.560 1600.310 597.920 1600.450 ;
        RECT 593.560 24.810 593.700 1600.310 ;
        RECT 597.640 1600.000 597.920 1600.310 ;
        RECT 365.340 24.490 365.600 24.810 ;
        RECT 593.500 24.490 593.760 24.810 ;
        RECT 365.400 2.400 365.540 24.490 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 25.400 383.570 25.460 ;
        RECT 607.730 25.400 608.050 25.460 ;
        RECT 383.250 25.260 608.050 25.400 ;
        RECT 383.250 25.200 383.570 25.260 ;
        RECT 607.730 25.200 608.050 25.260 ;
      LAYER via ;
        RECT 383.280 25.200 383.540 25.460 ;
        RECT 607.760 25.200 608.020 25.460 ;
      LAYER met2 ;
        RECT 612.360 1600.450 612.640 1604.000 ;
        RECT 607.820 1600.310 612.640 1600.450 ;
        RECT 607.820 25.490 607.960 1600.310 ;
        RECT 612.360 1600.000 612.640 1600.310 ;
        RECT 383.280 25.170 383.540 25.490 ;
        RECT 607.760 25.170 608.020 25.490 ;
        RECT 383.340 2.400 383.480 25.170 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 621.605 1497.445 621.775 1545.555 ;
        RECT 621.605 1449.165 621.775 1463.275 ;
        RECT 621.605 786.505 621.775 821.015 ;
        RECT 621.605 689.605 621.775 724.455 ;
        RECT 621.605 593.045 621.775 627.895 ;
        RECT 621.605 496.485 621.775 531.335 ;
        RECT 621.605 386.325 621.775 434.775 ;
        RECT 621.605 338.045 621.775 385.815 ;
        RECT 621.605 241.485 621.775 289.595 ;
        RECT 621.605 96.645 621.775 144.755 ;
      LAYER mcon ;
        RECT 621.605 1545.385 621.775 1545.555 ;
        RECT 621.605 1463.105 621.775 1463.275 ;
        RECT 621.605 820.845 621.775 821.015 ;
        RECT 621.605 724.285 621.775 724.455 ;
        RECT 621.605 627.725 621.775 627.895 ;
        RECT 621.605 531.165 621.775 531.335 ;
        RECT 621.605 434.605 621.775 434.775 ;
        RECT 621.605 385.645 621.775 385.815 ;
        RECT 621.605 289.425 621.775 289.595 ;
        RECT 621.605 144.585 621.775 144.755 ;
      LAYER met1 ;
        RECT 621.070 1559.140 621.390 1559.200 ;
        RECT 621.990 1559.140 622.310 1559.200 ;
        RECT 621.070 1559.000 622.310 1559.140 ;
        RECT 621.070 1558.940 621.390 1559.000 ;
        RECT 621.990 1558.940 622.310 1559.000 ;
        RECT 621.545 1545.540 621.835 1545.585 ;
        RECT 621.990 1545.540 622.310 1545.600 ;
        RECT 621.545 1545.400 622.310 1545.540 ;
        RECT 621.545 1545.355 621.835 1545.400 ;
        RECT 621.990 1545.340 622.310 1545.400 ;
        RECT 621.530 1497.600 621.850 1497.660 ;
        RECT 621.335 1497.460 621.850 1497.600 ;
        RECT 621.530 1497.400 621.850 1497.460 ;
        RECT 621.530 1463.260 621.850 1463.320 ;
        RECT 621.335 1463.120 621.850 1463.260 ;
        RECT 621.530 1463.060 621.850 1463.120 ;
        RECT 621.530 1449.320 621.850 1449.380 ;
        RECT 621.335 1449.180 621.850 1449.320 ;
        RECT 621.530 1449.120 621.850 1449.180 ;
        RECT 621.070 1318.080 621.390 1318.140 ;
        RECT 621.990 1318.080 622.310 1318.140 ;
        RECT 621.070 1317.940 622.310 1318.080 ;
        RECT 621.070 1317.880 621.390 1317.940 ;
        RECT 621.990 1317.880 622.310 1317.940 ;
        RECT 621.070 1221.520 621.390 1221.580 ;
        RECT 621.990 1221.520 622.310 1221.580 ;
        RECT 621.070 1221.380 622.310 1221.520 ;
        RECT 621.070 1221.320 621.390 1221.380 ;
        RECT 621.990 1221.320 622.310 1221.380 ;
        RECT 621.070 1124.960 621.390 1125.020 ;
        RECT 621.990 1124.960 622.310 1125.020 ;
        RECT 621.070 1124.820 622.310 1124.960 ;
        RECT 621.070 1124.760 621.390 1124.820 ;
        RECT 621.990 1124.760 622.310 1124.820 ;
        RECT 621.070 1028.400 621.390 1028.460 ;
        RECT 621.990 1028.400 622.310 1028.460 ;
        RECT 621.070 1028.260 622.310 1028.400 ;
        RECT 621.070 1028.200 621.390 1028.260 ;
        RECT 621.990 1028.200 622.310 1028.260 ;
        RECT 621.070 931.840 621.390 931.900 ;
        RECT 621.990 931.840 622.310 931.900 ;
        RECT 621.070 931.700 622.310 931.840 ;
        RECT 621.070 931.640 621.390 931.700 ;
        RECT 621.990 931.640 622.310 931.700 ;
        RECT 621.990 869.620 622.310 869.680 ;
        RECT 622.910 869.620 623.230 869.680 ;
        RECT 621.990 869.480 623.230 869.620 ;
        RECT 621.990 869.420 622.310 869.480 ;
        RECT 622.910 869.420 623.230 869.480 ;
        RECT 621.070 835.280 621.390 835.340 ;
        RECT 621.990 835.280 622.310 835.340 ;
        RECT 621.070 835.140 622.310 835.280 ;
        RECT 621.070 835.080 621.390 835.140 ;
        RECT 621.990 835.080 622.310 835.140 ;
        RECT 621.530 821.000 621.850 821.060 ;
        RECT 621.335 820.860 621.850 821.000 ;
        RECT 621.530 820.800 621.850 820.860 ;
        RECT 621.530 786.660 621.850 786.720 ;
        RECT 621.335 786.520 621.850 786.660 ;
        RECT 621.530 786.460 621.850 786.520 ;
        RECT 621.070 738.380 621.390 738.440 ;
        RECT 621.990 738.380 622.310 738.440 ;
        RECT 621.070 738.240 622.310 738.380 ;
        RECT 621.070 738.180 621.390 738.240 ;
        RECT 621.990 738.180 622.310 738.240 ;
        RECT 621.530 724.440 621.850 724.500 ;
        RECT 621.335 724.300 621.850 724.440 ;
        RECT 621.530 724.240 621.850 724.300 ;
        RECT 621.530 689.760 621.850 689.820 ;
        RECT 621.335 689.620 621.850 689.760 ;
        RECT 621.530 689.560 621.850 689.620 ;
        RECT 621.070 641.820 621.390 641.880 ;
        RECT 621.990 641.820 622.310 641.880 ;
        RECT 621.070 641.680 622.310 641.820 ;
        RECT 621.070 641.620 621.390 641.680 ;
        RECT 621.990 641.620 622.310 641.680 ;
        RECT 621.530 627.880 621.850 627.940 ;
        RECT 621.335 627.740 621.850 627.880 ;
        RECT 621.530 627.680 621.850 627.740 ;
        RECT 621.530 593.200 621.850 593.260 ;
        RECT 621.335 593.060 621.850 593.200 ;
        RECT 621.530 593.000 621.850 593.060 ;
        RECT 621.070 545.260 621.390 545.320 ;
        RECT 621.990 545.260 622.310 545.320 ;
        RECT 621.070 545.120 622.310 545.260 ;
        RECT 621.070 545.060 621.390 545.120 ;
        RECT 621.990 545.060 622.310 545.120 ;
        RECT 621.530 531.320 621.850 531.380 ;
        RECT 621.335 531.180 621.850 531.320 ;
        RECT 621.530 531.120 621.850 531.180 ;
        RECT 621.530 496.640 621.850 496.700 ;
        RECT 621.335 496.500 621.850 496.640 ;
        RECT 621.530 496.440 621.850 496.500 ;
        RECT 621.070 448.700 621.390 448.760 ;
        RECT 621.990 448.700 622.310 448.760 ;
        RECT 621.070 448.560 622.310 448.700 ;
        RECT 621.070 448.500 621.390 448.560 ;
        RECT 621.990 448.500 622.310 448.560 ;
        RECT 621.530 434.760 621.850 434.820 ;
        RECT 621.335 434.620 621.850 434.760 ;
        RECT 621.530 434.560 621.850 434.620 ;
        RECT 621.545 386.480 621.835 386.525 ;
        RECT 621.990 386.480 622.310 386.540 ;
        RECT 621.545 386.340 622.310 386.480 ;
        RECT 621.545 386.295 621.835 386.340 ;
        RECT 621.990 386.280 622.310 386.340 ;
        RECT 621.545 385.800 621.835 385.845 ;
        RECT 621.990 385.800 622.310 385.860 ;
        RECT 621.545 385.660 622.310 385.800 ;
        RECT 621.545 385.615 621.835 385.660 ;
        RECT 621.990 385.600 622.310 385.660 ;
        RECT 621.530 338.200 621.850 338.260 ;
        RECT 621.335 338.060 621.850 338.200 ;
        RECT 621.530 338.000 621.850 338.060 ;
        RECT 621.545 289.580 621.835 289.625 ;
        RECT 621.990 289.580 622.310 289.640 ;
        RECT 621.545 289.440 622.310 289.580 ;
        RECT 621.545 289.395 621.835 289.440 ;
        RECT 621.990 289.380 622.310 289.440 ;
        RECT 621.530 241.640 621.850 241.700 ;
        RECT 621.335 241.500 621.850 241.640 ;
        RECT 621.530 241.440 621.850 241.500 ;
        RECT 621.530 144.740 621.850 144.800 ;
        RECT 621.335 144.600 621.850 144.740 ;
        RECT 621.530 144.540 621.850 144.600 ;
        RECT 621.545 96.800 621.835 96.845 ;
        RECT 622.450 96.800 622.770 96.860 ;
        RECT 621.545 96.660 622.770 96.800 ;
        RECT 621.545 96.615 621.835 96.660 ;
        RECT 622.450 96.600 622.770 96.660 ;
        RECT 401.190 17.920 401.510 17.980 ;
        RECT 620.610 17.920 620.930 17.980 ;
        RECT 401.190 17.780 620.930 17.920 ;
        RECT 401.190 17.720 401.510 17.780 ;
        RECT 620.610 17.720 620.930 17.780 ;
      LAYER via ;
        RECT 621.100 1558.940 621.360 1559.200 ;
        RECT 622.020 1558.940 622.280 1559.200 ;
        RECT 622.020 1545.340 622.280 1545.600 ;
        RECT 621.560 1497.400 621.820 1497.660 ;
        RECT 621.560 1463.060 621.820 1463.320 ;
        RECT 621.560 1449.120 621.820 1449.380 ;
        RECT 621.100 1317.880 621.360 1318.140 ;
        RECT 622.020 1317.880 622.280 1318.140 ;
        RECT 621.100 1221.320 621.360 1221.580 ;
        RECT 622.020 1221.320 622.280 1221.580 ;
        RECT 621.100 1124.760 621.360 1125.020 ;
        RECT 622.020 1124.760 622.280 1125.020 ;
        RECT 621.100 1028.200 621.360 1028.460 ;
        RECT 622.020 1028.200 622.280 1028.460 ;
        RECT 621.100 931.640 621.360 931.900 ;
        RECT 622.020 931.640 622.280 931.900 ;
        RECT 622.020 869.420 622.280 869.680 ;
        RECT 622.940 869.420 623.200 869.680 ;
        RECT 621.100 835.080 621.360 835.340 ;
        RECT 622.020 835.080 622.280 835.340 ;
        RECT 621.560 820.800 621.820 821.060 ;
        RECT 621.560 786.460 621.820 786.720 ;
        RECT 621.100 738.180 621.360 738.440 ;
        RECT 622.020 738.180 622.280 738.440 ;
        RECT 621.560 724.240 621.820 724.500 ;
        RECT 621.560 689.560 621.820 689.820 ;
        RECT 621.100 641.620 621.360 641.880 ;
        RECT 622.020 641.620 622.280 641.880 ;
        RECT 621.560 627.680 621.820 627.940 ;
        RECT 621.560 593.000 621.820 593.260 ;
        RECT 621.100 545.060 621.360 545.320 ;
        RECT 622.020 545.060 622.280 545.320 ;
        RECT 621.560 531.120 621.820 531.380 ;
        RECT 621.560 496.440 621.820 496.700 ;
        RECT 621.100 448.500 621.360 448.760 ;
        RECT 622.020 448.500 622.280 448.760 ;
        RECT 621.560 434.560 621.820 434.820 ;
        RECT 622.020 386.280 622.280 386.540 ;
        RECT 622.020 385.600 622.280 385.860 ;
        RECT 621.560 338.000 621.820 338.260 ;
        RECT 622.020 289.380 622.280 289.640 ;
        RECT 621.560 241.440 621.820 241.700 ;
        RECT 621.560 144.540 621.820 144.800 ;
        RECT 622.480 96.600 622.740 96.860 ;
        RECT 401.220 17.720 401.480 17.980 ;
        RECT 620.640 17.720 620.900 17.980 ;
      LAYER met2 ;
        RECT 626.620 1601.130 626.900 1604.000 ;
        RECT 622.540 1600.990 626.900 1601.130 ;
        RECT 622.540 1580.050 622.680 1600.990 ;
        RECT 626.620 1600.000 626.900 1600.990 ;
        RECT 621.160 1579.910 622.680 1580.050 ;
        RECT 621.160 1559.230 621.300 1579.910 ;
        RECT 621.100 1558.910 621.360 1559.230 ;
        RECT 622.020 1558.910 622.280 1559.230 ;
        RECT 622.080 1545.630 622.220 1558.910 ;
        RECT 622.020 1545.310 622.280 1545.630 ;
        RECT 621.560 1497.370 621.820 1497.690 ;
        RECT 621.620 1463.350 621.760 1497.370 ;
        RECT 621.560 1463.030 621.820 1463.350 ;
        RECT 621.560 1449.090 621.820 1449.410 ;
        RECT 621.620 1414.810 621.760 1449.090 ;
        RECT 621.620 1414.670 622.220 1414.810 ;
        RECT 622.080 1318.170 622.220 1414.670 ;
        RECT 621.100 1317.850 621.360 1318.170 ;
        RECT 622.020 1317.850 622.280 1318.170 ;
        RECT 621.160 1317.570 621.300 1317.850 ;
        RECT 621.160 1317.430 621.760 1317.570 ;
        RECT 621.620 1269.970 621.760 1317.430 ;
        RECT 621.620 1269.830 622.220 1269.970 ;
        RECT 622.080 1221.610 622.220 1269.830 ;
        RECT 621.100 1221.290 621.360 1221.610 ;
        RECT 622.020 1221.290 622.280 1221.610 ;
        RECT 621.160 1221.010 621.300 1221.290 ;
        RECT 621.160 1220.870 621.760 1221.010 ;
        RECT 621.620 1173.410 621.760 1220.870 ;
        RECT 621.620 1173.270 622.220 1173.410 ;
        RECT 622.080 1125.050 622.220 1173.270 ;
        RECT 621.100 1124.730 621.360 1125.050 ;
        RECT 622.020 1124.730 622.280 1125.050 ;
        RECT 621.160 1124.450 621.300 1124.730 ;
        RECT 621.160 1124.310 621.760 1124.450 ;
        RECT 621.620 1076.850 621.760 1124.310 ;
        RECT 621.620 1076.710 622.220 1076.850 ;
        RECT 622.080 1028.490 622.220 1076.710 ;
        RECT 621.100 1028.170 621.360 1028.490 ;
        RECT 622.020 1028.170 622.280 1028.490 ;
        RECT 621.160 1027.890 621.300 1028.170 ;
        RECT 621.160 1027.750 621.760 1027.890 ;
        RECT 621.620 980.290 621.760 1027.750 ;
        RECT 621.620 980.150 622.220 980.290 ;
        RECT 622.080 931.930 622.220 980.150 ;
        RECT 621.100 931.610 621.360 931.930 ;
        RECT 622.020 931.610 622.280 931.930 ;
        RECT 621.160 931.330 621.300 931.610 ;
        RECT 621.160 931.190 621.760 931.330 ;
        RECT 621.620 917.845 621.760 931.190 ;
        RECT 621.550 917.475 621.830 917.845 ;
        RECT 622.930 917.475 623.210 917.845 ;
        RECT 623.000 869.710 623.140 917.475 ;
        RECT 622.020 869.390 622.280 869.710 ;
        RECT 622.940 869.390 623.200 869.710 ;
        RECT 622.080 835.370 622.220 869.390 ;
        RECT 621.100 835.050 621.360 835.370 ;
        RECT 622.020 835.050 622.280 835.370 ;
        RECT 621.160 834.770 621.300 835.050 ;
        RECT 621.160 834.630 621.760 834.770 ;
        RECT 621.620 821.090 621.760 834.630 ;
        RECT 621.560 820.770 621.820 821.090 ;
        RECT 621.560 786.430 621.820 786.750 ;
        RECT 621.620 772.890 621.760 786.430 ;
        RECT 621.620 772.750 622.220 772.890 ;
        RECT 622.080 738.470 622.220 772.750 ;
        RECT 621.100 738.210 621.360 738.470 ;
        RECT 621.100 738.150 621.760 738.210 ;
        RECT 622.020 738.150 622.280 738.470 ;
        RECT 621.160 738.070 621.760 738.150 ;
        RECT 621.620 724.530 621.760 738.070 ;
        RECT 621.560 724.210 621.820 724.530 ;
        RECT 621.560 689.530 621.820 689.850 ;
        RECT 621.620 676.330 621.760 689.530 ;
        RECT 621.620 676.190 622.220 676.330 ;
        RECT 622.080 641.910 622.220 676.190 ;
        RECT 621.100 641.650 621.360 641.910 ;
        RECT 621.100 641.590 621.760 641.650 ;
        RECT 622.020 641.590 622.280 641.910 ;
        RECT 621.160 641.510 621.760 641.590 ;
        RECT 621.620 627.970 621.760 641.510 ;
        RECT 621.560 627.650 621.820 627.970 ;
        RECT 621.560 592.970 621.820 593.290 ;
        RECT 621.620 579.770 621.760 592.970 ;
        RECT 621.620 579.630 622.220 579.770 ;
        RECT 622.080 545.350 622.220 579.630 ;
        RECT 621.100 545.090 621.360 545.350 ;
        RECT 621.100 545.030 621.760 545.090 ;
        RECT 622.020 545.030 622.280 545.350 ;
        RECT 621.160 544.950 621.760 545.030 ;
        RECT 621.620 531.410 621.760 544.950 ;
        RECT 621.560 531.090 621.820 531.410 ;
        RECT 621.560 496.410 621.820 496.730 ;
        RECT 621.620 483.210 621.760 496.410 ;
        RECT 621.620 483.070 622.220 483.210 ;
        RECT 622.080 448.790 622.220 483.070 ;
        RECT 621.100 448.530 621.360 448.790 ;
        RECT 621.100 448.470 621.760 448.530 ;
        RECT 622.020 448.470 622.280 448.790 ;
        RECT 621.160 448.390 621.760 448.470 ;
        RECT 621.620 434.850 621.760 448.390 ;
        RECT 621.560 434.530 621.820 434.850 ;
        RECT 622.020 386.250 622.280 386.570 ;
        RECT 622.080 385.890 622.220 386.250 ;
        RECT 622.020 385.570 622.280 385.890 ;
        RECT 621.560 337.970 621.820 338.290 ;
        RECT 621.620 303.690 621.760 337.970 ;
        RECT 621.620 303.550 622.220 303.690 ;
        RECT 622.080 289.670 622.220 303.550 ;
        RECT 622.020 289.350 622.280 289.670 ;
        RECT 621.560 241.410 621.820 241.730 ;
        RECT 621.620 207.130 621.760 241.410 ;
        RECT 621.620 206.990 622.220 207.130 ;
        RECT 622.080 158.850 622.220 206.990 ;
        RECT 621.160 158.710 622.220 158.850 ;
        RECT 621.160 158.170 621.300 158.710 ;
        RECT 621.160 158.030 621.760 158.170 ;
        RECT 621.620 144.830 621.760 158.030 ;
        RECT 621.560 144.510 621.820 144.830 ;
        RECT 622.480 96.570 622.740 96.890 ;
        RECT 622.540 39.850 622.680 96.570 ;
        RECT 621.160 39.710 622.680 39.850 ;
        RECT 621.160 19.450 621.300 39.710 ;
        RECT 620.700 19.310 621.300 19.450 ;
        RECT 620.700 18.010 620.840 19.310 ;
        RECT 401.220 17.690 401.480 18.010 ;
        RECT 620.640 17.690 620.900 18.010 ;
        RECT 401.280 2.400 401.420 17.690 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 621.550 917.520 621.830 917.800 ;
        RECT 622.930 917.520 623.210 917.800 ;
      LAYER met3 ;
        RECT 621.525 917.810 621.855 917.825 ;
        RECT 622.905 917.810 623.235 917.825 ;
        RECT 621.525 917.510 623.235 917.810 ;
        RECT 621.525 917.495 621.855 917.510 ;
        RECT 622.905 917.495 623.235 917.510 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 345.605 1497.445 345.775 1545.555 ;
        RECT 345.605 1352.605 345.775 1400.715 ;
        RECT 345.605 1256.045 345.775 1304.155 ;
        RECT 345.605 338.045 345.775 386.155 ;
        RECT 345.605 241.485 345.775 289.595 ;
        RECT 345.605 144.925 345.775 193.035 ;
      LAYER mcon ;
        RECT 345.605 1545.385 345.775 1545.555 ;
        RECT 345.605 1400.545 345.775 1400.715 ;
        RECT 345.605 1303.985 345.775 1304.155 ;
        RECT 345.605 385.985 345.775 386.155 ;
        RECT 345.605 289.425 345.775 289.595 ;
        RECT 345.605 192.865 345.775 193.035 ;
      LAYER met1 ;
        RECT 345.545 1545.540 345.835 1545.585 ;
        RECT 345.990 1545.540 346.310 1545.600 ;
        RECT 345.545 1545.400 346.310 1545.540 ;
        RECT 345.545 1545.355 345.835 1545.400 ;
        RECT 345.990 1545.340 346.310 1545.400 ;
        RECT 345.530 1497.600 345.850 1497.660 ;
        RECT 345.335 1497.460 345.850 1497.600 ;
        RECT 345.530 1497.400 345.850 1497.460 ;
        RECT 345.530 1400.700 345.850 1400.760 ;
        RECT 345.335 1400.560 345.850 1400.700 ;
        RECT 345.530 1400.500 345.850 1400.560 ;
        RECT 345.545 1352.760 345.835 1352.805 ;
        RECT 345.990 1352.760 346.310 1352.820 ;
        RECT 345.545 1352.620 346.310 1352.760 ;
        RECT 345.545 1352.575 345.835 1352.620 ;
        RECT 345.990 1352.560 346.310 1352.620 ;
        RECT 345.530 1304.140 345.850 1304.200 ;
        RECT 345.335 1304.000 345.850 1304.140 ;
        RECT 345.530 1303.940 345.850 1304.000 ;
        RECT 345.545 1256.200 345.835 1256.245 ;
        RECT 345.990 1256.200 346.310 1256.260 ;
        RECT 345.545 1256.060 346.310 1256.200 ;
        RECT 345.545 1256.015 345.835 1256.060 ;
        RECT 345.990 1256.000 346.310 1256.060 ;
        RECT 345.990 1159.300 346.310 1159.360 ;
        RECT 346.910 1159.300 347.230 1159.360 ;
        RECT 345.990 1159.160 347.230 1159.300 ;
        RECT 345.990 1159.100 346.310 1159.160 ;
        RECT 346.910 1159.100 347.230 1159.160 ;
        RECT 345.990 1062.740 346.310 1062.800 ;
        RECT 346.910 1062.740 347.230 1062.800 ;
        RECT 345.990 1062.600 347.230 1062.740 ;
        RECT 345.990 1062.540 346.310 1062.600 ;
        RECT 346.910 1062.540 347.230 1062.600 ;
        RECT 345.990 966.180 346.310 966.240 ;
        RECT 346.910 966.180 347.230 966.240 ;
        RECT 345.990 966.040 347.230 966.180 ;
        RECT 345.990 965.980 346.310 966.040 ;
        RECT 346.910 965.980 347.230 966.040 ;
        RECT 345.990 869.620 346.310 869.680 ;
        RECT 346.910 869.620 347.230 869.680 ;
        RECT 345.990 869.480 347.230 869.620 ;
        RECT 345.990 869.420 346.310 869.480 ;
        RECT 346.910 869.420 347.230 869.480 ;
        RECT 345.530 821.000 345.850 821.060 ;
        RECT 346.910 821.000 347.230 821.060 ;
        RECT 345.530 820.860 347.230 821.000 ;
        RECT 345.530 820.800 345.850 820.860 ;
        RECT 346.910 820.800 347.230 820.860 ;
        RECT 345.530 689.900 345.850 690.160 ;
        RECT 345.070 689.760 345.390 689.820 ;
        RECT 345.620 689.760 345.760 689.900 ;
        RECT 345.070 689.620 345.760 689.760 ;
        RECT 345.070 689.560 345.390 689.620 ;
        RECT 345.530 593.340 345.850 593.600 ;
        RECT 345.070 593.200 345.390 593.260 ;
        RECT 345.620 593.200 345.760 593.340 ;
        RECT 345.070 593.060 345.760 593.200 ;
        RECT 345.070 593.000 345.390 593.060 ;
        RECT 345.530 496.780 345.850 497.040 ;
        RECT 345.070 496.640 345.390 496.700 ;
        RECT 345.620 496.640 345.760 496.780 ;
        RECT 345.070 496.500 345.760 496.640 ;
        RECT 345.070 496.440 345.390 496.500 ;
        RECT 345.530 400.220 345.850 400.480 ;
        RECT 345.620 400.080 345.760 400.220 ;
        RECT 345.990 400.080 346.310 400.140 ;
        RECT 345.620 399.940 346.310 400.080 ;
        RECT 345.990 399.880 346.310 399.940 ;
        RECT 345.545 386.140 345.835 386.185 ;
        RECT 345.990 386.140 346.310 386.200 ;
        RECT 345.545 386.000 346.310 386.140 ;
        RECT 345.545 385.955 345.835 386.000 ;
        RECT 345.990 385.940 346.310 386.000 ;
        RECT 345.530 338.200 345.850 338.260 ;
        RECT 345.335 338.060 345.850 338.200 ;
        RECT 345.530 338.000 345.850 338.060 ;
        RECT 344.150 303.520 344.470 303.580 ;
        RECT 345.990 303.520 346.310 303.580 ;
        RECT 344.150 303.380 346.310 303.520 ;
        RECT 344.150 303.320 344.470 303.380 ;
        RECT 345.990 303.320 346.310 303.380 ;
        RECT 345.545 289.580 345.835 289.625 ;
        RECT 345.990 289.580 346.310 289.640 ;
        RECT 345.545 289.440 346.310 289.580 ;
        RECT 345.545 289.395 345.835 289.440 ;
        RECT 345.990 289.380 346.310 289.440 ;
        RECT 345.530 241.640 345.850 241.700 ;
        RECT 345.335 241.500 345.850 241.640 ;
        RECT 345.530 241.440 345.850 241.500 ;
        RECT 345.070 206.960 345.390 207.020 ;
        RECT 345.990 206.960 346.310 207.020 ;
        RECT 345.070 206.820 346.310 206.960 ;
        RECT 345.070 206.760 345.390 206.820 ;
        RECT 345.990 206.760 346.310 206.820 ;
        RECT 345.545 193.020 345.835 193.065 ;
        RECT 345.990 193.020 346.310 193.080 ;
        RECT 345.545 192.880 346.310 193.020 ;
        RECT 345.545 192.835 345.835 192.880 ;
        RECT 345.990 192.820 346.310 192.880 ;
        RECT 345.530 145.080 345.850 145.140 ;
        RECT 345.335 144.940 345.850 145.080 ;
        RECT 345.530 144.880 345.850 144.940 ;
        RECT 62.170 25.400 62.490 25.460 ;
        RECT 345.990 25.400 346.310 25.460 ;
        RECT 62.170 25.260 346.310 25.400 ;
        RECT 62.170 25.200 62.490 25.260 ;
        RECT 345.990 25.200 346.310 25.260 ;
      LAYER via ;
        RECT 346.020 1545.340 346.280 1545.600 ;
        RECT 345.560 1497.400 345.820 1497.660 ;
        RECT 345.560 1400.500 345.820 1400.760 ;
        RECT 346.020 1352.560 346.280 1352.820 ;
        RECT 345.560 1303.940 345.820 1304.200 ;
        RECT 346.020 1256.000 346.280 1256.260 ;
        RECT 346.020 1159.100 346.280 1159.360 ;
        RECT 346.940 1159.100 347.200 1159.360 ;
        RECT 346.020 1062.540 346.280 1062.800 ;
        RECT 346.940 1062.540 347.200 1062.800 ;
        RECT 346.020 965.980 346.280 966.240 ;
        RECT 346.940 965.980 347.200 966.240 ;
        RECT 346.020 869.420 346.280 869.680 ;
        RECT 346.940 869.420 347.200 869.680 ;
        RECT 345.560 820.800 345.820 821.060 ;
        RECT 346.940 820.800 347.200 821.060 ;
        RECT 345.560 689.900 345.820 690.160 ;
        RECT 345.100 689.560 345.360 689.820 ;
        RECT 345.560 593.340 345.820 593.600 ;
        RECT 345.100 593.000 345.360 593.260 ;
        RECT 345.560 496.780 345.820 497.040 ;
        RECT 345.100 496.440 345.360 496.700 ;
        RECT 345.560 400.220 345.820 400.480 ;
        RECT 346.020 399.880 346.280 400.140 ;
        RECT 346.020 385.940 346.280 386.200 ;
        RECT 345.560 338.000 345.820 338.260 ;
        RECT 344.180 303.320 344.440 303.580 ;
        RECT 346.020 303.320 346.280 303.580 ;
        RECT 346.020 289.380 346.280 289.640 ;
        RECT 345.560 241.440 345.820 241.700 ;
        RECT 345.100 206.760 345.360 207.020 ;
        RECT 346.020 206.760 346.280 207.020 ;
        RECT 346.020 192.820 346.280 193.080 ;
        RECT 345.560 144.880 345.820 145.140 ;
        RECT 62.200 25.200 62.460 25.460 ;
        RECT 346.020 25.200 346.280 25.460 ;
      LAYER met2 ;
        RECT 350.620 1601.130 350.900 1604.000 ;
        RECT 346.080 1600.990 350.900 1601.130 ;
        RECT 346.080 1545.630 346.220 1600.990 ;
        RECT 350.620 1600.000 350.900 1600.990 ;
        RECT 346.020 1545.310 346.280 1545.630 ;
        RECT 345.560 1497.370 345.820 1497.690 ;
        RECT 345.620 1473.290 345.760 1497.370 ;
        RECT 345.620 1473.150 346.220 1473.290 ;
        RECT 346.080 1414.130 346.220 1473.150 ;
        RECT 345.620 1413.990 346.220 1414.130 ;
        RECT 345.620 1400.790 345.760 1413.990 ;
        RECT 345.560 1400.470 345.820 1400.790 ;
        RECT 346.020 1352.530 346.280 1352.850 ;
        RECT 346.080 1317.570 346.220 1352.530 ;
        RECT 345.620 1317.430 346.220 1317.570 ;
        RECT 345.620 1304.230 345.760 1317.430 ;
        RECT 345.560 1303.910 345.820 1304.230 ;
        RECT 346.020 1255.970 346.280 1256.290 ;
        RECT 346.080 1221.010 346.220 1255.970 ;
        RECT 345.620 1220.870 346.220 1221.010 ;
        RECT 345.620 1207.525 345.760 1220.870 ;
        RECT 345.550 1207.155 345.830 1207.525 ;
        RECT 346.930 1207.155 347.210 1207.525 ;
        RECT 347.000 1159.390 347.140 1207.155 ;
        RECT 346.020 1159.070 346.280 1159.390 ;
        RECT 346.940 1159.070 347.200 1159.390 ;
        RECT 346.080 1124.450 346.220 1159.070 ;
        RECT 345.620 1124.310 346.220 1124.450 ;
        RECT 345.620 1110.965 345.760 1124.310 ;
        RECT 345.550 1110.595 345.830 1110.965 ;
        RECT 346.930 1110.595 347.210 1110.965 ;
        RECT 347.000 1062.830 347.140 1110.595 ;
        RECT 346.020 1062.510 346.280 1062.830 ;
        RECT 346.940 1062.510 347.200 1062.830 ;
        RECT 346.080 1027.890 346.220 1062.510 ;
        RECT 345.620 1027.750 346.220 1027.890 ;
        RECT 345.620 1014.405 345.760 1027.750 ;
        RECT 345.550 1014.035 345.830 1014.405 ;
        RECT 346.930 1014.035 347.210 1014.405 ;
        RECT 347.000 966.270 347.140 1014.035 ;
        RECT 346.020 965.950 346.280 966.270 ;
        RECT 346.940 965.950 347.200 966.270 ;
        RECT 346.080 931.330 346.220 965.950 ;
        RECT 345.620 931.190 346.220 931.330 ;
        RECT 345.620 917.845 345.760 931.190 ;
        RECT 345.550 917.475 345.830 917.845 ;
        RECT 346.930 917.475 347.210 917.845 ;
        RECT 347.000 869.710 347.140 917.475 ;
        RECT 346.020 869.390 346.280 869.710 ;
        RECT 346.940 869.390 347.200 869.710 ;
        RECT 346.080 834.770 346.220 869.390 ;
        RECT 345.620 834.630 346.220 834.770 ;
        RECT 345.620 821.090 345.760 834.630 ;
        RECT 345.560 820.770 345.820 821.090 ;
        RECT 346.940 820.770 347.200 821.090 ;
        RECT 347.000 773.005 347.140 820.770 ;
        RECT 346.010 772.635 346.290 773.005 ;
        RECT 346.930 772.635 347.210 773.005 ;
        RECT 346.080 738.210 346.220 772.635 ;
        RECT 345.620 738.070 346.220 738.210 ;
        RECT 345.620 690.190 345.760 738.070 ;
        RECT 345.560 689.870 345.820 690.190 ;
        RECT 345.100 689.530 345.360 689.850 ;
        RECT 345.160 676.445 345.300 689.530 ;
        RECT 345.090 676.075 345.370 676.445 ;
        RECT 346.010 676.075 346.290 676.445 ;
        RECT 346.080 641.650 346.220 676.075 ;
        RECT 345.620 641.510 346.220 641.650 ;
        RECT 345.620 593.630 345.760 641.510 ;
        RECT 345.560 593.310 345.820 593.630 ;
        RECT 345.100 592.970 345.360 593.290 ;
        RECT 345.160 579.885 345.300 592.970 ;
        RECT 345.090 579.515 345.370 579.885 ;
        RECT 346.010 579.515 346.290 579.885 ;
        RECT 346.080 545.090 346.220 579.515 ;
        RECT 345.620 544.950 346.220 545.090 ;
        RECT 345.620 497.070 345.760 544.950 ;
        RECT 345.560 496.750 345.820 497.070 ;
        RECT 345.100 496.410 345.360 496.730 ;
        RECT 345.160 483.325 345.300 496.410 ;
        RECT 345.090 482.955 345.370 483.325 ;
        RECT 346.010 482.955 346.290 483.325 ;
        RECT 346.080 448.530 346.220 482.955 ;
        RECT 345.620 448.390 346.220 448.530 ;
        RECT 345.620 400.510 345.760 448.390 ;
        RECT 345.560 400.190 345.820 400.510 ;
        RECT 346.020 399.850 346.280 400.170 ;
        RECT 346.080 386.230 346.220 399.850 ;
        RECT 346.020 385.910 346.280 386.230 ;
        RECT 345.560 337.970 345.820 338.290 ;
        RECT 344.170 337.435 344.450 337.805 ;
        RECT 345.090 337.690 345.370 337.805 ;
        RECT 345.620 337.690 345.760 337.970 ;
        RECT 345.090 337.550 345.760 337.690 ;
        RECT 345.090 337.435 345.370 337.550 ;
        RECT 344.240 303.610 344.380 337.435 ;
        RECT 344.180 303.290 344.440 303.610 ;
        RECT 346.020 303.290 346.280 303.610 ;
        RECT 346.080 289.670 346.220 303.290 ;
        RECT 346.020 289.350 346.280 289.670 ;
        RECT 345.560 241.410 345.820 241.730 ;
        RECT 345.620 207.130 345.760 241.410 ;
        RECT 345.160 207.050 345.760 207.130 ;
        RECT 345.100 206.990 345.760 207.050 ;
        RECT 345.100 206.730 345.360 206.990 ;
        RECT 346.020 206.730 346.280 207.050 ;
        RECT 346.080 193.110 346.220 206.730 ;
        RECT 346.020 192.790 346.280 193.110 ;
        RECT 345.560 144.850 345.820 145.170 ;
        RECT 345.620 120.770 345.760 144.850 ;
        RECT 345.620 120.630 346.220 120.770 ;
        RECT 346.080 25.490 346.220 120.630 ;
        RECT 62.200 25.170 62.460 25.490 ;
        RECT 346.020 25.170 346.280 25.490 ;
        RECT 62.260 2.400 62.400 25.170 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 345.550 1207.200 345.830 1207.480 ;
        RECT 346.930 1207.200 347.210 1207.480 ;
        RECT 345.550 1110.640 345.830 1110.920 ;
        RECT 346.930 1110.640 347.210 1110.920 ;
        RECT 345.550 1014.080 345.830 1014.360 ;
        RECT 346.930 1014.080 347.210 1014.360 ;
        RECT 345.550 917.520 345.830 917.800 ;
        RECT 346.930 917.520 347.210 917.800 ;
        RECT 346.010 772.680 346.290 772.960 ;
        RECT 346.930 772.680 347.210 772.960 ;
        RECT 345.090 676.120 345.370 676.400 ;
        RECT 346.010 676.120 346.290 676.400 ;
        RECT 345.090 579.560 345.370 579.840 ;
        RECT 346.010 579.560 346.290 579.840 ;
        RECT 345.090 483.000 345.370 483.280 ;
        RECT 346.010 483.000 346.290 483.280 ;
        RECT 344.170 337.480 344.450 337.760 ;
        RECT 345.090 337.480 345.370 337.760 ;
      LAYER met3 ;
        RECT 345.525 1207.490 345.855 1207.505 ;
        RECT 346.905 1207.490 347.235 1207.505 ;
        RECT 345.525 1207.190 347.235 1207.490 ;
        RECT 345.525 1207.175 345.855 1207.190 ;
        RECT 346.905 1207.175 347.235 1207.190 ;
        RECT 345.525 1110.930 345.855 1110.945 ;
        RECT 346.905 1110.930 347.235 1110.945 ;
        RECT 345.525 1110.630 347.235 1110.930 ;
        RECT 345.525 1110.615 345.855 1110.630 ;
        RECT 346.905 1110.615 347.235 1110.630 ;
        RECT 345.525 1014.370 345.855 1014.385 ;
        RECT 346.905 1014.370 347.235 1014.385 ;
        RECT 345.525 1014.070 347.235 1014.370 ;
        RECT 345.525 1014.055 345.855 1014.070 ;
        RECT 346.905 1014.055 347.235 1014.070 ;
        RECT 345.525 917.810 345.855 917.825 ;
        RECT 346.905 917.810 347.235 917.825 ;
        RECT 345.525 917.510 347.235 917.810 ;
        RECT 345.525 917.495 345.855 917.510 ;
        RECT 346.905 917.495 347.235 917.510 ;
        RECT 345.985 772.970 346.315 772.985 ;
        RECT 346.905 772.970 347.235 772.985 ;
        RECT 345.985 772.670 347.235 772.970 ;
        RECT 345.985 772.655 346.315 772.670 ;
        RECT 346.905 772.655 347.235 772.670 ;
        RECT 345.065 676.410 345.395 676.425 ;
        RECT 345.985 676.410 346.315 676.425 ;
        RECT 345.065 676.110 346.315 676.410 ;
        RECT 345.065 676.095 345.395 676.110 ;
        RECT 345.985 676.095 346.315 676.110 ;
        RECT 345.065 579.850 345.395 579.865 ;
        RECT 345.985 579.850 346.315 579.865 ;
        RECT 345.065 579.550 346.315 579.850 ;
        RECT 345.065 579.535 345.395 579.550 ;
        RECT 345.985 579.535 346.315 579.550 ;
        RECT 345.065 483.290 345.395 483.305 ;
        RECT 345.985 483.290 346.315 483.305 ;
        RECT 345.065 482.990 346.315 483.290 ;
        RECT 345.065 482.975 345.395 482.990 ;
        RECT 345.985 482.975 346.315 482.990 ;
        RECT 344.145 337.770 344.475 337.785 ;
        RECT 345.065 337.770 345.395 337.785 ;
        RECT 344.145 337.470 345.395 337.770 ;
        RECT 344.145 337.455 344.475 337.470 ;
        RECT 345.065 337.455 345.395 337.470 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 635.405 1497.445 635.575 1545.555 ;
        RECT 635.405 1459.365 635.575 1463.275 ;
        RECT 635.405 786.505 635.575 821.015 ;
        RECT 635.405 689.605 635.575 724.455 ;
        RECT 635.405 593.045 635.575 627.895 ;
        RECT 635.405 496.485 635.575 531.335 ;
        RECT 635.405 386.325 635.575 434.775 ;
        RECT 635.405 241.485 635.575 289.595 ;
        RECT 635.405 144.925 635.575 193.035 ;
      LAYER mcon ;
        RECT 635.405 1545.385 635.575 1545.555 ;
        RECT 635.405 1463.105 635.575 1463.275 ;
        RECT 635.405 820.845 635.575 821.015 ;
        RECT 635.405 724.285 635.575 724.455 ;
        RECT 635.405 627.725 635.575 627.895 ;
        RECT 635.405 531.165 635.575 531.335 ;
        RECT 635.405 434.605 635.575 434.775 ;
        RECT 635.405 289.425 635.575 289.595 ;
        RECT 635.405 192.865 635.575 193.035 ;
      LAYER met1 ;
        RECT 634.870 1559.140 635.190 1559.200 ;
        RECT 635.790 1559.140 636.110 1559.200 ;
        RECT 634.870 1559.000 636.110 1559.140 ;
        RECT 634.870 1558.940 635.190 1559.000 ;
        RECT 635.790 1558.940 636.110 1559.000 ;
        RECT 635.345 1545.540 635.635 1545.585 ;
        RECT 635.790 1545.540 636.110 1545.600 ;
        RECT 635.345 1545.400 636.110 1545.540 ;
        RECT 635.345 1545.355 635.635 1545.400 ;
        RECT 635.790 1545.340 636.110 1545.400 ;
        RECT 635.330 1497.600 635.650 1497.660 ;
        RECT 635.135 1497.460 635.650 1497.600 ;
        RECT 635.330 1497.400 635.650 1497.460 ;
        RECT 635.330 1463.260 635.650 1463.320 ;
        RECT 635.135 1463.120 635.650 1463.260 ;
        RECT 635.330 1463.060 635.650 1463.120 ;
        RECT 635.330 1459.520 635.650 1459.580 ;
        RECT 635.135 1459.380 635.650 1459.520 ;
        RECT 635.330 1459.320 635.650 1459.380 ;
        RECT 634.870 1318.080 635.190 1318.140 ;
        RECT 635.790 1318.080 636.110 1318.140 ;
        RECT 634.870 1317.940 636.110 1318.080 ;
        RECT 634.870 1317.880 635.190 1317.940 ;
        RECT 635.790 1317.880 636.110 1317.940 ;
        RECT 634.870 1221.520 635.190 1221.580 ;
        RECT 635.790 1221.520 636.110 1221.580 ;
        RECT 634.870 1221.380 636.110 1221.520 ;
        RECT 634.870 1221.320 635.190 1221.380 ;
        RECT 635.790 1221.320 636.110 1221.380 ;
        RECT 634.870 1124.960 635.190 1125.020 ;
        RECT 635.790 1124.960 636.110 1125.020 ;
        RECT 634.870 1124.820 636.110 1124.960 ;
        RECT 634.870 1124.760 635.190 1124.820 ;
        RECT 635.790 1124.760 636.110 1124.820 ;
        RECT 634.870 1028.400 635.190 1028.460 ;
        RECT 635.790 1028.400 636.110 1028.460 ;
        RECT 634.870 1028.260 636.110 1028.400 ;
        RECT 634.870 1028.200 635.190 1028.260 ;
        RECT 635.790 1028.200 636.110 1028.260 ;
        RECT 634.870 931.840 635.190 931.900 ;
        RECT 635.790 931.840 636.110 931.900 ;
        RECT 634.870 931.700 636.110 931.840 ;
        RECT 634.870 931.640 635.190 931.700 ;
        RECT 635.790 931.640 636.110 931.700 ;
        RECT 634.410 869.620 634.730 869.680 ;
        RECT 635.790 869.620 636.110 869.680 ;
        RECT 634.410 869.480 636.110 869.620 ;
        RECT 634.410 869.420 634.730 869.480 ;
        RECT 635.790 869.420 636.110 869.480 ;
        RECT 634.870 835.280 635.190 835.340 ;
        RECT 635.790 835.280 636.110 835.340 ;
        RECT 634.870 835.140 636.110 835.280 ;
        RECT 634.870 835.080 635.190 835.140 ;
        RECT 635.790 835.080 636.110 835.140 ;
        RECT 635.330 821.000 635.650 821.060 ;
        RECT 635.135 820.860 635.650 821.000 ;
        RECT 635.330 820.800 635.650 820.860 ;
        RECT 635.330 786.660 635.650 786.720 ;
        RECT 635.135 786.520 635.650 786.660 ;
        RECT 635.330 786.460 635.650 786.520 ;
        RECT 634.870 738.380 635.190 738.440 ;
        RECT 635.790 738.380 636.110 738.440 ;
        RECT 634.870 738.240 636.110 738.380 ;
        RECT 634.870 738.180 635.190 738.240 ;
        RECT 635.790 738.180 636.110 738.240 ;
        RECT 635.330 724.440 635.650 724.500 ;
        RECT 635.135 724.300 635.650 724.440 ;
        RECT 635.330 724.240 635.650 724.300 ;
        RECT 635.330 689.760 635.650 689.820 ;
        RECT 635.135 689.620 635.650 689.760 ;
        RECT 635.330 689.560 635.650 689.620 ;
        RECT 634.870 641.820 635.190 641.880 ;
        RECT 635.790 641.820 636.110 641.880 ;
        RECT 634.870 641.680 636.110 641.820 ;
        RECT 634.870 641.620 635.190 641.680 ;
        RECT 635.790 641.620 636.110 641.680 ;
        RECT 635.330 627.880 635.650 627.940 ;
        RECT 635.135 627.740 635.650 627.880 ;
        RECT 635.330 627.680 635.650 627.740 ;
        RECT 635.330 593.200 635.650 593.260 ;
        RECT 635.135 593.060 635.650 593.200 ;
        RECT 635.330 593.000 635.650 593.060 ;
        RECT 634.870 545.260 635.190 545.320 ;
        RECT 635.790 545.260 636.110 545.320 ;
        RECT 634.870 545.120 636.110 545.260 ;
        RECT 634.870 545.060 635.190 545.120 ;
        RECT 635.790 545.060 636.110 545.120 ;
        RECT 635.330 531.320 635.650 531.380 ;
        RECT 635.135 531.180 635.650 531.320 ;
        RECT 635.330 531.120 635.650 531.180 ;
        RECT 635.330 496.640 635.650 496.700 ;
        RECT 635.135 496.500 635.650 496.640 ;
        RECT 635.330 496.440 635.650 496.500 ;
        RECT 634.870 448.700 635.190 448.760 ;
        RECT 635.790 448.700 636.110 448.760 ;
        RECT 634.870 448.560 636.110 448.700 ;
        RECT 634.870 448.500 635.190 448.560 ;
        RECT 635.790 448.500 636.110 448.560 ;
        RECT 635.330 434.760 635.650 434.820 ;
        RECT 635.135 434.620 635.650 434.760 ;
        RECT 635.330 434.560 635.650 434.620 ;
        RECT 635.345 386.480 635.635 386.525 ;
        RECT 635.790 386.480 636.110 386.540 ;
        RECT 635.345 386.340 636.110 386.480 ;
        RECT 635.345 386.295 635.635 386.340 ;
        RECT 635.790 386.280 636.110 386.340 ;
        RECT 634.870 352.140 635.190 352.200 ;
        RECT 634.870 352.000 635.560 352.140 ;
        RECT 634.870 351.940 635.190 352.000 ;
        RECT 635.420 351.860 635.560 352.000 ;
        RECT 635.330 351.600 635.650 351.860 ;
        RECT 635.345 289.580 635.635 289.625 ;
        RECT 635.790 289.580 636.110 289.640 ;
        RECT 635.345 289.440 636.110 289.580 ;
        RECT 635.345 289.395 635.635 289.440 ;
        RECT 635.790 289.380 636.110 289.440 ;
        RECT 635.330 241.640 635.650 241.700 ;
        RECT 635.135 241.500 635.650 241.640 ;
        RECT 635.330 241.440 635.650 241.500 ;
        RECT 635.345 193.020 635.635 193.065 ;
        RECT 635.790 193.020 636.110 193.080 ;
        RECT 635.345 192.880 636.110 193.020 ;
        RECT 635.345 192.835 635.635 192.880 ;
        RECT 635.790 192.820 636.110 192.880 ;
        RECT 635.330 145.080 635.650 145.140 ;
        RECT 635.135 144.940 635.650 145.080 ;
        RECT 635.330 144.880 635.650 144.940 ;
        RECT 419.130 17.240 419.450 17.300 ;
        RECT 634.870 17.240 635.190 17.300 ;
        RECT 419.130 17.100 635.190 17.240 ;
        RECT 419.130 17.040 419.450 17.100 ;
        RECT 634.870 17.040 635.190 17.100 ;
      LAYER via ;
        RECT 634.900 1558.940 635.160 1559.200 ;
        RECT 635.820 1558.940 636.080 1559.200 ;
        RECT 635.820 1545.340 636.080 1545.600 ;
        RECT 635.360 1497.400 635.620 1497.660 ;
        RECT 635.360 1463.060 635.620 1463.320 ;
        RECT 635.360 1459.320 635.620 1459.580 ;
        RECT 634.900 1317.880 635.160 1318.140 ;
        RECT 635.820 1317.880 636.080 1318.140 ;
        RECT 634.900 1221.320 635.160 1221.580 ;
        RECT 635.820 1221.320 636.080 1221.580 ;
        RECT 634.900 1124.760 635.160 1125.020 ;
        RECT 635.820 1124.760 636.080 1125.020 ;
        RECT 634.900 1028.200 635.160 1028.460 ;
        RECT 635.820 1028.200 636.080 1028.460 ;
        RECT 634.900 931.640 635.160 931.900 ;
        RECT 635.820 931.640 636.080 931.900 ;
        RECT 634.440 869.420 634.700 869.680 ;
        RECT 635.820 869.420 636.080 869.680 ;
        RECT 634.900 835.080 635.160 835.340 ;
        RECT 635.820 835.080 636.080 835.340 ;
        RECT 635.360 820.800 635.620 821.060 ;
        RECT 635.360 786.460 635.620 786.720 ;
        RECT 634.900 738.180 635.160 738.440 ;
        RECT 635.820 738.180 636.080 738.440 ;
        RECT 635.360 724.240 635.620 724.500 ;
        RECT 635.360 689.560 635.620 689.820 ;
        RECT 634.900 641.620 635.160 641.880 ;
        RECT 635.820 641.620 636.080 641.880 ;
        RECT 635.360 627.680 635.620 627.940 ;
        RECT 635.360 593.000 635.620 593.260 ;
        RECT 634.900 545.060 635.160 545.320 ;
        RECT 635.820 545.060 636.080 545.320 ;
        RECT 635.360 531.120 635.620 531.380 ;
        RECT 635.360 496.440 635.620 496.700 ;
        RECT 634.900 448.500 635.160 448.760 ;
        RECT 635.820 448.500 636.080 448.760 ;
        RECT 635.360 434.560 635.620 434.820 ;
        RECT 635.820 386.280 636.080 386.540 ;
        RECT 634.900 351.940 635.160 352.200 ;
        RECT 635.360 351.600 635.620 351.860 ;
        RECT 635.820 289.380 636.080 289.640 ;
        RECT 635.360 241.440 635.620 241.700 ;
        RECT 635.820 192.820 636.080 193.080 ;
        RECT 635.360 144.880 635.620 145.140 ;
        RECT 419.160 17.040 419.420 17.300 ;
        RECT 634.900 17.040 635.160 17.300 ;
      LAYER met2 ;
        RECT 641.340 1601.130 641.620 1604.000 ;
        RECT 636.800 1600.990 641.620 1601.130 ;
        RECT 636.800 1580.050 636.940 1600.990 ;
        RECT 641.340 1600.000 641.620 1600.990 ;
        RECT 634.960 1579.910 636.940 1580.050 ;
        RECT 634.960 1559.230 635.100 1579.910 ;
        RECT 634.900 1558.910 635.160 1559.230 ;
        RECT 635.820 1558.910 636.080 1559.230 ;
        RECT 635.880 1545.630 636.020 1558.910 ;
        RECT 635.820 1545.310 636.080 1545.630 ;
        RECT 635.360 1497.370 635.620 1497.690 ;
        RECT 635.420 1463.350 635.560 1497.370 ;
        RECT 635.360 1463.030 635.620 1463.350 ;
        RECT 635.360 1459.290 635.620 1459.610 ;
        RECT 635.420 1414.810 635.560 1459.290 ;
        RECT 635.420 1414.670 636.020 1414.810 ;
        RECT 635.880 1318.170 636.020 1414.670 ;
        RECT 634.900 1317.850 635.160 1318.170 ;
        RECT 635.820 1317.850 636.080 1318.170 ;
        RECT 634.960 1317.570 635.100 1317.850 ;
        RECT 634.960 1317.430 635.560 1317.570 ;
        RECT 635.420 1269.970 635.560 1317.430 ;
        RECT 635.420 1269.830 636.020 1269.970 ;
        RECT 635.880 1221.610 636.020 1269.830 ;
        RECT 634.900 1221.290 635.160 1221.610 ;
        RECT 635.820 1221.290 636.080 1221.610 ;
        RECT 634.960 1221.010 635.100 1221.290 ;
        RECT 634.960 1220.870 635.560 1221.010 ;
        RECT 635.420 1173.410 635.560 1220.870 ;
        RECT 635.420 1173.270 636.020 1173.410 ;
        RECT 635.880 1125.050 636.020 1173.270 ;
        RECT 634.900 1124.730 635.160 1125.050 ;
        RECT 635.820 1124.730 636.080 1125.050 ;
        RECT 634.960 1124.450 635.100 1124.730 ;
        RECT 634.960 1124.310 635.560 1124.450 ;
        RECT 635.420 1076.850 635.560 1124.310 ;
        RECT 635.420 1076.710 636.020 1076.850 ;
        RECT 635.880 1028.490 636.020 1076.710 ;
        RECT 634.900 1028.170 635.160 1028.490 ;
        RECT 635.820 1028.170 636.080 1028.490 ;
        RECT 634.960 1027.890 635.100 1028.170 ;
        RECT 634.960 1027.750 635.560 1027.890 ;
        RECT 635.420 980.290 635.560 1027.750 ;
        RECT 635.420 980.150 636.020 980.290 ;
        RECT 635.880 931.930 636.020 980.150 ;
        RECT 634.900 931.610 635.160 931.930 ;
        RECT 635.820 931.610 636.080 931.930 ;
        RECT 634.960 931.330 635.100 931.610 ;
        RECT 634.960 931.190 635.560 931.330 ;
        RECT 635.420 917.845 635.560 931.190 ;
        RECT 634.430 917.475 634.710 917.845 ;
        RECT 635.350 917.475 635.630 917.845 ;
        RECT 634.500 869.710 634.640 917.475 ;
        RECT 634.440 869.390 634.700 869.710 ;
        RECT 635.820 869.390 636.080 869.710 ;
        RECT 635.880 835.370 636.020 869.390 ;
        RECT 634.900 835.050 635.160 835.370 ;
        RECT 635.820 835.050 636.080 835.370 ;
        RECT 634.960 834.770 635.100 835.050 ;
        RECT 634.960 834.630 635.560 834.770 ;
        RECT 635.420 821.090 635.560 834.630 ;
        RECT 635.360 820.770 635.620 821.090 ;
        RECT 635.360 786.430 635.620 786.750 ;
        RECT 635.420 772.890 635.560 786.430 ;
        RECT 635.420 772.750 636.020 772.890 ;
        RECT 635.880 738.470 636.020 772.750 ;
        RECT 634.900 738.210 635.160 738.470 ;
        RECT 634.900 738.150 635.560 738.210 ;
        RECT 635.820 738.150 636.080 738.470 ;
        RECT 634.960 738.070 635.560 738.150 ;
        RECT 635.420 724.530 635.560 738.070 ;
        RECT 635.360 724.210 635.620 724.530 ;
        RECT 635.360 689.530 635.620 689.850 ;
        RECT 635.420 676.330 635.560 689.530 ;
        RECT 635.420 676.190 636.020 676.330 ;
        RECT 635.880 641.910 636.020 676.190 ;
        RECT 634.900 641.650 635.160 641.910 ;
        RECT 634.900 641.590 635.560 641.650 ;
        RECT 635.820 641.590 636.080 641.910 ;
        RECT 634.960 641.510 635.560 641.590 ;
        RECT 635.420 627.970 635.560 641.510 ;
        RECT 635.360 627.650 635.620 627.970 ;
        RECT 635.360 592.970 635.620 593.290 ;
        RECT 635.420 579.770 635.560 592.970 ;
        RECT 635.420 579.630 636.020 579.770 ;
        RECT 635.880 545.350 636.020 579.630 ;
        RECT 634.900 545.090 635.160 545.350 ;
        RECT 634.900 545.030 635.560 545.090 ;
        RECT 635.820 545.030 636.080 545.350 ;
        RECT 634.960 544.950 635.560 545.030 ;
        RECT 635.420 531.410 635.560 544.950 ;
        RECT 635.360 531.090 635.620 531.410 ;
        RECT 635.360 496.410 635.620 496.730 ;
        RECT 635.420 483.210 635.560 496.410 ;
        RECT 635.420 483.070 636.020 483.210 ;
        RECT 635.880 448.790 636.020 483.070 ;
        RECT 634.900 448.530 635.160 448.790 ;
        RECT 634.900 448.470 635.560 448.530 ;
        RECT 635.820 448.470 636.080 448.790 ;
        RECT 634.960 448.390 635.560 448.470 ;
        RECT 635.420 434.850 635.560 448.390 ;
        RECT 635.360 434.530 635.620 434.850 ;
        RECT 635.820 386.250 636.080 386.570 ;
        RECT 635.880 386.085 636.020 386.250 ;
        RECT 634.890 385.715 635.170 386.085 ;
        RECT 635.810 385.715 636.090 386.085 ;
        RECT 634.960 352.230 635.100 385.715 ;
        RECT 634.900 351.910 635.160 352.230 ;
        RECT 635.360 351.570 635.620 351.890 ;
        RECT 635.420 303.690 635.560 351.570 ;
        RECT 635.420 303.550 636.020 303.690 ;
        RECT 635.880 289.670 636.020 303.550 ;
        RECT 635.820 289.350 636.080 289.670 ;
        RECT 635.360 241.410 635.620 241.730 ;
        RECT 635.420 207.130 635.560 241.410 ;
        RECT 635.420 206.990 636.020 207.130 ;
        RECT 635.880 193.110 636.020 206.990 ;
        RECT 635.820 192.790 636.080 193.110 ;
        RECT 635.360 144.850 635.620 145.170 ;
        RECT 635.420 110.570 635.560 144.850 ;
        RECT 635.420 110.430 636.020 110.570 ;
        RECT 635.880 62.290 636.020 110.430 ;
        RECT 634.960 62.150 636.020 62.290 ;
        RECT 634.960 17.330 635.100 62.150 ;
        RECT 419.160 17.010 419.420 17.330 ;
        RECT 634.900 17.010 635.160 17.330 ;
        RECT 419.220 2.400 419.360 17.010 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 634.430 917.520 634.710 917.800 ;
        RECT 635.350 917.520 635.630 917.800 ;
        RECT 634.890 385.760 635.170 386.040 ;
        RECT 635.810 385.760 636.090 386.040 ;
      LAYER met3 ;
        RECT 634.405 917.810 634.735 917.825 ;
        RECT 635.325 917.810 635.655 917.825 ;
        RECT 634.405 917.510 635.655 917.810 ;
        RECT 634.405 917.495 634.735 917.510 ;
        RECT 635.325 917.495 635.655 917.510 ;
        RECT 634.865 386.050 635.195 386.065 ;
        RECT 635.785 386.050 636.115 386.065 ;
        RECT 634.865 385.750 636.115 386.050 ;
        RECT 634.865 385.735 635.195 385.750 ;
        RECT 635.785 385.735 636.115 385.750 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 26.080 436.930 26.140 ;
        RECT 656.030 26.080 656.350 26.140 ;
        RECT 436.610 25.940 656.350 26.080 ;
        RECT 436.610 25.880 436.930 25.940 ;
        RECT 656.030 25.880 656.350 25.940 ;
      LAYER via ;
        RECT 436.640 25.880 436.900 26.140 ;
        RECT 656.060 25.880 656.320 26.140 ;
      LAYER met2 ;
        RECT 655.600 1600.450 655.880 1604.000 ;
        RECT 655.600 1600.310 656.260 1600.450 ;
        RECT 655.600 1600.000 655.880 1600.310 ;
        RECT 656.120 26.170 656.260 1600.310 ;
        RECT 436.640 25.850 436.900 26.170 ;
        RECT 656.060 25.850 656.320 26.170 ;
        RECT 436.700 2.400 436.840 25.850 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 455.010 25.740 455.330 25.800 ;
        RECT 669.830 25.740 670.150 25.800 ;
        RECT 455.010 25.600 670.150 25.740 ;
        RECT 455.010 25.540 455.330 25.600 ;
        RECT 669.830 25.540 670.150 25.600 ;
      LAYER via ;
        RECT 455.040 25.540 455.300 25.800 ;
        RECT 669.860 25.540 670.120 25.800 ;
      LAYER met2 ;
        RECT 670.320 1600.450 670.600 1604.000 ;
        RECT 669.920 1600.310 670.600 1600.450 ;
        RECT 669.920 25.830 670.060 1600.310 ;
        RECT 670.320 1600.000 670.600 1600.310 ;
        RECT 455.040 25.510 455.300 25.830 ;
        RECT 669.860 25.510 670.120 25.830 ;
        RECT 455.100 13.330 455.240 25.510 ;
        RECT 454.640 13.190 455.240 13.330 ;
        RECT 454.640 2.400 454.780 13.190 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 26.420 472.810 26.480 ;
        RECT 683.630 26.420 683.950 26.480 ;
        RECT 472.490 26.280 683.950 26.420 ;
        RECT 472.490 26.220 472.810 26.280 ;
        RECT 683.630 26.220 683.950 26.280 ;
      LAYER via ;
        RECT 472.520 26.220 472.780 26.480 ;
        RECT 683.660 26.220 683.920 26.480 ;
      LAYER met2 ;
        RECT 685.040 1600.450 685.320 1604.000 ;
        RECT 683.720 1600.310 685.320 1600.450 ;
        RECT 683.720 26.510 683.860 1600.310 ;
        RECT 685.040 1600.000 685.320 1600.310 ;
        RECT 472.520 26.190 472.780 26.510 ;
        RECT 683.660 26.190 683.920 26.510 ;
        RECT 472.580 2.400 472.720 26.190 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 679.490 1589.060 679.810 1589.120 ;
        RECT 699.270 1589.060 699.590 1589.120 ;
        RECT 679.490 1588.920 699.590 1589.060 ;
        RECT 679.490 1588.860 679.810 1588.920 ;
        RECT 699.270 1588.860 699.590 1588.920 ;
        RECT 490.430 19.280 490.750 19.340 ;
        RECT 676.270 19.280 676.590 19.340 ;
        RECT 490.430 19.140 676.590 19.280 ;
        RECT 490.430 19.080 490.750 19.140 ;
        RECT 676.270 19.080 676.590 19.140 ;
      LAYER via ;
        RECT 679.520 1588.860 679.780 1589.120 ;
        RECT 699.300 1588.860 699.560 1589.120 ;
        RECT 490.460 19.080 490.720 19.340 ;
        RECT 676.300 19.080 676.560 19.340 ;
      LAYER met2 ;
        RECT 699.300 1600.000 699.580 1604.000 ;
        RECT 699.360 1589.150 699.500 1600.000 ;
        RECT 679.520 1588.830 679.780 1589.150 ;
        RECT 699.300 1588.830 699.560 1589.150 ;
        RECT 679.580 19.565 679.720 1588.830 ;
        RECT 490.460 19.050 490.720 19.370 ;
        RECT 676.290 19.195 676.570 19.565 ;
        RECT 679.510 19.195 679.790 19.565 ;
        RECT 676.300 19.050 676.560 19.195 ;
        RECT 490.520 2.400 490.660 19.050 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 676.290 19.240 676.570 19.520 ;
        RECT 679.510 19.240 679.790 19.520 ;
      LAYER met3 ;
        RECT 676.265 19.530 676.595 19.545 ;
        RECT 679.485 19.530 679.815 19.545 ;
        RECT 676.265 19.230 679.815 19.530 ;
        RECT 676.265 19.215 676.595 19.230 ;
        RECT 679.485 19.215 679.815 19.230 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 676.345 18.445 677.435 18.615 ;
      LAYER mcon ;
        RECT 677.265 18.445 677.435 18.615 ;
      LAYER met1 ;
        RECT 700.190 1587.360 700.510 1587.420 ;
        RECT 712.150 1587.360 712.470 1587.420 ;
        RECT 700.190 1587.220 712.470 1587.360 ;
        RECT 700.190 1587.160 700.510 1587.220 ;
        RECT 712.150 1587.160 712.470 1587.220 ;
        RECT 507.910 18.600 508.230 18.660 ;
        RECT 676.285 18.600 676.575 18.645 ;
        RECT 507.910 18.460 676.575 18.600 ;
        RECT 507.910 18.400 508.230 18.460 ;
        RECT 676.285 18.415 676.575 18.460 ;
        RECT 677.205 18.600 677.495 18.645 ;
        RECT 700.190 18.600 700.510 18.660 ;
        RECT 677.205 18.460 700.510 18.600 ;
        RECT 677.205 18.415 677.495 18.460 ;
        RECT 700.190 18.400 700.510 18.460 ;
      LAYER via ;
        RECT 700.220 1587.160 700.480 1587.420 ;
        RECT 712.180 1587.160 712.440 1587.420 ;
        RECT 507.940 18.400 508.200 18.660 ;
        RECT 700.220 18.400 700.480 18.660 ;
      LAYER met2 ;
        RECT 714.020 1600.450 714.300 1604.000 ;
        RECT 712.240 1600.310 714.300 1600.450 ;
        RECT 712.240 1587.450 712.380 1600.310 ;
        RECT 714.020 1600.000 714.300 1600.310 ;
        RECT 700.220 1587.130 700.480 1587.450 ;
        RECT 712.180 1587.130 712.440 1587.450 ;
        RECT 700.280 18.690 700.420 1587.130 ;
        RECT 507.940 18.370 508.200 18.690 ;
        RECT 700.220 18.370 700.480 18.690 ;
        RECT 508.000 2.400 508.140 18.370 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 26.760 526.170 26.820 ;
        RECT 724.570 26.760 724.890 26.820 ;
        RECT 525.850 26.620 724.890 26.760 ;
        RECT 525.850 26.560 526.170 26.620 ;
        RECT 724.570 26.560 724.890 26.620 ;
      LAYER via ;
        RECT 525.880 26.560 526.140 26.820 ;
        RECT 724.600 26.560 724.860 26.820 ;
      LAYER met2 ;
        RECT 728.280 1600.450 728.560 1604.000 ;
        RECT 724.660 1600.310 728.560 1600.450 ;
        RECT 724.660 26.850 724.800 1600.310 ;
        RECT 728.280 1600.000 728.560 1600.310 ;
        RECT 525.880 26.530 526.140 26.850 ;
        RECT 724.600 26.530 724.860 26.850 ;
        RECT 525.940 2.400 526.080 26.530 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 676.805 19.465 676.975 23.375 ;
      LAYER mcon ;
        RECT 676.805 23.205 676.975 23.375 ;
      LAYER met1 ;
        RECT 713.990 1588.720 714.310 1588.780 ;
        RECT 742.970 1588.720 743.290 1588.780 ;
        RECT 713.990 1588.580 743.290 1588.720 ;
        RECT 713.990 1588.520 714.310 1588.580 ;
        RECT 742.970 1588.520 743.290 1588.580 ;
        RECT 676.745 23.360 677.035 23.405 ;
        RECT 713.990 23.360 714.310 23.420 ;
        RECT 676.745 23.220 714.310 23.360 ;
        RECT 676.745 23.175 677.035 23.220 ;
        RECT 713.990 23.160 714.310 23.220 ;
        RECT 543.790 19.620 544.110 19.680 ;
        RECT 676.745 19.620 677.035 19.665 ;
        RECT 543.790 19.480 677.035 19.620 ;
        RECT 543.790 19.420 544.110 19.480 ;
        RECT 676.745 19.435 677.035 19.480 ;
      LAYER via ;
        RECT 714.020 1588.520 714.280 1588.780 ;
        RECT 743.000 1588.520 743.260 1588.780 ;
        RECT 714.020 23.160 714.280 23.420 ;
        RECT 543.820 19.420 544.080 19.680 ;
      LAYER met2 ;
        RECT 743.000 1600.000 743.280 1604.000 ;
        RECT 743.060 1588.810 743.200 1600.000 ;
        RECT 714.020 1588.490 714.280 1588.810 ;
        RECT 743.000 1588.490 743.260 1588.810 ;
        RECT 714.080 23.450 714.220 1588.490 ;
        RECT 714.020 23.130 714.280 23.450 ;
        RECT 543.820 19.390 544.080 19.710 ;
        RECT 543.880 2.400 544.020 19.390 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 752.705 1207.425 752.875 1255.875 ;
        RECT 752.245 565.845 752.415 613.955 ;
        RECT 752.245 510.765 752.415 524.875 ;
        RECT 753.165 421.005 753.335 496.995 ;
        RECT 753.625 331.245 753.795 396.695 ;
        RECT 676.805 17.425 677.895 17.595 ;
      LAYER mcon ;
        RECT 752.705 1255.705 752.875 1255.875 ;
        RECT 752.245 613.785 752.415 613.955 ;
        RECT 752.245 524.705 752.415 524.875 ;
        RECT 753.165 496.825 753.335 496.995 ;
        RECT 753.625 396.525 753.795 396.695 ;
        RECT 677.725 17.425 677.895 17.595 ;
      LAYER met1 ;
        RECT 752.630 1497.260 752.950 1497.320 ;
        RECT 753.550 1497.260 753.870 1497.320 ;
        RECT 752.630 1497.120 753.870 1497.260 ;
        RECT 752.630 1497.060 752.950 1497.120 ;
        RECT 753.550 1497.060 753.870 1497.120 ;
        RECT 752.630 1400.700 752.950 1400.760 ;
        RECT 753.550 1400.700 753.870 1400.760 ;
        RECT 752.630 1400.560 753.870 1400.700 ;
        RECT 752.630 1400.500 752.950 1400.560 ;
        RECT 753.550 1400.500 753.870 1400.560 ;
        RECT 752.630 1317.400 752.950 1317.460 ;
        RECT 753.550 1317.400 753.870 1317.460 ;
        RECT 752.630 1317.260 753.870 1317.400 ;
        RECT 752.630 1317.200 752.950 1317.260 ;
        RECT 753.550 1317.200 753.870 1317.260 ;
        RECT 752.630 1304.140 752.950 1304.200 ;
        RECT 753.550 1304.140 753.870 1304.200 ;
        RECT 752.630 1304.000 753.870 1304.140 ;
        RECT 752.630 1303.940 752.950 1304.000 ;
        RECT 753.550 1303.940 753.870 1304.000 ;
        RECT 752.630 1255.860 752.950 1255.920 ;
        RECT 752.435 1255.720 752.950 1255.860 ;
        RECT 752.630 1255.660 752.950 1255.720 ;
        RECT 752.645 1207.580 752.935 1207.625 ;
        RECT 753.550 1207.580 753.870 1207.640 ;
        RECT 752.645 1207.440 753.870 1207.580 ;
        RECT 752.645 1207.395 752.935 1207.440 ;
        RECT 753.550 1207.380 753.870 1207.440 ;
        RECT 752.630 1159.300 752.950 1159.360 ;
        RECT 753.550 1159.300 753.870 1159.360 ;
        RECT 752.630 1159.160 753.870 1159.300 ;
        RECT 752.630 1159.100 752.950 1159.160 ;
        RECT 753.550 1159.100 753.870 1159.160 ;
        RECT 752.630 1062.740 752.950 1062.800 ;
        RECT 753.550 1062.740 753.870 1062.800 ;
        RECT 752.630 1062.600 753.870 1062.740 ;
        RECT 752.630 1062.540 752.950 1062.600 ;
        RECT 753.550 1062.540 753.870 1062.600 ;
        RECT 753.550 966.180 753.870 966.240 ;
        RECT 754.470 966.180 754.790 966.240 ;
        RECT 753.550 966.040 754.790 966.180 ;
        RECT 753.550 965.980 753.870 966.040 ;
        RECT 754.470 965.980 754.790 966.040 ;
        RECT 753.550 869.620 753.870 869.680 ;
        RECT 754.470 869.620 754.790 869.680 ;
        RECT 753.550 869.480 754.790 869.620 ;
        RECT 753.550 869.420 753.870 869.480 ;
        RECT 754.470 869.420 754.790 869.480 ;
        RECT 752.630 821.000 752.950 821.060 ;
        RECT 754.470 821.000 754.790 821.060 ;
        RECT 752.630 820.860 754.790 821.000 ;
        RECT 752.630 820.800 752.950 820.860 ;
        RECT 754.470 820.800 754.790 820.860 ;
        RECT 752.170 621.420 752.490 621.480 ;
        RECT 753.090 621.420 753.410 621.480 ;
        RECT 752.170 621.280 753.410 621.420 ;
        RECT 752.170 621.220 752.490 621.280 ;
        RECT 753.090 621.220 753.410 621.280 ;
        RECT 752.170 613.940 752.490 614.000 ;
        RECT 751.975 613.800 752.490 613.940 ;
        RECT 752.170 613.740 752.490 613.800 ;
        RECT 752.185 566.000 752.475 566.045 ;
        RECT 752.630 566.000 752.950 566.060 ;
        RECT 752.185 565.860 752.950 566.000 ;
        RECT 752.185 565.815 752.475 565.860 ;
        RECT 752.630 565.800 752.950 565.860 ;
        RECT 752.185 524.860 752.475 524.905 ;
        RECT 752.630 524.860 752.950 524.920 ;
        RECT 752.185 524.720 752.950 524.860 ;
        RECT 752.185 524.675 752.475 524.720 ;
        RECT 752.630 524.660 752.950 524.720 ;
        RECT 752.170 510.920 752.490 510.980 ;
        RECT 752.170 510.780 752.685 510.920 ;
        RECT 752.170 510.720 752.490 510.780 ;
        RECT 752.170 496.980 752.490 497.040 ;
        RECT 753.105 496.980 753.395 497.025 ;
        RECT 752.170 496.840 753.395 496.980 ;
        RECT 752.170 496.780 752.490 496.840 ;
        RECT 753.105 496.795 753.395 496.840 ;
        RECT 753.090 421.160 753.410 421.220 ;
        RECT 752.895 421.020 753.410 421.160 ;
        RECT 753.090 420.960 753.410 421.020 ;
        RECT 753.090 396.680 753.410 396.740 ;
        RECT 753.565 396.680 753.855 396.725 ;
        RECT 753.090 396.540 753.855 396.680 ;
        RECT 753.090 396.480 753.410 396.540 ;
        RECT 753.565 396.495 753.855 396.540 ;
        RECT 753.550 331.400 753.870 331.460 ;
        RECT 753.355 331.260 753.870 331.400 ;
        RECT 753.550 331.200 753.870 331.260 ;
        RECT 753.090 255.720 753.410 255.980 ;
        RECT 753.180 255.300 753.320 255.720 ;
        RECT 753.090 255.040 753.410 255.300 ;
        RECT 752.630 241.300 752.950 241.360 ;
        RECT 753.550 241.300 753.870 241.360 ;
        RECT 752.630 241.160 753.870 241.300 ;
        RECT 752.630 241.100 752.950 241.160 ;
        RECT 753.550 241.100 753.870 241.160 ;
        RECT 753.090 159.160 753.410 159.420 ;
        RECT 753.180 158.740 753.320 159.160 ;
        RECT 753.090 158.480 753.410 158.740 ;
        RECT 752.630 144.740 752.950 144.800 ;
        RECT 753.550 144.740 753.870 144.800 ;
        RECT 752.630 144.600 753.870 144.740 ;
        RECT 752.630 144.540 752.950 144.600 ;
        RECT 753.550 144.540 753.870 144.600 ;
        RECT 561.730 17.580 562.050 17.640 ;
        RECT 676.745 17.580 677.035 17.625 ;
        RECT 561.730 17.440 677.035 17.580 ;
        RECT 561.730 17.380 562.050 17.440 ;
        RECT 676.745 17.395 677.035 17.440 ;
        RECT 677.665 17.580 677.955 17.625 ;
        RECT 753.550 17.580 753.870 17.640 ;
        RECT 677.665 17.440 753.870 17.580 ;
        RECT 677.665 17.395 677.955 17.440 ;
        RECT 753.550 17.380 753.870 17.440 ;
      LAYER via ;
        RECT 752.660 1497.060 752.920 1497.320 ;
        RECT 753.580 1497.060 753.840 1497.320 ;
        RECT 752.660 1400.500 752.920 1400.760 ;
        RECT 753.580 1400.500 753.840 1400.760 ;
        RECT 752.660 1317.200 752.920 1317.460 ;
        RECT 753.580 1317.200 753.840 1317.460 ;
        RECT 752.660 1303.940 752.920 1304.200 ;
        RECT 753.580 1303.940 753.840 1304.200 ;
        RECT 752.660 1255.660 752.920 1255.920 ;
        RECT 753.580 1207.380 753.840 1207.640 ;
        RECT 752.660 1159.100 752.920 1159.360 ;
        RECT 753.580 1159.100 753.840 1159.360 ;
        RECT 752.660 1062.540 752.920 1062.800 ;
        RECT 753.580 1062.540 753.840 1062.800 ;
        RECT 753.580 965.980 753.840 966.240 ;
        RECT 754.500 965.980 754.760 966.240 ;
        RECT 753.580 869.420 753.840 869.680 ;
        RECT 754.500 869.420 754.760 869.680 ;
        RECT 752.660 820.800 752.920 821.060 ;
        RECT 754.500 820.800 754.760 821.060 ;
        RECT 752.200 621.220 752.460 621.480 ;
        RECT 753.120 621.220 753.380 621.480 ;
        RECT 752.200 613.740 752.460 614.000 ;
        RECT 752.660 565.800 752.920 566.060 ;
        RECT 752.660 524.660 752.920 524.920 ;
        RECT 752.200 510.720 752.460 510.980 ;
        RECT 752.200 496.780 752.460 497.040 ;
        RECT 753.120 420.960 753.380 421.220 ;
        RECT 753.120 396.480 753.380 396.740 ;
        RECT 753.580 331.200 753.840 331.460 ;
        RECT 753.120 255.720 753.380 255.980 ;
        RECT 753.120 255.040 753.380 255.300 ;
        RECT 752.660 241.100 752.920 241.360 ;
        RECT 753.580 241.100 753.840 241.360 ;
        RECT 753.120 159.160 753.380 159.420 ;
        RECT 753.120 158.480 753.380 158.740 ;
        RECT 752.660 144.540 752.920 144.800 ;
        RECT 753.580 144.540 753.840 144.800 ;
        RECT 561.760 17.380 562.020 17.640 ;
        RECT 753.580 17.380 753.840 17.640 ;
      LAYER met2 ;
        RECT 757.720 1600.450 758.000 1604.000 ;
        RECT 753.180 1600.310 758.000 1600.450 ;
        RECT 753.180 1580.050 753.320 1600.310 ;
        RECT 757.720 1600.000 758.000 1600.310 ;
        RECT 752.720 1579.910 753.320 1580.050 ;
        RECT 752.720 1510.690 752.860 1579.910 ;
        RECT 752.720 1510.550 753.780 1510.690 ;
        RECT 753.640 1497.350 753.780 1510.550 ;
        RECT 752.660 1497.030 752.920 1497.350 ;
        RECT 753.580 1497.030 753.840 1497.350 ;
        RECT 752.720 1414.130 752.860 1497.030 ;
        RECT 752.720 1413.990 753.780 1414.130 ;
        RECT 753.640 1400.790 753.780 1413.990 ;
        RECT 752.660 1400.470 752.920 1400.790 ;
        RECT 753.580 1400.470 753.840 1400.790 ;
        RECT 752.720 1317.490 752.860 1400.470 ;
        RECT 752.660 1317.170 752.920 1317.490 ;
        RECT 753.580 1317.170 753.840 1317.490 ;
        RECT 753.640 1304.230 753.780 1317.170 ;
        RECT 752.660 1303.910 752.920 1304.230 ;
        RECT 753.580 1303.910 753.840 1304.230 ;
        RECT 752.720 1255.950 752.860 1303.910 ;
        RECT 752.660 1255.630 752.920 1255.950 ;
        RECT 753.580 1207.350 753.840 1207.670 ;
        RECT 753.640 1159.390 753.780 1207.350 ;
        RECT 752.660 1159.070 752.920 1159.390 ;
        RECT 753.580 1159.070 753.840 1159.390 ;
        RECT 752.720 1124.450 752.860 1159.070 ;
        RECT 752.720 1124.310 753.780 1124.450 ;
        RECT 753.640 1062.830 753.780 1124.310 ;
        RECT 752.660 1062.510 752.920 1062.830 ;
        RECT 753.580 1062.510 753.840 1062.830 ;
        RECT 752.720 1014.405 752.860 1062.510 ;
        RECT 752.650 1014.035 752.930 1014.405 ;
        RECT 754.490 1014.035 754.770 1014.405 ;
        RECT 754.560 966.270 754.700 1014.035 ;
        RECT 753.580 965.950 753.840 966.270 ;
        RECT 754.500 965.950 754.760 966.270 ;
        RECT 753.640 931.330 753.780 965.950 ;
        RECT 752.720 931.190 753.780 931.330 ;
        RECT 752.720 917.845 752.860 931.190 ;
        RECT 752.650 917.475 752.930 917.845 ;
        RECT 754.490 917.475 754.770 917.845 ;
        RECT 754.560 869.710 754.700 917.475 ;
        RECT 753.580 869.390 753.840 869.710 ;
        RECT 754.500 869.390 754.760 869.710 ;
        RECT 753.640 834.770 753.780 869.390 ;
        RECT 752.720 834.630 753.780 834.770 ;
        RECT 752.720 821.090 752.860 834.630 ;
        RECT 752.660 820.770 752.920 821.090 ;
        RECT 754.500 820.770 754.760 821.090 ;
        RECT 754.560 773.005 754.700 820.770 ;
        RECT 753.570 772.635 753.850 773.005 ;
        RECT 754.490 772.635 754.770 773.005 ;
        RECT 753.640 738.210 753.780 772.635 ;
        RECT 753.180 738.070 753.780 738.210 ;
        RECT 753.180 690.725 753.320 738.070 ;
        RECT 753.110 690.355 753.390 690.725 ;
        RECT 752.650 669.275 752.930 669.645 ;
        RECT 752.720 645.730 752.860 669.275 ;
        RECT 752.720 645.590 753.320 645.730 ;
        RECT 753.180 621.510 753.320 645.590 ;
        RECT 752.200 621.190 752.460 621.510 ;
        RECT 753.120 621.190 753.380 621.510 ;
        RECT 752.260 614.030 752.400 621.190 ;
        RECT 752.200 613.710 752.460 614.030 ;
        RECT 752.660 565.770 752.920 566.090 ;
        RECT 752.720 524.950 752.860 565.770 ;
        RECT 752.660 524.630 752.920 524.950 ;
        RECT 752.200 510.690 752.460 511.010 ;
        RECT 752.260 510.525 752.400 510.690 ;
        RECT 752.190 510.155 752.470 510.525 ;
        RECT 752.190 509.475 752.470 509.845 ;
        RECT 752.260 497.070 752.400 509.475 ;
        RECT 752.200 496.750 752.460 497.070 ;
        RECT 753.120 420.930 753.380 421.250 ;
        RECT 753.180 396.770 753.320 420.930 ;
        RECT 753.120 396.450 753.380 396.770 ;
        RECT 753.580 331.170 753.840 331.490 ;
        RECT 753.640 303.690 753.780 331.170 ;
        RECT 752.720 303.550 753.780 303.690 ;
        RECT 752.720 266.290 752.860 303.550 ;
        RECT 752.720 266.150 753.320 266.290 ;
        RECT 753.180 256.010 753.320 266.150 ;
        RECT 753.120 255.690 753.380 256.010 ;
        RECT 753.120 255.010 753.380 255.330 ;
        RECT 753.180 241.810 753.320 255.010 ;
        RECT 753.180 241.670 753.780 241.810 ;
        RECT 753.640 241.390 753.780 241.670 ;
        RECT 752.660 241.070 752.920 241.390 ;
        RECT 753.580 241.070 753.840 241.390 ;
        RECT 752.720 175.850 752.860 241.070 ;
        RECT 752.720 175.710 753.320 175.850 ;
        RECT 753.180 159.450 753.320 175.710 ;
        RECT 753.120 159.130 753.380 159.450 ;
        RECT 753.120 158.450 753.380 158.770 ;
        RECT 753.180 145.250 753.320 158.450 ;
        RECT 753.180 145.110 753.780 145.250 ;
        RECT 753.640 144.830 753.780 145.110 ;
        RECT 752.660 144.510 752.920 144.830 ;
        RECT 753.580 144.510 753.840 144.830 ;
        RECT 752.720 62.290 752.860 144.510 ;
        RECT 752.720 62.150 753.780 62.290 ;
        RECT 753.640 17.670 753.780 62.150 ;
        RECT 561.760 17.350 562.020 17.670 ;
        RECT 753.580 17.350 753.840 17.670 ;
        RECT 561.820 2.400 561.960 17.350 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 752.650 1014.080 752.930 1014.360 ;
        RECT 754.490 1014.080 754.770 1014.360 ;
        RECT 752.650 917.520 752.930 917.800 ;
        RECT 754.490 917.520 754.770 917.800 ;
        RECT 753.570 772.680 753.850 772.960 ;
        RECT 754.490 772.680 754.770 772.960 ;
        RECT 753.110 690.400 753.390 690.680 ;
        RECT 752.650 669.320 752.930 669.600 ;
        RECT 752.190 510.200 752.470 510.480 ;
        RECT 752.190 509.520 752.470 509.800 ;
      LAYER met3 ;
        RECT 752.625 1014.370 752.955 1014.385 ;
        RECT 754.465 1014.370 754.795 1014.385 ;
        RECT 752.625 1014.070 754.795 1014.370 ;
        RECT 752.625 1014.055 752.955 1014.070 ;
        RECT 754.465 1014.055 754.795 1014.070 ;
        RECT 752.625 917.810 752.955 917.825 ;
        RECT 754.465 917.810 754.795 917.825 ;
        RECT 752.625 917.510 754.795 917.810 ;
        RECT 752.625 917.495 752.955 917.510 ;
        RECT 754.465 917.495 754.795 917.510 ;
        RECT 753.545 772.970 753.875 772.985 ;
        RECT 754.465 772.970 754.795 772.985 ;
        RECT 753.545 772.670 754.795 772.970 ;
        RECT 753.545 772.655 753.875 772.670 ;
        RECT 754.465 772.655 754.795 772.670 ;
        RECT 753.085 690.700 753.415 690.705 ;
        RECT 752.830 690.690 753.415 690.700 ;
        RECT 752.630 690.390 753.415 690.690 ;
        RECT 752.830 690.380 753.415 690.390 ;
        RECT 753.085 690.375 753.415 690.380 ;
        RECT 752.625 669.620 752.955 669.625 ;
        RECT 752.625 669.610 753.210 669.620 ;
        RECT 752.625 669.310 753.410 669.610 ;
        RECT 752.625 669.300 753.210 669.310 ;
        RECT 752.625 669.295 752.955 669.300 ;
        RECT 752.165 510.490 752.495 510.505 ;
        RECT 751.950 510.175 752.495 510.490 ;
        RECT 751.950 509.825 752.250 510.175 ;
        RECT 751.950 509.510 752.495 509.825 ;
        RECT 752.165 509.495 752.495 509.510 ;
      LAYER via3 ;
        RECT 752.860 690.380 753.180 690.700 ;
        RECT 752.860 669.300 753.180 669.620 ;
      LAYER met4 ;
        RECT 752.855 690.375 753.185 690.705 ;
        RECT 752.870 669.625 753.170 690.375 ;
        RECT 752.855 669.295 753.185 669.625 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 766.505 1207.425 766.675 1255.875 ;
        RECT 766.505 662.405 766.675 710.515 ;
        RECT 766.045 565.845 766.215 613.955 ;
        RECT 766.045 427.805 766.215 475.915 ;
        RECT 766.045 379.525 766.215 422.875 ;
        RECT 676.805 18.105 677.895 18.275 ;
      LAYER mcon ;
        RECT 766.505 1255.705 766.675 1255.875 ;
        RECT 766.505 710.345 766.675 710.515 ;
        RECT 766.045 613.785 766.215 613.955 ;
        RECT 766.045 475.745 766.215 475.915 ;
        RECT 766.045 422.705 766.215 422.875 ;
        RECT 677.725 18.105 677.895 18.275 ;
      LAYER met1 ;
        RECT 766.430 1497.260 766.750 1497.320 ;
        RECT 767.350 1497.260 767.670 1497.320 ;
        RECT 766.430 1497.120 767.670 1497.260 ;
        RECT 766.430 1497.060 766.750 1497.120 ;
        RECT 767.350 1497.060 767.670 1497.120 ;
        RECT 766.430 1413.960 766.750 1414.020 ;
        RECT 767.350 1413.960 767.670 1414.020 ;
        RECT 766.430 1413.820 767.670 1413.960 ;
        RECT 766.430 1413.760 766.750 1413.820 ;
        RECT 767.350 1413.760 767.670 1413.820 ;
        RECT 766.430 1400.700 766.750 1400.760 ;
        RECT 767.350 1400.700 767.670 1400.760 ;
        RECT 766.430 1400.560 767.670 1400.700 ;
        RECT 766.430 1400.500 766.750 1400.560 ;
        RECT 767.350 1400.500 767.670 1400.560 ;
        RECT 766.430 1304.140 766.750 1304.200 ;
        RECT 767.350 1304.140 767.670 1304.200 ;
        RECT 766.430 1304.000 767.670 1304.140 ;
        RECT 766.430 1303.940 766.750 1304.000 ;
        RECT 767.350 1303.940 767.670 1304.000 ;
        RECT 766.430 1255.860 766.750 1255.920 ;
        RECT 766.235 1255.720 766.750 1255.860 ;
        RECT 766.430 1255.660 766.750 1255.720 ;
        RECT 766.445 1207.580 766.735 1207.625 ;
        RECT 767.350 1207.580 767.670 1207.640 ;
        RECT 766.445 1207.440 767.670 1207.580 ;
        RECT 766.445 1207.395 766.735 1207.440 ;
        RECT 767.350 1207.380 767.670 1207.440 ;
        RECT 766.430 1159.300 766.750 1159.360 ;
        RECT 767.810 1159.300 768.130 1159.360 ;
        RECT 766.430 1159.160 768.130 1159.300 ;
        RECT 766.430 1159.100 766.750 1159.160 ;
        RECT 767.810 1159.100 768.130 1159.160 ;
        RECT 767.350 1111.020 767.670 1111.080 ;
        RECT 767.810 1111.020 768.130 1111.080 ;
        RECT 767.350 1110.880 768.130 1111.020 ;
        RECT 767.350 1110.820 767.670 1110.880 ;
        RECT 767.810 1110.820 768.130 1110.880 ;
        RECT 766.430 1086.880 766.750 1086.940 ;
        RECT 767.810 1086.880 768.130 1086.940 ;
        RECT 766.430 1086.740 768.130 1086.880 ;
        RECT 766.430 1086.680 766.750 1086.740 ;
        RECT 767.810 1086.680 768.130 1086.740 ;
        RECT 767.350 966.180 767.670 966.240 ;
        RECT 768.270 966.180 768.590 966.240 ;
        RECT 767.350 966.040 768.590 966.180 ;
        RECT 767.350 965.980 767.670 966.040 ;
        RECT 768.270 965.980 768.590 966.040 ;
        RECT 767.350 869.620 767.670 869.680 ;
        RECT 768.270 869.620 768.590 869.680 ;
        RECT 767.350 869.480 768.590 869.620 ;
        RECT 767.350 869.420 767.670 869.480 ;
        RECT 768.270 869.420 768.590 869.480 ;
        RECT 766.430 821.000 766.750 821.060 ;
        RECT 768.270 821.000 768.590 821.060 ;
        RECT 766.430 820.860 768.590 821.000 ;
        RECT 766.430 820.800 766.750 820.860 ;
        RECT 768.270 820.800 768.590 820.860 ;
        RECT 766.890 738.040 767.210 738.100 ;
        RECT 767.350 738.040 767.670 738.100 ;
        RECT 766.890 737.900 767.670 738.040 ;
        RECT 766.890 737.840 767.210 737.900 ;
        RECT 767.350 737.840 767.670 737.900 ;
        RECT 766.445 710.500 766.735 710.545 ;
        RECT 766.890 710.500 767.210 710.560 ;
        RECT 766.445 710.360 767.210 710.500 ;
        RECT 766.445 710.315 766.735 710.360 ;
        RECT 766.890 710.300 767.210 710.360 ;
        RECT 766.430 662.560 766.750 662.620 ;
        RECT 766.235 662.420 766.750 662.560 ;
        RECT 766.430 662.360 766.750 662.420 ;
        RECT 766.430 642.160 766.750 642.220 ;
        RECT 766.060 642.020 766.750 642.160 ;
        RECT 766.060 641.540 766.200 642.020 ;
        RECT 766.430 641.960 766.750 642.020 ;
        RECT 765.970 641.280 766.290 641.540 ;
        RECT 765.970 613.940 766.290 614.000 ;
        RECT 765.775 613.800 766.290 613.940 ;
        RECT 765.970 613.740 766.290 613.800 ;
        RECT 765.985 566.000 766.275 566.045 ;
        RECT 766.430 566.000 766.750 566.060 ;
        RECT 765.985 565.860 766.750 566.000 ;
        RECT 765.985 565.815 766.275 565.860 ;
        RECT 766.430 565.800 766.750 565.860 ;
        RECT 766.430 545.600 766.750 545.660 ;
        RECT 766.060 545.460 766.750 545.600 ;
        RECT 766.060 544.980 766.200 545.460 ;
        RECT 766.430 545.400 766.750 545.460 ;
        RECT 765.970 544.720 766.290 544.980 ;
        RECT 765.985 475.900 766.275 475.945 ;
        RECT 766.430 475.900 766.750 475.960 ;
        RECT 765.985 475.760 766.750 475.900 ;
        RECT 765.985 475.715 766.275 475.760 ;
        RECT 766.430 475.700 766.750 475.760 ;
        RECT 765.970 427.960 766.290 428.020 ;
        RECT 765.970 427.820 766.485 427.960 ;
        RECT 765.970 427.760 766.290 427.820 ;
        RECT 765.970 422.860 766.290 422.920 ;
        RECT 765.970 422.720 766.485 422.860 ;
        RECT 765.970 422.660 766.290 422.720 ;
        RECT 765.985 379.680 766.275 379.725 ;
        RECT 767.350 379.680 767.670 379.740 ;
        RECT 765.985 379.540 767.670 379.680 ;
        RECT 765.985 379.495 766.275 379.540 ;
        RECT 767.350 379.480 767.670 379.540 ;
        RECT 766.430 241.300 766.750 241.360 ;
        RECT 767.350 241.300 767.670 241.360 ;
        RECT 766.430 241.160 767.670 241.300 ;
        RECT 766.430 241.100 766.750 241.160 ;
        RECT 767.350 241.100 767.670 241.160 ;
        RECT 766.890 159.020 767.210 159.080 ;
        RECT 766.890 158.880 767.580 159.020 ;
        RECT 766.890 158.820 767.210 158.880 ;
        RECT 767.440 158.400 767.580 158.880 ;
        RECT 767.350 158.140 767.670 158.400 ;
        RECT 766.430 144.740 766.750 144.800 ;
        RECT 767.350 144.740 767.670 144.800 ;
        RECT 766.430 144.600 767.670 144.740 ;
        RECT 766.430 144.540 766.750 144.600 ;
        RECT 767.350 144.540 767.670 144.600 ;
        RECT 579.670 18.260 579.990 18.320 ;
        RECT 676.745 18.260 677.035 18.305 ;
        RECT 579.670 18.120 677.035 18.260 ;
        RECT 579.670 18.060 579.990 18.120 ;
        RECT 676.745 18.075 677.035 18.120 ;
        RECT 677.665 18.260 677.955 18.305 ;
        RECT 767.350 18.260 767.670 18.320 ;
        RECT 677.665 18.120 767.670 18.260 ;
        RECT 677.665 18.075 677.955 18.120 ;
        RECT 767.350 18.060 767.670 18.120 ;
      LAYER via ;
        RECT 766.460 1497.060 766.720 1497.320 ;
        RECT 767.380 1497.060 767.640 1497.320 ;
        RECT 766.460 1413.760 766.720 1414.020 ;
        RECT 767.380 1413.760 767.640 1414.020 ;
        RECT 766.460 1400.500 766.720 1400.760 ;
        RECT 767.380 1400.500 767.640 1400.760 ;
        RECT 766.460 1303.940 766.720 1304.200 ;
        RECT 767.380 1303.940 767.640 1304.200 ;
        RECT 766.460 1255.660 766.720 1255.920 ;
        RECT 767.380 1207.380 767.640 1207.640 ;
        RECT 766.460 1159.100 766.720 1159.360 ;
        RECT 767.840 1159.100 768.100 1159.360 ;
        RECT 767.380 1110.820 767.640 1111.080 ;
        RECT 767.840 1110.820 768.100 1111.080 ;
        RECT 766.460 1086.680 766.720 1086.940 ;
        RECT 767.840 1086.680 768.100 1086.940 ;
        RECT 767.380 965.980 767.640 966.240 ;
        RECT 768.300 965.980 768.560 966.240 ;
        RECT 767.380 869.420 767.640 869.680 ;
        RECT 768.300 869.420 768.560 869.680 ;
        RECT 766.460 820.800 766.720 821.060 ;
        RECT 768.300 820.800 768.560 821.060 ;
        RECT 766.920 737.840 767.180 738.100 ;
        RECT 767.380 737.840 767.640 738.100 ;
        RECT 766.920 710.300 767.180 710.560 ;
        RECT 766.460 662.360 766.720 662.620 ;
        RECT 766.460 641.960 766.720 642.220 ;
        RECT 766.000 641.280 766.260 641.540 ;
        RECT 766.000 613.740 766.260 614.000 ;
        RECT 766.460 565.800 766.720 566.060 ;
        RECT 766.460 545.400 766.720 545.660 ;
        RECT 766.000 544.720 766.260 544.980 ;
        RECT 766.460 475.700 766.720 475.960 ;
        RECT 766.000 427.760 766.260 428.020 ;
        RECT 766.000 422.660 766.260 422.920 ;
        RECT 767.380 379.480 767.640 379.740 ;
        RECT 766.460 241.100 766.720 241.360 ;
        RECT 767.380 241.100 767.640 241.360 ;
        RECT 766.920 158.820 767.180 159.080 ;
        RECT 767.380 158.140 767.640 158.400 ;
        RECT 766.460 144.540 766.720 144.800 ;
        RECT 767.380 144.540 767.640 144.800 ;
        RECT 579.700 18.060 579.960 18.320 ;
        RECT 767.380 18.060 767.640 18.320 ;
      LAYER met2 ;
        RECT 771.980 1601.130 772.260 1604.000 ;
        RECT 767.900 1600.990 772.260 1601.130 ;
        RECT 767.900 1580.050 768.040 1600.990 ;
        RECT 771.980 1600.000 772.260 1600.990 ;
        RECT 766.520 1579.910 768.040 1580.050 ;
        RECT 766.520 1510.690 766.660 1579.910 ;
        RECT 766.520 1510.550 767.580 1510.690 ;
        RECT 767.440 1497.350 767.580 1510.550 ;
        RECT 766.460 1497.030 766.720 1497.350 ;
        RECT 767.380 1497.030 767.640 1497.350 ;
        RECT 766.520 1414.050 766.660 1497.030 ;
        RECT 766.460 1413.730 766.720 1414.050 ;
        RECT 767.380 1413.730 767.640 1414.050 ;
        RECT 767.440 1400.790 767.580 1413.730 ;
        RECT 766.460 1400.470 766.720 1400.790 ;
        RECT 767.380 1400.470 767.640 1400.790 ;
        RECT 766.520 1317.570 766.660 1400.470 ;
        RECT 766.520 1317.430 767.580 1317.570 ;
        RECT 767.440 1304.230 767.580 1317.430 ;
        RECT 766.460 1303.910 766.720 1304.230 ;
        RECT 767.380 1303.910 767.640 1304.230 ;
        RECT 766.520 1255.950 766.660 1303.910 ;
        RECT 766.460 1255.630 766.720 1255.950 ;
        RECT 767.440 1207.670 767.580 1207.825 ;
        RECT 767.380 1207.410 767.640 1207.670 ;
        RECT 767.380 1207.350 768.040 1207.410 ;
        RECT 767.440 1207.270 768.040 1207.350 ;
        RECT 767.900 1159.390 768.040 1207.270 ;
        RECT 766.460 1159.245 766.720 1159.390 ;
        RECT 767.840 1159.245 768.100 1159.390 ;
        RECT 766.450 1158.875 766.730 1159.245 ;
        RECT 767.830 1158.875 768.110 1159.245 ;
        RECT 767.440 1111.110 767.580 1111.265 ;
        RECT 767.900 1111.110 768.040 1158.875 ;
        RECT 767.380 1110.850 767.640 1111.110 ;
        RECT 767.840 1110.850 768.100 1111.110 ;
        RECT 767.380 1110.790 768.100 1110.850 ;
        RECT 767.440 1110.710 768.040 1110.790 ;
        RECT 767.900 1086.970 768.040 1110.710 ;
        RECT 766.460 1086.650 766.720 1086.970 ;
        RECT 767.840 1086.650 768.100 1086.970 ;
        RECT 766.520 1028.570 766.660 1086.650 ;
        RECT 766.520 1028.430 767.120 1028.570 ;
        RECT 766.980 1027.890 767.120 1028.430 ;
        RECT 766.520 1027.750 767.120 1027.890 ;
        RECT 766.520 1014.405 766.660 1027.750 ;
        RECT 766.450 1014.035 766.730 1014.405 ;
        RECT 768.290 1014.035 768.570 1014.405 ;
        RECT 768.360 966.270 768.500 1014.035 ;
        RECT 767.380 965.950 767.640 966.270 ;
        RECT 768.300 965.950 768.560 966.270 ;
        RECT 767.440 931.330 767.580 965.950 ;
        RECT 766.520 931.190 767.580 931.330 ;
        RECT 766.520 917.845 766.660 931.190 ;
        RECT 766.450 917.475 766.730 917.845 ;
        RECT 768.290 917.475 768.570 917.845 ;
        RECT 768.360 869.710 768.500 917.475 ;
        RECT 767.380 869.390 767.640 869.710 ;
        RECT 768.300 869.390 768.560 869.710 ;
        RECT 767.440 834.770 767.580 869.390 ;
        RECT 766.520 834.630 767.580 834.770 ;
        RECT 766.520 821.090 766.660 834.630 ;
        RECT 766.460 820.770 766.720 821.090 ;
        RECT 768.300 820.770 768.560 821.090 ;
        RECT 768.360 773.005 768.500 820.770 ;
        RECT 767.370 772.635 767.650 773.005 ;
        RECT 768.290 772.635 768.570 773.005 ;
        RECT 767.440 738.130 767.580 772.635 ;
        RECT 766.920 737.810 767.180 738.130 ;
        RECT 767.380 737.810 767.640 738.130 ;
        RECT 766.980 710.590 767.120 737.810 ;
        RECT 766.920 710.270 767.180 710.590 ;
        RECT 766.460 662.330 766.720 662.650 ;
        RECT 766.520 642.250 766.660 662.330 ;
        RECT 766.460 641.930 766.720 642.250 ;
        RECT 766.000 641.250 766.260 641.570 ;
        RECT 766.060 614.030 766.200 641.250 ;
        RECT 766.000 613.710 766.260 614.030 ;
        RECT 766.460 565.770 766.720 566.090 ;
        RECT 766.520 545.690 766.660 565.770 ;
        RECT 766.460 545.370 766.720 545.690 ;
        RECT 766.000 544.690 766.260 545.010 ;
        RECT 766.060 524.125 766.200 544.690 ;
        RECT 765.990 523.755 766.270 524.125 ;
        RECT 766.450 495.875 766.730 496.245 ;
        RECT 766.520 475.990 766.660 495.875 ;
        RECT 766.460 475.670 766.720 475.990 ;
        RECT 766.000 427.730 766.260 428.050 ;
        RECT 766.060 422.950 766.200 427.730 ;
        RECT 766.000 422.630 766.260 422.950 ;
        RECT 767.380 379.450 767.640 379.770 ;
        RECT 767.440 303.690 767.580 379.450 ;
        RECT 766.520 303.550 767.580 303.690 ;
        RECT 766.520 266.290 766.660 303.550 ;
        RECT 766.520 266.150 767.120 266.290 ;
        RECT 766.980 264.930 767.120 266.150 ;
        RECT 766.520 264.790 767.120 264.930 ;
        RECT 766.520 254.730 766.660 264.790 ;
        RECT 766.520 254.590 767.580 254.730 ;
        RECT 767.440 241.390 767.580 254.590 ;
        RECT 766.460 241.070 766.720 241.390 ;
        RECT 767.380 241.070 767.640 241.390 ;
        RECT 766.520 175.850 766.660 241.070 ;
        RECT 766.520 175.710 767.120 175.850 ;
        RECT 766.980 159.110 767.120 175.710 ;
        RECT 766.920 158.790 767.180 159.110 ;
        RECT 767.380 158.110 767.640 158.430 ;
        RECT 767.440 144.830 767.580 158.110 ;
        RECT 766.460 144.510 766.720 144.830 ;
        RECT 767.380 144.510 767.640 144.830 ;
        RECT 766.520 62.290 766.660 144.510 ;
        RECT 766.520 62.150 767.580 62.290 ;
        RECT 767.440 18.350 767.580 62.150 ;
        RECT 579.700 18.030 579.960 18.350 ;
        RECT 767.380 18.030 767.640 18.350 ;
        RECT 579.760 2.400 579.900 18.030 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 766.450 1158.920 766.730 1159.200 ;
        RECT 767.830 1158.920 768.110 1159.200 ;
        RECT 766.450 1014.080 766.730 1014.360 ;
        RECT 768.290 1014.080 768.570 1014.360 ;
        RECT 766.450 917.520 766.730 917.800 ;
        RECT 768.290 917.520 768.570 917.800 ;
        RECT 767.370 772.680 767.650 772.960 ;
        RECT 768.290 772.680 768.570 772.960 ;
        RECT 765.990 523.800 766.270 524.080 ;
        RECT 766.450 495.920 766.730 496.200 ;
      LAYER met3 ;
        RECT 766.425 1159.210 766.755 1159.225 ;
        RECT 767.805 1159.210 768.135 1159.225 ;
        RECT 766.425 1158.910 768.135 1159.210 ;
        RECT 766.425 1158.895 766.755 1158.910 ;
        RECT 767.805 1158.895 768.135 1158.910 ;
        RECT 766.425 1014.370 766.755 1014.385 ;
        RECT 768.265 1014.370 768.595 1014.385 ;
        RECT 766.425 1014.070 768.595 1014.370 ;
        RECT 766.425 1014.055 766.755 1014.070 ;
        RECT 768.265 1014.055 768.595 1014.070 ;
        RECT 766.425 917.810 766.755 917.825 ;
        RECT 768.265 917.810 768.595 917.825 ;
        RECT 766.425 917.510 768.595 917.810 ;
        RECT 766.425 917.495 766.755 917.510 ;
        RECT 768.265 917.495 768.595 917.510 ;
        RECT 767.345 772.970 767.675 772.985 ;
        RECT 768.265 772.970 768.595 772.985 ;
        RECT 767.345 772.670 768.595 772.970 ;
        RECT 767.345 772.655 767.675 772.670 ;
        RECT 768.265 772.655 768.595 772.670 ;
        RECT 765.965 524.100 766.295 524.105 ;
        RECT 765.710 524.090 766.295 524.100 ;
        RECT 765.710 523.790 766.520 524.090 ;
        RECT 765.710 523.780 766.295 523.790 ;
        RECT 765.965 523.775 766.295 523.780 ;
        RECT 765.710 496.210 766.090 496.220 ;
        RECT 766.425 496.210 766.755 496.225 ;
        RECT 765.710 495.910 766.755 496.210 ;
        RECT 765.710 495.900 766.090 495.910 ;
        RECT 766.425 495.895 766.755 495.910 ;
      LAYER via3 ;
        RECT 765.740 523.780 766.060 524.100 ;
        RECT 765.740 495.900 766.060 496.220 ;
      LAYER met4 ;
        RECT 765.735 523.775 766.065 524.105 ;
        RECT 765.750 496.225 766.050 523.775 ;
        RECT 765.735 495.895 766.065 496.225 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 25.740 86.410 25.800 ;
        RECT 365.770 25.740 366.090 25.800 ;
        RECT 86.090 25.600 366.090 25.740 ;
        RECT 86.090 25.540 86.410 25.600 ;
        RECT 365.770 25.540 366.090 25.600 ;
      LAYER via ;
        RECT 86.120 25.540 86.380 25.800 ;
        RECT 365.800 25.540 366.060 25.800 ;
      LAYER met2 ;
        RECT 369.940 1600.450 370.220 1604.000 ;
        RECT 365.860 1600.310 370.220 1600.450 ;
        RECT 365.860 25.830 366.000 1600.310 ;
        RECT 369.940 1600.000 370.220 1600.310 ;
        RECT 86.120 25.510 86.380 25.830 ;
        RECT 365.800 25.510 366.060 25.830 ;
        RECT 86.180 2.400 86.320 25.510 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 24.040 597.470 24.100 ;
        RECT 787.130 24.040 787.450 24.100 ;
        RECT 597.150 23.900 787.450 24.040 ;
        RECT 597.150 23.840 597.470 23.900 ;
        RECT 787.130 23.840 787.450 23.900 ;
      LAYER via ;
        RECT 597.180 23.840 597.440 24.100 ;
        RECT 787.160 23.840 787.420 24.100 ;
      LAYER met2 ;
        RECT 786.700 1600.450 786.980 1604.000 ;
        RECT 786.700 1600.310 787.360 1600.450 ;
        RECT 786.700 1600.000 786.980 1600.310 ;
        RECT 787.220 24.130 787.360 1600.310 ;
        RECT 597.180 23.810 597.440 24.130 ;
        RECT 787.160 23.810 787.420 24.130 ;
        RECT 597.240 2.400 597.380 23.810 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 1591.440 620.930 1591.500 ;
        RECT 800.930 1591.440 801.250 1591.500 ;
        RECT 620.610 1591.300 801.250 1591.440 ;
        RECT 620.610 1591.240 620.930 1591.300 ;
        RECT 800.930 1591.240 801.250 1591.300 ;
        RECT 615.090 20.640 615.410 20.700 ;
        RECT 620.610 20.640 620.930 20.700 ;
        RECT 615.090 20.500 620.930 20.640 ;
        RECT 615.090 20.440 615.410 20.500 ;
        RECT 620.610 20.440 620.930 20.500 ;
      LAYER via ;
        RECT 620.640 1591.240 620.900 1591.500 ;
        RECT 800.960 1591.240 801.220 1591.500 ;
        RECT 615.120 20.440 615.380 20.700 ;
        RECT 620.640 20.440 620.900 20.700 ;
      LAYER met2 ;
        RECT 800.960 1600.000 801.240 1604.000 ;
        RECT 801.020 1591.530 801.160 1600.000 ;
        RECT 620.640 1591.210 620.900 1591.530 ;
        RECT 800.960 1591.210 801.220 1591.530 ;
        RECT 620.700 20.730 620.840 1591.210 ;
        RECT 615.120 20.410 615.380 20.730 ;
        RECT 620.640 20.410 620.900 20.730 ;
        RECT 615.180 2.400 615.320 20.410 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 26.080 110.330 26.140 ;
        RECT 386.470 26.080 386.790 26.140 ;
        RECT 110.010 25.940 386.790 26.080 ;
        RECT 110.010 25.880 110.330 25.940 ;
        RECT 386.470 25.880 386.790 25.940 ;
      LAYER via ;
        RECT 110.040 25.880 110.300 26.140 ;
        RECT 386.500 25.880 386.760 26.140 ;
      LAYER met2 ;
        RECT 389.260 1600.450 389.540 1604.000 ;
        RECT 386.560 1600.310 389.540 1600.450 ;
        RECT 386.560 26.170 386.700 1600.310 ;
        RECT 389.260 1600.000 389.540 1600.310 ;
        RECT 110.040 25.850 110.300 26.170 ;
        RECT 386.500 25.850 386.760 26.170 ;
        RECT 110.100 13.330 110.240 25.850 ;
        RECT 109.640 13.190 110.240 13.330 ;
        RECT 109.640 2.400 109.780 13.190 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 26.760 133.790 26.820 ;
        RECT 407.630 26.760 407.950 26.820 ;
        RECT 133.470 26.620 407.950 26.760 ;
        RECT 133.470 26.560 133.790 26.620 ;
        RECT 407.630 26.560 407.950 26.620 ;
      LAYER via ;
        RECT 133.500 26.560 133.760 26.820 ;
        RECT 407.660 26.560 407.920 26.820 ;
      LAYER met2 ;
        RECT 408.580 1600.450 408.860 1604.000 ;
        RECT 407.720 1600.310 408.860 1600.450 ;
        RECT 407.720 26.850 407.860 1600.310 ;
        RECT 408.580 1600.000 408.860 1600.310 ;
        RECT 133.500 26.530 133.760 26.850 ;
        RECT 407.660 26.530 407.920 26.850 ;
        RECT 133.560 2.400 133.700 26.530 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 26.420 151.730 26.480 ;
        RECT 420.970 26.420 421.290 26.480 ;
        RECT 151.410 26.280 421.290 26.420 ;
        RECT 151.410 26.220 151.730 26.280 ;
        RECT 420.970 26.220 421.290 26.280 ;
      LAYER via ;
        RECT 151.440 26.220 151.700 26.480 ;
        RECT 421.000 26.220 421.260 26.480 ;
      LAYER met2 ;
        RECT 423.300 1600.450 423.580 1604.000 ;
        RECT 421.060 1600.310 423.580 1600.450 ;
        RECT 421.060 26.510 421.200 1600.310 ;
        RECT 423.300 1600.000 423.580 1600.310 ;
        RECT 151.440 26.190 151.700 26.510 ;
        RECT 421.000 26.190 421.260 26.510 ;
        RECT 151.500 2.400 151.640 26.190 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 27.100 169.670 27.160 ;
        RECT 434.770 27.100 435.090 27.160 ;
        RECT 169.350 26.960 435.090 27.100 ;
        RECT 169.350 26.900 169.670 26.960 ;
        RECT 434.770 26.900 435.090 26.960 ;
      LAYER via ;
        RECT 169.380 26.900 169.640 27.160 ;
        RECT 434.800 26.900 435.060 27.160 ;
      LAYER met2 ;
        RECT 437.560 1600.450 437.840 1604.000 ;
        RECT 434.860 1600.310 437.840 1600.450 ;
        RECT 434.860 27.190 435.000 1600.310 ;
        RECT 437.560 1600.000 437.840 1600.310 ;
        RECT 169.380 26.870 169.640 27.190 ;
        RECT 434.800 26.870 435.060 27.190 ;
        RECT 169.440 2.400 169.580 26.870 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 27.440 187.150 27.500 ;
        RECT 448.570 27.440 448.890 27.500 ;
        RECT 186.830 27.300 448.890 27.440 ;
        RECT 186.830 27.240 187.150 27.300 ;
        RECT 448.570 27.240 448.890 27.300 ;
      LAYER via ;
        RECT 186.860 27.240 187.120 27.500 ;
        RECT 448.600 27.240 448.860 27.500 ;
      LAYER met2 ;
        RECT 452.280 1600.450 452.560 1604.000 ;
        RECT 448.660 1600.310 452.560 1600.450 ;
        RECT 448.660 27.530 448.800 1600.310 ;
        RECT 452.280 1600.000 452.560 1600.310 ;
        RECT 186.860 27.210 187.120 27.530 ;
        RECT 448.600 27.210 448.860 27.530 ;
        RECT 186.920 2.400 187.060 27.210 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 210.290 1593.820 210.610 1593.880 ;
        RECT 466.970 1593.820 467.290 1593.880 ;
        RECT 210.290 1593.680 467.290 1593.820 ;
        RECT 210.290 1593.620 210.610 1593.680 ;
        RECT 466.970 1593.620 467.290 1593.680 ;
        RECT 204.770 18.260 205.090 18.320 ;
        RECT 210.290 18.260 210.610 18.320 ;
        RECT 204.770 18.120 210.610 18.260 ;
        RECT 204.770 18.060 205.090 18.120 ;
        RECT 210.290 18.060 210.610 18.120 ;
      LAYER via ;
        RECT 210.320 1593.620 210.580 1593.880 ;
        RECT 467.000 1593.620 467.260 1593.880 ;
        RECT 204.800 18.060 205.060 18.320 ;
        RECT 210.320 18.060 210.580 18.320 ;
      LAYER met2 ;
        RECT 467.000 1600.000 467.280 1604.000 ;
        RECT 467.060 1593.910 467.200 1600.000 ;
        RECT 210.320 1593.590 210.580 1593.910 ;
        RECT 467.000 1593.590 467.260 1593.910 ;
        RECT 210.380 18.350 210.520 1593.590 ;
        RECT 204.800 18.030 205.060 18.350 ;
        RECT 210.320 18.030 210.580 18.350 ;
        RECT 204.860 2.400 205.000 18.030 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 447.725 1587.545 447.895 1590.095 ;
      LAYER mcon ;
        RECT 447.725 1589.925 447.895 1590.095 ;
      LAYER met1 ;
        RECT 447.665 1590.080 447.955 1590.125 ;
        RECT 481.230 1590.080 481.550 1590.140 ;
        RECT 447.665 1589.940 481.550 1590.080 ;
        RECT 447.665 1589.895 447.955 1589.940 ;
        RECT 481.230 1589.880 481.550 1589.940 ;
        RECT 389.690 1587.700 390.010 1587.760 ;
        RECT 447.665 1587.700 447.955 1587.745 ;
        RECT 389.690 1587.560 447.955 1587.700 ;
        RECT 389.690 1587.500 390.010 1587.560 ;
        RECT 447.665 1587.515 447.955 1587.560 ;
        RECT 222.710 15.540 223.030 15.600 ;
        RECT 389.690 15.540 390.010 15.600 ;
        RECT 222.710 15.400 390.010 15.540 ;
        RECT 222.710 15.340 223.030 15.400 ;
        RECT 389.690 15.340 390.010 15.400 ;
      LAYER via ;
        RECT 481.260 1589.880 481.520 1590.140 ;
        RECT 389.720 1587.500 389.980 1587.760 ;
        RECT 222.740 15.340 223.000 15.600 ;
        RECT 389.720 15.340 389.980 15.600 ;
      LAYER met2 ;
        RECT 481.260 1600.000 481.540 1604.000 ;
        RECT 481.320 1590.170 481.460 1600.000 ;
        RECT 481.260 1589.850 481.520 1590.170 ;
        RECT 389.720 1587.470 389.980 1587.790 ;
        RECT 389.780 15.630 389.920 1587.470 ;
        RECT 222.740 15.310 223.000 15.630 ;
        RECT 389.720 15.310 389.980 15.630 ;
        RECT 222.800 2.400 222.940 15.310 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 120.590 1588.040 120.910 1588.100 ;
        RECT 120.590 1587.900 296.540 1588.040 ;
        RECT 120.590 1587.840 120.910 1587.900 ;
        RECT 296.400 1587.700 296.540 1587.900 ;
        RECT 313.330 1587.700 313.650 1587.760 ;
        RECT 296.400 1587.560 313.650 1587.700 ;
        RECT 313.330 1587.500 313.650 1587.560 ;
        RECT 20.310 17.920 20.630 17.980 ;
        RECT 120.590 17.920 120.910 17.980 ;
        RECT 20.310 17.780 120.910 17.920 ;
        RECT 20.310 17.720 20.630 17.780 ;
        RECT 120.590 17.720 120.910 17.780 ;
      LAYER via ;
        RECT 120.620 1587.840 120.880 1588.100 ;
        RECT 313.360 1587.500 313.620 1587.760 ;
        RECT 20.340 17.720 20.600 17.980 ;
        RECT 120.620 17.720 120.880 17.980 ;
      LAYER met2 ;
        RECT 316.580 1600.450 316.860 1604.000 ;
        RECT 313.420 1600.310 316.860 1600.450 ;
        RECT 120.620 1587.810 120.880 1588.130 ;
        RECT 120.680 18.010 120.820 1587.810 ;
        RECT 313.420 1587.790 313.560 1600.310 ;
        RECT 316.580 1600.000 316.860 1600.310 ;
        RECT 313.360 1587.470 313.620 1587.790 ;
        RECT 20.340 17.690 20.600 18.010 ;
        RECT 120.620 17.690 120.880 18.010 ;
        RECT 20.400 2.400 20.540 17.690 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 1591.100 48.230 1591.160 ;
        RECT 335.870 1591.100 336.190 1591.160 ;
        RECT 47.910 1590.960 336.190 1591.100 ;
        RECT 47.910 1590.900 48.230 1590.960 ;
        RECT 335.870 1590.900 336.190 1590.960 ;
        RECT 44.230 17.580 44.550 17.640 ;
        RECT 47.910 17.580 48.230 17.640 ;
        RECT 44.230 17.440 48.230 17.580 ;
        RECT 44.230 17.380 44.550 17.440 ;
        RECT 47.910 17.380 48.230 17.440 ;
      LAYER via ;
        RECT 47.940 1590.900 48.200 1591.160 ;
        RECT 335.900 1590.900 336.160 1591.160 ;
        RECT 44.260 17.380 44.520 17.640 ;
        RECT 47.940 17.380 48.200 17.640 ;
      LAYER met2 ;
        RECT 335.900 1600.000 336.180 1604.000 ;
        RECT 335.960 1591.190 336.100 1600.000 ;
        RECT 47.940 1590.870 48.200 1591.190 ;
        RECT 335.900 1590.870 336.160 1591.190 ;
        RECT 48.000 17.670 48.140 1590.870 ;
        RECT 44.260 17.350 44.520 17.670 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 44.320 2.400 44.460 17.350 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 417.290 1593.480 417.610 1593.540 ;
        RECT 500.550 1593.480 500.870 1593.540 ;
        RECT 417.290 1593.340 477.320 1593.480 ;
        RECT 417.290 1593.280 417.610 1593.340 ;
        RECT 477.180 1593.140 477.320 1593.340 ;
        RECT 487.760 1593.340 500.870 1593.480 ;
        RECT 487.760 1593.140 487.900 1593.340 ;
        RECT 500.550 1593.280 500.870 1593.340 ;
        RECT 477.180 1593.000 487.900 1593.140 ;
        RECT 246.630 15.880 246.950 15.940 ;
        RECT 417.290 15.880 417.610 15.940 ;
        RECT 246.630 15.740 417.610 15.880 ;
        RECT 246.630 15.680 246.950 15.740 ;
        RECT 417.290 15.680 417.610 15.740 ;
      LAYER via ;
        RECT 417.320 1593.280 417.580 1593.540 ;
        RECT 500.580 1593.280 500.840 1593.540 ;
        RECT 246.660 15.680 246.920 15.940 ;
        RECT 417.320 15.680 417.580 15.940 ;
      LAYER met2 ;
        RECT 500.580 1600.000 500.860 1604.000 ;
        RECT 500.640 1593.570 500.780 1600.000 ;
        RECT 417.320 1593.250 417.580 1593.570 ;
        RECT 500.580 1593.250 500.840 1593.570 ;
        RECT 417.380 15.970 417.520 1593.250 ;
        RECT 246.660 15.650 246.920 15.970 ;
        RECT 417.320 15.650 417.580 15.970 ;
        RECT 246.720 2.400 246.860 15.650 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 462.445 1588.225 462.615 1589.075 ;
      LAYER mcon ;
        RECT 462.445 1588.905 462.615 1589.075 ;
      LAYER met1 ;
        RECT 515.270 1589.400 515.590 1589.460 ;
        RECT 472.580 1589.260 515.590 1589.400 ;
        RECT 462.385 1589.060 462.675 1589.105 ;
        RECT 472.580 1589.060 472.720 1589.260 ;
        RECT 515.270 1589.200 515.590 1589.260 ;
        RECT 462.385 1588.920 472.720 1589.060 ;
        RECT 462.385 1588.875 462.675 1588.920 ;
        RECT 268.710 1588.380 269.030 1588.440 ;
        RECT 462.385 1588.380 462.675 1588.425 ;
        RECT 268.710 1588.240 462.675 1588.380 ;
        RECT 268.710 1588.180 269.030 1588.240 ;
        RECT 462.385 1588.195 462.675 1588.240 ;
        RECT 264.110 18.260 264.430 18.320 ;
        RECT 268.710 18.260 269.030 18.320 ;
        RECT 264.110 18.120 269.030 18.260 ;
        RECT 264.110 18.060 264.430 18.120 ;
        RECT 268.710 18.060 269.030 18.120 ;
      LAYER via ;
        RECT 515.300 1589.200 515.560 1589.460 ;
        RECT 268.740 1588.180 269.000 1588.440 ;
        RECT 264.140 18.060 264.400 18.320 ;
        RECT 268.740 18.060 269.000 18.320 ;
      LAYER met2 ;
        RECT 515.300 1600.000 515.580 1604.000 ;
        RECT 515.360 1589.490 515.500 1600.000 ;
        RECT 515.300 1589.170 515.560 1589.490 ;
        RECT 268.740 1588.150 269.000 1588.470 ;
        RECT 268.800 18.350 268.940 1588.150 ;
        RECT 264.140 18.030 264.400 18.350 ;
        RECT 268.740 18.030 269.000 18.350 ;
        RECT 264.200 2.400 264.340 18.030 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 473.025 1588.905 473.195 1591.795 ;
      LAYER mcon ;
        RECT 473.025 1591.625 473.195 1591.795 ;
      LAYER met1 ;
        RECT 431.090 1591.780 431.410 1591.840 ;
        RECT 472.965 1591.780 473.255 1591.825 ;
        RECT 431.090 1591.640 473.255 1591.780 ;
        RECT 431.090 1591.580 431.410 1591.640 ;
        RECT 472.965 1591.595 473.255 1591.640 ;
        RECT 472.965 1589.060 473.255 1589.105 ;
        RECT 529.990 1589.060 530.310 1589.120 ;
        RECT 472.965 1588.920 530.310 1589.060 ;
        RECT 472.965 1588.875 473.255 1588.920 ;
        RECT 529.990 1588.860 530.310 1588.920 ;
        RECT 282.050 14.860 282.370 14.920 ;
        RECT 431.090 14.860 431.410 14.920 ;
        RECT 282.050 14.720 431.410 14.860 ;
        RECT 282.050 14.660 282.370 14.720 ;
        RECT 431.090 14.660 431.410 14.720 ;
      LAYER via ;
        RECT 431.120 1591.580 431.380 1591.840 ;
        RECT 530.020 1588.860 530.280 1589.120 ;
        RECT 282.080 14.660 282.340 14.920 ;
        RECT 431.120 14.660 431.380 14.920 ;
      LAYER met2 ;
        RECT 530.020 1600.000 530.300 1604.000 ;
        RECT 431.120 1591.550 431.380 1591.870 ;
        RECT 431.180 14.950 431.320 1591.550 ;
        RECT 530.080 1589.150 530.220 1600.000 ;
        RECT 530.020 1588.830 530.280 1589.150 ;
        RECT 282.080 14.630 282.340 14.950 ;
        RECT 431.120 14.630 431.380 14.950 ;
        RECT 282.140 2.400 282.280 14.630 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 472.105 1588.395 472.275 1589.415 ;
        RECT 472.105 1588.225 472.735 1588.395 ;
        RECT 485.905 1588.225 486.075 1594.175 ;
      LAYER mcon ;
        RECT 485.905 1594.005 486.075 1594.175 ;
        RECT 472.105 1589.245 472.275 1589.415 ;
        RECT 472.565 1588.225 472.735 1588.395 ;
      LAYER met1 ;
        RECT 485.845 1594.160 486.135 1594.205 ;
        RECT 485.845 1594.020 487.440 1594.160 ;
        RECT 485.845 1593.975 486.135 1594.020 ;
        RECT 487.300 1593.820 487.440 1594.020 ;
        RECT 542.870 1593.820 543.190 1593.880 ;
        RECT 487.300 1593.680 543.190 1593.820 ;
        RECT 542.870 1593.620 543.190 1593.680 ;
        RECT 458.690 1589.400 459.010 1589.460 ;
        RECT 472.045 1589.400 472.335 1589.445 ;
        RECT 458.690 1589.260 472.335 1589.400 ;
        RECT 458.690 1589.200 459.010 1589.260 ;
        RECT 472.045 1589.215 472.335 1589.260 ;
        RECT 472.505 1588.380 472.795 1588.425 ;
        RECT 485.845 1588.380 486.135 1588.425 ;
        RECT 472.505 1588.240 486.135 1588.380 ;
        RECT 472.505 1588.195 472.795 1588.240 ;
        RECT 485.845 1588.195 486.135 1588.240 ;
        RECT 299.990 15.200 300.310 15.260 ;
        RECT 458.690 15.200 459.010 15.260 ;
        RECT 299.990 15.060 459.010 15.200 ;
        RECT 299.990 15.000 300.310 15.060 ;
        RECT 458.690 15.000 459.010 15.060 ;
      LAYER via ;
        RECT 542.900 1593.620 543.160 1593.880 ;
        RECT 458.720 1589.200 458.980 1589.460 ;
        RECT 300.020 15.000 300.280 15.260 ;
        RECT 458.720 15.000 458.980 15.260 ;
      LAYER met2 ;
        RECT 544.280 1600.450 544.560 1604.000 ;
        RECT 542.960 1600.310 544.560 1600.450 ;
        RECT 542.960 1593.910 543.100 1600.310 ;
        RECT 544.280 1600.000 544.560 1600.310 ;
        RECT 542.900 1593.590 543.160 1593.910 ;
        RECT 458.720 1589.170 458.980 1589.490 ;
        RECT 458.780 15.290 458.920 1589.170 ;
        RECT 300.020 14.970 300.280 15.290 ;
        RECT 458.720 14.970 458.980 15.290 ;
        RECT 300.080 2.400 300.220 14.970 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 545.245 1590.775 545.415 1591.115 ;
        RECT 544.325 1590.605 545.415 1590.775 ;
        RECT 544.325 1589.245 544.495 1590.605 ;
      LAYER mcon ;
        RECT 545.245 1590.945 545.415 1591.115 ;
      LAYER met1 ;
        RECT 545.185 1591.100 545.475 1591.145 ;
        RECT 558.970 1591.100 559.290 1591.160 ;
        RECT 545.185 1590.960 559.290 1591.100 ;
        RECT 545.185 1590.915 545.475 1590.960 ;
        RECT 558.970 1590.900 559.290 1590.960 ;
        RECT 479.390 1589.740 479.710 1589.800 ;
        RECT 479.390 1589.600 521.020 1589.740 ;
        RECT 479.390 1589.540 479.710 1589.600 ;
        RECT 520.880 1589.400 521.020 1589.600 ;
        RECT 544.265 1589.400 544.555 1589.445 ;
        RECT 520.880 1589.260 544.555 1589.400 ;
        RECT 544.265 1589.215 544.555 1589.260 ;
        RECT 317.930 16.560 318.250 16.620 ;
        RECT 479.390 16.560 479.710 16.620 ;
        RECT 317.930 16.420 479.710 16.560 ;
        RECT 317.930 16.360 318.250 16.420 ;
        RECT 479.390 16.360 479.710 16.420 ;
      LAYER via ;
        RECT 559.000 1590.900 559.260 1591.160 ;
        RECT 479.420 1589.540 479.680 1589.800 ;
        RECT 317.960 16.360 318.220 16.620 ;
        RECT 479.420 16.360 479.680 16.620 ;
      LAYER met2 ;
        RECT 559.000 1600.000 559.280 1604.000 ;
        RECT 559.060 1591.190 559.200 1600.000 ;
        RECT 559.000 1590.870 559.260 1591.190 ;
        RECT 479.420 1589.510 479.680 1589.830 ;
        RECT 479.480 16.650 479.620 1589.510 ;
        RECT 317.960 16.330 318.220 16.650 ;
        RECT 479.420 16.330 479.680 16.650 ;
        RECT 318.020 2.400 318.160 16.330 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 507.065 1590.945 507.235 1593.495 ;
      LAYER mcon ;
        RECT 507.065 1593.325 507.235 1593.495 ;
      LAYER met1 ;
        RECT 573.230 1593.820 573.550 1593.880 ;
        RECT 543.420 1593.680 573.550 1593.820 ;
        RECT 507.005 1593.480 507.295 1593.525 ;
        RECT 543.420 1593.480 543.560 1593.680 ;
        RECT 573.230 1593.620 573.550 1593.680 ;
        RECT 507.005 1593.340 543.560 1593.480 ;
        RECT 507.005 1593.295 507.295 1593.340 ;
        RECT 337.710 1591.100 338.030 1591.160 ;
        RECT 507.005 1591.100 507.295 1591.145 ;
        RECT 337.710 1590.960 507.295 1591.100 ;
        RECT 337.710 1590.900 338.030 1590.960 ;
        RECT 507.005 1590.915 507.295 1590.960 ;
      LAYER via ;
        RECT 573.260 1593.620 573.520 1593.880 ;
        RECT 337.740 1590.900 338.000 1591.160 ;
      LAYER met2 ;
        RECT 573.260 1600.000 573.540 1604.000 ;
        RECT 573.320 1593.910 573.460 1600.000 ;
        RECT 573.260 1593.590 573.520 1593.910 ;
        RECT 337.740 1590.870 338.000 1591.190 ;
        RECT 337.800 3.130 337.940 1590.870 ;
        RECT 335.960 2.990 337.940 3.130 ;
        RECT 335.960 2.400 336.100 2.990 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 493.190 1590.080 493.510 1590.140 ;
        RECT 587.950 1590.080 588.270 1590.140 ;
        RECT 493.190 1589.940 588.270 1590.080 ;
        RECT 493.190 1589.880 493.510 1589.940 ;
        RECT 587.950 1589.880 588.270 1589.940 ;
        RECT 353.350 14.520 353.670 14.580 ;
        RECT 493.190 14.520 493.510 14.580 ;
        RECT 353.350 14.380 493.510 14.520 ;
        RECT 353.350 14.320 353.670 14.380 ;
        RECT 493.190 14.320 493.510 14.380 ;
      LAYER via ;
        RECT 493.220 1589.880 493.480 1590.140 ;
        RECT 587.980 1589.880 588.240 1590.140 ;
        RECT 353.380 14.320 353.640 14.580 ;
        RECT 493.220 14.320 493.480 14.580 ;
      LAYER met2 ;
        RECT 587.980 1600.000 588.260 1604.000 ;
        RECT 588.040 1590.170 588.180 1600.000 ;
        RECT 493.220 1589.850 493.480 1590.170 ;
        RECT 587.980 1589.850 588.240 1590.170 ;
        RECT 493.280 14.610 493.420 1589.850 ;
        RECT 353.380 14.290 353.640 14.610 ;
        RECT 493.220 14.290 493.480 14.610 ;
        RECT 353.440 2.400 353.580 14.290 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 1590.760 372.530 1590.820 ;
        RECT 602.670 1590.760 602.990 1590.820 ;
        RECT 372.210 1590.620 602.990 1590.760 ;
        RECT 372.210 1590.560 372.530 1590.620 ;
        RECT 602.670 1590.560 602.990 1590.620 ;
        RECT 371.290 2.960 371.610 3.020 ;
        RECT 372.210 2.960 372.530 3.020 ;
        RECT 371.290 2.820 372.530 2.960 ;
        RECT 371.290 2.760 371.610 2.820 ;
        RECT 372.210 2.760 372.530 2.820 ;
      LAYER via ;
        RECT 372.240 1590.560 372.500 1590.820 ;
        RECT 602.700 1590.560 602.960 1590.820 ;
        RECT 371.320 2.760 371.580 3.020 ;
        RECT 372.240 2.760 372.500 3.020 ;
      LAYER met2 ;
        RECT 602.700 1600.000 602.980 1604.000 ;
        RECT 602.760 1590.850 602.900 1600.000 ;
        RECT 372.240 1590.530 372.500 1590.850 ;
        RECT 602.700 1590.530 602.960 1590.850 ;
        RECT 372.300 3.050 372.440 1590.530 ;
        RECT 371.320 2.730 371.580 3.050 ;
        RECT 372.240 2.730 372.500 3.050 ;
        RECT 371.380 2.400 371.520 2.730 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.450 1591.100 507.770 1591.160 ;
        RECT 544.710 1591.100 545.030 1591.160 ;
        RECT 507.450 1590.960 545.030 1591.100 ;
        RECT 507.450 1590.900 507.770 1590.960 ;
        RECT 544.710 1590.900 545.030 1590.960 ;
        RECT 544.710 1589.400 545.030 1589.460 ;
        RECT 616.930 1589.400 617.250 1589.460 ;
        RECT 544.710 1589.260 617.250 1589.400 ;
        RECT 544.710 1589.200 545.030 1589.260 ;
        RECT 616.930 1589.200 617.250 1589.260 ;
        RECT 389.230 14.180 389.550 14.240 ;
        RECT 507.450 14.180 507.770 14.240 ;
        RECT 389.230 14.040 507.770 14.180 ;
        RECT 389.230 13.980 389.550 14.040 ;
        RECT 507.450 13.980 507.770 14.040 ;
      LAYER via ;
        RECT 507.480 1590.900 507.740 1591.160 ;
        RECT 544.740 1590.900 545.000 1591.160 ;
        RECT 544.740 1589.200 545.000 1589.460 ;
        RECT 616.960 1589.200 617.220 1589.460 ;
        RECT 389.260 13.980 389.520 14.240 ;
        RECT 507.480 13.980 507.740 14.240 ;
      LAYER met2 ;
        RECT 616.960 1600.000 617.240 1604.000 ;
        RECT 507.480 1590.870 507.740 1591.190 ;
        RECT 544.740 1590.870 545.000 1591.190 ;
        RECT 507.540 14.270 507.680 1590.870 ;
        RECT 544.800 1589.490 544.940 1590.870 ;
        RECT 617.020 1589.490 617.160 1600.000 ;
        RECT 544.740 1589.170 545.000 1589.490 ;
        RECT 616.960 1589.170 617.220 1589.490 ;
        RECT 389.260 13.950 389.520 14.270 ;
        RECT 507.480 13.950 507.740 14.270 ;
        RECT 389.320 2.400 389.460 13.950 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 520.865 1587.545 521.035 1588.395 ;
      LAYER mcon ;
        RECT 520.865 1588.225 521.035 1588.395 ;
      LAYER met1 ;
        RECT 486.290 1588.380 486.610 1588.440 ;
        RECT 520.805 1588.380 521.095 1588.425 ;
        RECT 486.290 1588.240 521.095 1588.380 ;
        RECT 486.290 1588.180 486.610 1588.240 ;
        RECT 520.805 1588.195 521.095 1588.240 ;
        RECT 631.650 1588.040 631.970 1588.100 ;
        RECT 622.540 1587.900 631.970 1588.040 ;
        RECT 520.805 1587.700 521.095 1587.745 ;
        RECT 622.540 1587.700 622.680 1587.900 ;
        RECT 631.650 1587.840 631.970 1587.900 ;
        RECT 520.805 1587.560 622.680 1587.700 ;
        RECT 520.805 1587.515 521.095 1587.560 ;
        RECT 407.170 19.280 407.490 19.340 ;
        RECT 486.290 19.280 486.610 19.340 ;
        RECT 407.170 19.140 486.610 19.280 ;
        RECT 407.170 19.080 407.490 19.140 ;
        RECT 486.290 19.080 486.610 19.140 ;
      LAYER via ;
        RECT 486.320 1588.180 486.580 1588.440 ;
        RECT 631.680 1587.840 631.940 1588.100 ;
        RECT 407.200 19.080 407.460 19.340 ;
        RECT 486.320 19.080 486.580 19.340 ;
      LAYER met2 ;
        RECT 631.680 1600.000 631.960 1604.000 ;
        RECT 486.320 1588.150 486.580 1588.470 ;
        RECT 486.380 19.370 486.520 1588.150 ;
        RECT 631.740 1588.130 631.880 1600.000 ;
        RECT 631.680 1587.810 631.940 1588.130 ;
        RECT 407.200 19.050 407.460 19.370 ;
        RECT 486.320 19.050 486.580 19.370 ;
        RECT 407.260 2.400 407.400 19.050 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 1590.760 68.470 1590.820 ;
        RECT 355.190 1590.760 355.510 1590.820 ;
        RECT 68.150 1590.620 355.510 1590.760 ;
        RECT 68.150 1590.560 68.470 1590.620 ;
        RECT 355.190 1590.560 355.510 1590.620 ;
      LAYER via ;
        RECT 68.180 1590.560 68.440 1590.820 ;
        RECT 355.220 1590.560 355.480 1590.820 ;
      LAYER met2 ;
        RECT 355.220 1600.000 355.500 1604.000 ;
        RECT 355.280 1590.850 355.420 1600.000 ;
        RECT 68.180 1590.530 68.440 1590.850 ;
        RECT 355.220 1590.530 355.480 1590.850 ;
        RECT 68.240 2.400 68.380 1590.530 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 506.990 1587.700 507.310 1587.760 ;
        RECT 506.990 1587.560 520.560 1587.700 ;
        RECT 506.990 1587.500 507.310 1587.560 ;
        RECT 520.420 1587.360 520.560 1587.560 ;
        RECT 645.910 1587.360 646.230 1587.420 ;
        RECT 520.420 1587.220 646.230 1587.360 ;
        RECT 645.910 1587.160 646.230 1587.220 ;
        RECT 424.650 15.880 424.970 15.940 ;
        RECT 506.990 15.880 507.310 15.940 ;
        RECT 424.650 15.740 507.310 15.880 ;
        RECT 424.650 15.680 424.970 15.740 ;
        RECT 506.990 15.680 507.310 15.740 ;
      LAYER via ;
        RECT 507.020 1587.500 507.280 1587.760 ;
        RECT 645.940 1587.160 646.200 1587.420 ;
        RECT 424.680 15.680 424.940 15.940 ;
        RECT 507.020 15.680 507.280 15.940 ;
      LAYER met2 ;
        RECT 645.940 1600.000 646.220 1604.000 ;
        RECT 507.020 1587.470 507.280 1587.790 ;
        RECT 507.080 15.970 507.220 1587.470 ;
        RECT 646.000 1587.450 646.140 1600.000 ;
        RECT 645.940 1587.130 646.200 1587.450 ;
        RECT 424.680 15.650 424.940 15.970 ;
        RECT 507.020 15.650 507.280 15.970 ;
        RECT 424.740 2.400 424.880 15.650 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 458.765 1587.545 458.935 1592.815 ;
        RECT 468.425 1592.645 468.595 1593.835 ;
        RECT 486.825 1591.625 486.995 1593.835 ;
      LAYER mcon ;
        RECT 468.425 1593.665 468.595 1593.835 ;
        RECT 458.765 1592.645 458.935 1592.815 ;
        RECT 486.825 1593.665 486.995 1593.835 ;
      LAYER met1 ;
        RECT 468.365 1593.820 468.655 1593.865 ;
        RECT 486.765 1593.820 487.055 1593.865 ;
        RECT 468.365 1593.680 487.055 1593.820 ;
        RECT 468.365 1593.635 468.655 1593.680 ;
        RECT 486.765 1593.635 487.055 1593.680 ;
        RECT 458.705 1592.800 458.995 1592.845 ;
        RECT 468.365 1592.800 468.655 1592.845 ;
        RECT 458.705 1592.660 468.655 1592.800 ;
        RECT 458.705 1592.615 458.995 1592.660 ;
        RECT 468.365 1592.615 468.655 1592.660 ;
        RECT 486.765 1591.780 487.055 1591.825 ;
        RECT 660.630 1591.780 660.950 1591.840 ;
        RECT 486.765 1591.640 660.950 1591.780 ;
        RECT 486.765 1591.595 487.055 1591.640 ;
        RECT 660.630 1591.580 660.950 1591.640 ;
        RECT 448.110 1587.700 448.430 1587.760 ;
        RECT 458.705 1587.700 458.995 1587.745 ;
        RECT 448.110 1587.560 458.995 1587.700 ;
        RECT 448.110 1587.500 448.430 1587.560 ;
        RECT 458.705 1587.515 458.995 1587.560 ;
        RECT 442.590 18.600 442.910 18.660 ;
        RECT 448.110 18.600 448.430 18.660 ;
        RECT 442.590 18.460 448.430 18.600 ;
        RECT 442.590 18.400 442.910 18.460 ;
        RECT 448.110 18.400 448.430 18.460 ;
      LAYER via ;
        RECT 660.660 1591.580 660.920 1591.840 ;
        RECT 448.140 1587.500 448.400 1587.760 ;
        RECT 442.620 18.400 442.880 18.660 ;
        RECT 448.140 18.400 448.400 18.660 ;
      LAYER met2 ;
        RECT 660.660 1600.000 660.940 1604.000 ;
        RECT 660.720 1591.870 660.860 1600.000 ;
        RECT 660.660 1591.550 660.920 1591.870 ;
        RECT 448.140 1587.470 448.400 1587.790 ;
        RECT 448.200 18.690 448.340 1587.470 ;
        RECT 442.620 18.370 442.880 18.690 ;
        RECT 448.140 18.370 448.400 18.690 ;
        RECT 442.680 2.400 442.820 18.370 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.690 1588.380 528.010 1588.440 ;
        RECT 675.350 1588.380 675.670 1588.440 ;
        RECT 527.690 1588.240 675.670 1588.380 ;
        RECT 527.690 1588.180 528.010 1588.240 ;
        RECT 675.350 1588.180 675.670 1588.240 ;
        RECT 460.530 19.620 460.850 19.680 ;
        RECT 527.690 19.620 528.010 19.680 ;
        RECT 460.530 19.480 528.010 19.620 ;
        RECT 460.530 19.420 460.850 19.480 ;
        RECT 527.690 19.420 528.010 19.480 ;
      LAYER via ;
        RECT 527.720 1588.180 527.980 1588.440 ;
        RECT 675.380 1588.180 675.640 1588.440 ;
        RECT 460.560 19.420 460.820 19.680 ;
        RECT 527.720 19.420 527.980 19.680 ;
      LAYER met2 ;
        RECT 675.380 1600.000 675.660 1604.000 ;
        RECT 675.440 1588.470 675.580 1600.000 ;
        RECT 527.720 1588.150 527.980 1588.470 ;
        RECT 675.380 1588.150 675.640 1588.470 ;
        RECT 527.780 19.710 527.920 1588.150 ;
        RECT 460.560 19.390 460.820 19.710 ;
        RECT 527.720 19.390 527.980 19.710 ;
        RECT 460.620 2.400 460.760 19.390 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 541.565 1592.985 544.955 1593.155 ;
        RECT 521.325 1586.865 521.495 1589.755 ;
        RECT 541.565 1589.585 541.735 1592.985 ;
      LAYER mcon ;
        RECT 544.785 1592.985 544.955 1593.155 ;
        RECT 521.325 1589.585 521.495 1589.755 ;
      LAYER met1 ;
        RECT 544.725 1593.140 545.015 1593.185 ;
        RECT 689.610 1593.140 689.930 1593.200 ;
        RECT 544.725 1593.000 689.930 1593.140 ;
        RECT 544.725 1592.955 545.015 1593.000 ;
        RECT 689.610 1592.940 689.930 1593.000 ;
        RECT 521.265 1589.740 521.555 1589.785 ;
        RECT 541.505 1589.740 541.795 1589.785 ;
        RECT 521.265 1589.600 541.795 1589.740 ;
        RECT 521.265 1589.555 521.555 1589.600 ;
        RECT 541.505 1589.555 541.795 1589.600 ;
        RECT 482.610 1587.360 482.930 1587.420 ;
        RECT 482.610 1587.220 513.660 1587.360 ;
        RECT 482.610 1587.160 482.930 1587.220 ;
        RECT 513.520 1587.020 513.660 1587.220 ;
        RECT 521.265 1587.020 521.555 1587.065 ;
        RECT 513.520 1586.880 521.555 1587.020 ;
        RECT 521.265 1586.835 521.555 1586.880 ;
        RECT 478.470 14.860 478.790 14.920 ;
        RECT 482.610 14.860 482.930 14.920 ;
        RECT 478.470 14.720 482.930 14.860 ;
        RECT 478.470 14.660 478.790 14.720 ;
        RECT 482.610 14.660 482.930 14.720 ;
      LAYER via ;
        RECT 689.640 1592.940 689.900 1593.200 ;
        RECT 482.640 1587.160 482.900 1587.420 ;
        RECT 478.500 14.660 478.760 14.920 ;
        RECT 482.640 14.660 482.900 14.920 ;
      LAYER met2 ;
        RECT 689.640 1600.000 689.920 1604.000 ;
        RECT 689.700 1593.230 689.840 1600.000 ;
        RECT 689.640 1592.910 689.900 1593.230 ;
        RECT 482.640 1587.130 482.900 1587.450 ;
        RECT 482.700 14.950 482.840 1587.130 ;
        RECT 478.500 14.630 478.760 14.950 ;
        RECT 482.640 14.630 482.900 14.950 ;
        RECT 478.560 2.400 478.700 14.630 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 679.105 1588.225 679.275 1589.075 ;
      LAYER mcon ;
        RECT 679.105 1588.905 679.275 1589.075 ;
      LAYER met1 ;
        RECT 541.490 1589.060 541.810 1589.120 ;
        RECT 679.045 1589.060 679.335 1589.105 ;
        RECT 541.490 1588.920 679.335 1589.060 ;
        RECT 541.490 1588.860 541.810 1588.920 ;
        RECT 679.045 1588.875 679.335 1588.920 ;
        RECT 679.045 1588.380 679.335 1588.425 ;
        RECT 704.330 1588.380 704.650 1588.440 ;
        RECT 679.045 1588.240 704.650 1588.380 ;
        RECT 679.045 1588.195 679.335 1588.240 ;
        RECT 704.330 1588.180 704.650 1588.240 ;
        RECT 496.410 20.640 496.730 20.700 ;
        RECT 541.490 20.640 541.810 20.700 ;
        RECT 496.410 20.500 541.810 20.640 ;
        RECT 496.410 20.440 496.730 20.500 ;
        RECT 541.490 20.440 541.810 20.500 ;
      LAYER via ;
        RECT 541.520 1588.860 541.780 1589.120 ;
        RECT 704.360 1588.180 704.620 1588.440 ;
        RECT 496.440 20.440 496.700 20.700 ;
        RECT 541.520 20.440 541.780 20.700 ;
      LAYER met2 ;
        RECT 704.360 1600.000 704.640 1604.000 ;
        RECT 541.520 1588.830 541.780 1589.150 ;
        RECT 541.580 20.730 541.720 1588.830 ;
        RECT 704.420 1588.470 704.560 1600.000 ;
        RECT 704.360 1588.150 704.620 1588.470 ;
        RECT 496.440 20.410 496.700 20.730 ;
        RECT 541.520 20.410 541.780 20.730 ;
        RECT 496.500 2.400 496.640 20.410 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 541.950 1589.740 542.270 1589.800 ;
        RECT 718.590 1589.740 718.910 1589.800 ;
        RECT 541.950 1589.600 718.910 1589.740 ;
        RECT 541.950 1589.540 542.270 1589.600 ;
        RECT 718.590 1589.540 718.910 1589.600 ;
        RECT 513.890 15.200 514.210 15.260 ;
        RECT 541.950 15.200 542.270 15.260 ;
        RECT 513.890 15.060 542.270 15.200 ;
        RECT 513.890 15.000 514.210 15.060 ;
        RECT 541.950 15.000 542.270 15.060 ;
      LAYER via ;
        RECT 541.980 1589.540 542.240 1589.800 ;
        RECT 718.620 1589.540 718.880 1589.800 ;
        RECT 513.920 15.000 514.180 15.260 ;
        RECT 541.980 15.000 542.240 15.260 ;
      LAYER met2 ;
        RECT 718.620 1600.000 718.900 1604.000 ;
        RECT 718.680 1589.830 718.820 1600.000 ;
        RECT 541.980 1589.510 542.240 1589.830 ;
        RECT 718.620 1589.510 718.880 1589.830 ;
        RECT 542.040 15.290 542.180 1589.510 ;
        RECT 513.920 14.970 514.180 15.290 ;
        RECT 541.980 14.970 542.240 15.290 ;
        RECT 513.980 2.400 514.120 14.970 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 575.990 1588.720 576.310 1588.780 ;
        RECT 575.990 1588.580 713.760 1588.720 ;
        RECT 575.990 1588.520 576.310 1588.580 ;
        RECT 713.620 1588.380 713.760 1588.580 ;
        RECT 733.310 1588.380 733.630 1588.440 ;
        RECT 713.620 1588.240 733.630 1588.380 ;
        RECT 733.310 1588.180 733.630 1588.240 ;
        RECT 531.830 18.260 532.150 18.320 ;
        RECT 575.990 18.260 576.310 18.320 ;
        RECT 531.830 18.120 576.310 18.260 ;
        RECT 531.830 18.060 532.150 18.120 ;
        RECT 575.990 18.060 576.310 18.120 ;
      LAYER via ;
        RECT 576.020 1588.520 576.280 1588.780 ;
        RECT 733.340 1588.180 733.600 1588.440 ;
        RECT 531.860 18.060 532.120 18.320 ;
        RECT 576.020 18.060 576.280 18.320 ;
      LAYER met2 ;
        RECT 733.340 1600.000 733.620 1604.000 ;
        RECT 576.020 1588.490 576.280 1588.810 ;
        RECT 576.080 18.350 576.220 1588.490 ;
        RECT 733.400 1588.470 733.540 1600.000 ;
        RECT 733.340 1588.150 733.600 1588.470 ;
        RECT 531.860 18.030 532.120 18.350 ;
        RECT 576.020 18.030 576.280 18.350 ;
        RECT 531.920 2.400 532.060 18.030 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 707.090 1591.780 707.410 1591.840 ;
        RECT 748.030 1591.780 748.350 1591.840 ;
        RECT 707.090 1591.640 748.350 1591.780 ;
        RECT 707.090 1591.580 707.410 1591.640 ;
        RECT 748.030 1591.580 748.350 1591.640 ;
        RECT 549.770 16.220 550.090 16.280 ;
        RECT 707.090 16.220 707.410 16.280 ;
        RECT 549.770 16.080 707.410 16.220 ;
        RECT 549.770 16.020 550.090 16.080 ;
        RECT 707.090 16.020 707.410 16.080 ;
      LAYER via ;
        RECT 707.120 1591.580 707.380 1591.840 ;
        RECT 748.060 1591.580 748.320 1591.840 ;
        RECT 549.800 16.020 550.060 16.280 ;
        RECT 707.120 16.020 707.380 16.280 ;
      LAYER met2 ;
        RECT 748.060 1600.000 748.340 1604.000 ;
        RECT 748.120 1591.870 748.260 1600.000 ;
        RECT 707.120 1591.550 707.380 1591.870 ;
        RECT 748.060 1591.550 748.320 1591.870 ;
        RECT 707.180 16.310 707.320 1591.550 ;
        RECT 549.800 15.990 550.060 16.310 ;
        RECT 707.120 15.990 707.380 16.310 ;
        RECT 549.860 2.400 550.000 15.990 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 621.145 15.045 621.315 20.655 ;
      LAYER mcon ;
        RECT 621.145 20.485 621.315 20.655 ;
      LAYER met1 ;
        RECT 762.290 1588.040 762.610 1588.100 ;
        RECT 750.420 1587.900 762.610 1588.040 ;
        RECT 734.690 1587.360 735.010 1587.420 ;
        RECT 750.420 1587.360 750.560 1587.900 ;
        RECT 762.290 1587.840 762.610 1587.900 ;
        RECT 734.690 1587.220 750.560 1587.360 ;
        RECT 734.690 1587.160 735.010 1587.220 ;
        RECT 621.085 20.640 621.375 20.685 ;
        RECT 734.690 20.640 735.010 20.700 ;
        RECT 621.085 20.500 735.010 20.640 ;
        RECT 621.085 20.455 621.375 20.500 ;
        RECT 734.690 20.440 735.010 20.500 ;
        RECT 567.710 15.200 568.030 15.260 ;
        RECT 621.085 15.200 621.375 15.245 ;
        RECT 567.710 15.060 621.375 15.200 ;
        RECT 567.710 15.000 568.030 15.060 ;
        RECT 621.085 15.015 621.375 15.060 ;
      LAYER via ;
        RECT 734.720 1587.160 734.980 1587.420 ;
        RECT 762.320 1587.840 762.580 1588.100 ;
        RECT 734.720 20.440 734.980 20.700 ;
        RECT 567.740 15.000 568.000 15.260 ;
      LAYER met2 ;
        RECT 762.320 1600.000 762.600 1604.000 ;
        RECT 762.380 1588.130 762.520 1600.000 ;
        RECT 762.320 1587.810 762.580 1588.130 ;
        RECT 734.720 1587.130 734.980 1587.450 ;
        RECT 734.780 20.730 734.920 1587.130 ;
        RECT 734.720 20.410 734.980 20.730 ;
        RECT 567.740 14.970 568.000 15.290 ;
        RECT 567.800 2.400 567.940 14.970 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 593.010 1591.100 593.330 1591.160 ;
        RECT 777.010 1591.100 777.330 1591.160 ;
        RECT 593.010 1590.960 777.330 1591.100 ;
        RECT 593.010 1590.900 593.330 1590.960 ;
        RECT 777.010 1590.900 777.330 1590.960 ;
        RECT 589.790 1590.080 590.110 1590.140 ;
        RECT 593.010 1590.080 593.330 1590.140 ;
        RECT 589.790 1589.940 593.330 1590.080 ;
        RECT 589.790 1589.880 590.110 1589.940 ;
        RECT 593.010 1589.880 593.330 1589.940 ;
        RECT 585.650 16.900 585.970 16.960 ;
        RECT 589.790 16.900 590.110 16.960 ;
        RECT 585.650 16.760 590.110 16.900 ;
        RECT 585.650 16.700 585.970 16.760 ;
        RECT 589.790 16.700 590.110 16.760 ;
      LAYER via ;
        RECT 593.040 1590.900 593.300 1591.160 ;
        RECT 777.040 1590.900 777.300 1591.160 ;
        RECT 589.820 1589.880 590.080 1590.140 ;
        RECT 593.040 1589.880 593.300 1590.140 ;
        RECT 585.680 16.700 585.940 16.960 ;
        RECT 589.820 16.700 590.080 16.960 ;
      LAYER met2 ;
        RECT 777.040 1600.000 777.320 1604.000 ;
        RECT 777.100 1591.190 777.240 1600.000 ;
        RECT 593.040 1590.870 593.300 1591.190 ;
        RECT 777.040 1590.870 777.300 1591.190 ;
        RECT 593.100 1590.170 593.240 1590.870 ;
        RECT 589.820 1589.850 590.080 1590.170 ;
        RECT 593.040 1589.850 593.300 1590.170 ;
        RECT 589.880 16.990 590.020 1589.850 ;
        RECT 585.680 16.670 585.940 16.990 ;
        RECT 589.820 16.670 590.080 16.990 ;
        RECT 585.740 2.400 585.880 16.670 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 327.665 1587.205 328.755 1587.375 ;
      LAYER mcon ;
        RECT 328.585 1587.205 328.755 1587.375 ;
      LAYER met1 ;
        RECT 314.250 1587.360 314.570 1587.420 ;
        RECT 327.605 1587.360 327.895 1587.405 ;
        RECT 314.250 1587.220 327.895 1587.360 ;
        RECT 314.250 1587.160 314.570 1587.220 ;
        RECT 327.605 1587.175 327.895 1587.220 ;
        RECT 328.525 1587.360 328.815 1587.405 ;
        RECT 374.510 1587.360 374.830 1587.420 ;
        RECT 328.525 1587.220 374.830 1587.360 ;
        RECT 328.525 1587.175 328.815 1587.220 ;
        RECT 374.510 1587.160 374.830 1587.220 ;
        RECT 91.610 16.560 91.930 16.620 ;
        RECT 314.250 16.560 314.570 16.620 ;
        RECT 91.610 16.420 314.570 16.560 ;
        RECT 91.610 16.360 91.930 16.420 ;
        RECT 314.250 16.360 314.570 16.420 ;
      LAYER via ;
        RECT 314.280 1587.160 314.540 1587.420 ;
        RECT 374.540 1587.160 374.800 1587.420 ;
        RECT 91.640 16.360 91.900 16.620 ;
        RECT 314.280 16.360 314.540 16.620 ;
      LAYER met2 ;
        RECT 374.540 1600.000 374.820 1604.000 ;
        RECT 374.600 1587.450 374.740 1600.000 ;
        RECT 314.280 1587.130 314.540 1587.450 ;
        RECT 374.540 1587.130 374.800 1587.450 ;
        RECT 314.340 16.650 314.480 1587.130 ;
        RECT 91.640 16.330 91.900 16.650 ;
        RECT 314.280 16.330 314.540 16.650 ;
        RECT 91.700 2.400 91.840 16.330 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 1590.080 607.130 1590.140 ;
        RECT 791.270 1590.080 791.590 1590.140 ;
        RECT 606.810 1589.940 791.590 1590.080 ;
        RECT 606.810 1589.880 607.130 1589.940 ;
        RECT 791.270 1589.880 791.590 1589.940 ;
        RECT 603.130 20.640 603.450 20.700 ;
        RECT 606.810 20.640 607.130 20.700 ;
        RECT 603.130 20.500 607.130 20.640 ;
        RECT 603.130 20.440 603.450 20.500 ;
        RECT 606.810 20.440 607.130 20.500 ;
      LAYER via ;
        RECT 606.840 1589.880 607.100 1590.140 ;
        RECT 791.300 1589.880 791.560 1590.140 ;
        RECT 603.160 20.440 603.420 20.700 ;
        RECT 606.840 20.440 607.100 20.700 ;
      LAYER met2 ;
        RECT 791.300 1600.000 791.580 1604.000 ;
        RECT 791.360 1590.170 791.500 1600.000 ;
        RECT 606.840 1589.850 607.100 1590.170 ;
        RECT 791.300 1589.850 791.560 1590.170 ;
        RECT 606.900 20.730 607.040 1589.850 ;
        RECT 603.160 20.410 603.420 20.730 ;
        RECT 606.840 20.410 607.100 20.730 ;
        RECT 603.220 2.400 603.360 20.410 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.510 1589.400 627.830 1589.460 ;
        RECT 805.990 1589.400 806.310 1589.460 ;
        RECT 627.510 1589.260 806.310 1589.400 ;
        RECT 627.510 1589.200 627.830 1589.260 ;
        RECT 805.990 1589.200 806.310 1589.260 ;
        RECT 621.070 17.920 621.390 17.980 ;
        RECT 627.510 17.920 627.830 17.980 ;
        RECT 621.070 17.780 627.830 17.920 ;
        RECT 621.070 17.720 621.390 17.780 ;
        RECT 627.510 17.720 627.830 17.780 ;
      LAYER via ;
        RECT 627.540 1589.200 627.800 1589.460 ;
        RECT 806.020 1589.200 806.280 1589.460 ;
        RECT 621.100 17.720 621.360 17.980 ;
        RECT 627.540 17.720 627.800 17.980 ;
      LAYER met2 ;
        RECT 806.020 1600.000 806.300 1604.000 ;
        RECT 806.080 1589.490 806.220 1600.000 ;
        RECT 627.540 1589.170 627.800 1589.490 ;
        RECT 806.020 1589.170 806.280 1589.490 ;
        RECT 627.600 18.010 627.740 1589.170 ;
        RECT 621.100 17.690 621.360 18.010 ;
        RECT 627.540 17.690 627.800 18.010 ;
        RECT 621.160 2.400 621.300 17.690 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 141.290 1593.480 141.610 1593.540 ;
        RECT 394.290 1593.480 394.610 1593.540 ;
        RECT 141.290 1593.340 394.610 1593.480 ;
        RECT 141.290 1593.280 141.610 1593.340 ;
        RECT 394.290 1593.280 394.610 1593.340 ;
        RECT 115.530 20.640 115.850 20.700 ;
        RECT 141.290 20.640 141.610 20.700 ;
        RECT 115.530 20.500 141.610 20.640 ;
        RECT 115.530 20.440 115.850 20.500 ;
        RECT 141.290 20.440 141.610 20.500 ;
      LAYER via ;
        RECT 141.320 1593.280 141.580 1593.540 ;
        RECT 394.320 1593.280 394.580 1593.540 ;
        RECT 115.560 20.440 115.820 20.700 ;
        RECT 141.320 20.440 141.580 20.700 ;
      LAYER met2 ;
        RECT 394.320 1600.000 394.600 1604.000 ;
        RECT 394.380 1593.570 394.520 1600.000 ;
        RECT 141.320 1593.250 141.580 1593.570 ;
        RECT 394.320 1593.250 394.580 1593.570 ;
        RECT 141.380 20.730 141.520 1593.250 ;
        RECT 115.560 20.410 115.820 20.730 ;
        RECT 141.320 20.410 141.580 20.730 ;
        RECT 115.620 2.400 115.760 20.410 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 396.590 1590.080 396.910 1590.140 ;
        RECT 413.610 1590.080 413.930 1590.140 ;
        RECT 396.590 1589.940 413.930 1590.080 ;
        RECT 396.590 1589.880 396.910 1589.940 ;
        RECT 413.610 1589.880 413.930 1589.940 ;
        RECT 139.450 18.260 139.770 18.320 ;
        RECT 139.450 18.120 162.680 18.260 ;
        RECT 139.450 18.060 139.770 18.120 ;
        RECT 162.540 17.920 162.680 18.120 ;
        RECT 396.590 17.920 396.910 17.980 ;
        RECT 162.540 17.780 396.910 17.920 ;
        RECT 396.590 17.720 396.910 17.780 ;
      LAYER via ;
        RECT 396.620 1589.880 396.880 1590.140 ;
        RECT 413.640 1589.880 413.900 1590.140 ;
        RECT 139.480 18.060 139.740 18.320 ;
        RECT 396.620 17.720 396.880 17.980 ;
      LAYER met2 ;
        RECT 413.640 1600.000 413.920 1604.000 ;
        RECT 413.700 1590.170 413.840 1600.000 ;
        RECT 396.620 1589.850 396.880 1590.170 ;
        RECT 413.640 1589.850 413.900 1590.170 ;
        RECT 139.480 18.030 139.740 18.350 ;
        RECT 139.540 2.400 139.680 18.030 ;
        RECT 396.680 18.010 396.820 1589.850 ;
        RECT 396.620 17.690 396.880 18.010 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 1591.780 158.630 1591.840 ;
        RECT 427.870 1591.780 428.190 1591.840 ;
        RECT 158.310 1591.640 428.190 1591.780 ;
        RECT 158.310 1591.580 158.630 1591.640 ;
        RECT 427.870 1591.580 428.190 1591.640 ;
      LAYER via ;
        RECT 158.340 1591.580 158.600 1591.840 ;
        RECT 427.900 1591.580 428.160 1591.840 ;
      LAYER met2 ;
        RECT 427.900 1600.000 428.180 1604.000 ;
        RECT 427.960 1591.870 428.100 1600.000 ;
        RECT 158.340 1591.550 158.600 1591.870 ;
        RECT 427.900 1591.550 428.160 1591.870 ;
        RECT 158.400 16.900 158.540 1591.550 ;
        RECT 157.480 16.760 158.540 16.900 ;
        RECT 157.480 2.400 157.620 16.760 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 410.390 1592.460 410.710 1592.520 ;
        RECT 442.590 1592.460 442.910 1592.520 ;
        RECT 410.390 1592.320 442.910 1592.460 ;
        RECT 410.390 1592.260 410.710 1592.320 ;
        RECT 442.590 1592.260 442.910 1592.320 ;
        RECT 174.870 20.300 175.190 20.360 ;
        RECT 410.390 20.300 410.710 20.360 ;
        RECT 174.870 20.160 410.710 20.300 ;
        RECT 174.870 20.100 175.190 20.160 ;
        RECT 410.390 20.100 410.710 20.160 ;
      LAYER via ;
        RECT 410.420 1592.260 410.680 1592.520 ;
        RECT 442.620 1592.260 442.880 1592.520 ;
        RECT 174.900 20.100 175.160 20.360 ;
        RECT 410.420 20.100 410.680 20.360 ;
      LAYER met2 ;
        RECT 442.620 1600.000 442.900 1604.000 ;
        RECT 442.680 1592.550 442.820 1600.000 ;
        RECT 410.420 1592.230 410.680 1592.550 ;
        RECT 442.620 1592.230 442.880 1592.550 ;
        RECT 410.480 20.390 410.620 1592.230 ;
        RECT 174.900 20.070 175.160 20.390 ;
        RECT 410.420 20.070 410.680 20.390 ;
        RECT 174.960 2.400 175.100 20.070 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.350 1592.800 192.670 1592.860 ;
        RECT 457.310 1592.800 457.630 1592.860 ;
        RECT 192.350 1592.660 457.630 1592.800 ;
        RECT 192.350 1592.600 192.670 1592.660 ;
        RECT 457.310 1592.600 457.630 1592.660 ;
      LAYER via ;
        RECT 192.380 1592.600 192.640 1592.860 ;
        RECT 457.340 1592.600 457.600 1592.860 ;
      LAYER met2 ;
        RECT 457.340 1600.000 457.620 1604.000 ;
        RECT 457.400 1592.890 457.540 1600.000 ;
        RECT 192.380 1592.570 192.640 1592.890 ;
        RECT 457.340 1592.570 457.600 1592.890 ;
        RECT 192.440 17.410 192.580 1592.570 ;
        RECT 192.440 17.270 193.040 17.410 ;
        RECT 192.900 2.400 193.040 17.270 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 276.145 14.025 276.315 20.655 ;
        RECT 345.145 14.025 345.315 20.655 ;
        RECT 372.745 19.805 372.915 20.655 ;
      LAYER mcon ;
        RECT 276.145 20.485 276.315 20.655 ;
        RECT 345.145 20.485 345.315 20.655 ;
        RECT 372.745 20.485 372.915 20.655 ;
      LAYER met1 ;
        RECT 444.890 1587.360 445.210 1587.420 ;
        RECT 471.570 1587.360 471.890 1587.420 ;
        RECT 444.890 1587.220 471.890 1587.360 ;
        RECT 444.890 1587.160 445.210 1587.220 ;
        RECT 471.570 1587.160 471.890 1587.220 ;
        RECT 210.750 20.640 211.070 20.700 ;
        RECT 276.085 20.640 276.375 20.685 ;
        RECT 210.750 20.500 276.375 20.640 ;
        RECT 210.750 20.440 211.070 20.500 ;
        RECT 276.085 20.455 276.375 20.500 ;
        RECT 345.085 20.640 345.375 20.685 ;
        RECT 372.685 20.640 372.975 20.685 ;
        RECT 345.085 20.500 372.975 20.640 ;
        RECT 345.085 20.455 345.375 20.500 ;
        RECT 372.685 20.455 372.975 20.500 ;
        RECT 372.685 19.960 372.975 20.005 ;
        RECT 444.890 19.960 445.210 20.020 ;
        RECT 372.685 19.820 445.210 19.960 ;
        RECT 372.685 19.775 372.975 19.820 ;
        RECT 444.890 19.760 445.210 19.820 ;
        RECT 276.085 14.180 276.375 14.225 ;
        RECT 345.085 14.180 345.375 14.225 ;
        RECT 276.085 14.040 345.375 14.180 ;
        RECT 276.085 13.995 276.375 14.040 ;
        RECT 345.085 13.995 345.375 14.040 ;
      LAYER via ;
        RECT 444.920 1587.160 445.180 1587.420 ;
        RECT 471.600 1587.160 471.860 1587.420 ;
        RECT 210.780 20.440 211.040 20.700 ;
        RECT 444.920 19.760 445.180 20.020 ;
      LAYER met2 ;
        RECT 471.600 1600.000 471.880 1604.000 ;
        RECT 471.660 1587.450 471.800 1600.000 ;
        RECT 444.920 1587.130 445.180 1587.450 ;
        RECT 471.600 1587.130 471.860 1587.450 ;
        RECT 210.780 20.410 211.040 20.730 ;
        RECT 210.840 2.400 210.980 20.410 ;
        RECT 444.980 20.050 445.120 1587.130 ;
        RECT 444.920 19.730 445.180 20.050 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 473.485 1589.585 473.655 1591.795 ;
      LAYER mcon ;
        RECT 473.485 1591.625 473.655 1591.795 ;
      LAYER met1 ;
        RECT 473.425 1591.780 473.715 1591.825 ;
        RECT 486.290 1591.780 486.610 1591.840 ;
        RECT 473.425 1591.640 486.610 1591.780 ;
        RECT 473.425 1591.595 473.715 1591.640 ;
        RECT 486.290 1591.580 486.610 1591.640 ;
        RECT 473.425 1589.740 473.715 1589.785 ;
        RECT 458.320 1589.600 473.715 1589.740 ;
        RECT 234.210 1589.400 234.530 1589.460 ;
        RECT 458.320 1589.400 458.460 1589.600 ;
        RECT 473.425 1589.555 473.715 1589.600 ;
        RECT 234.210 1589.260 458.460 1589.400 ;
        RECT 234.210 1589.200 234.530 1589.260 ;
        RECT 228.690 18.260 229.010 18.320 ;
        RECT 234.210 18.260 234.530 18.320 ;
        RECT 228.690 18.120 234.530 18.260 ;
        RECT 228.690 18.060 229.010 18.120 ;
        RECT 234.210 18.060 234.530 18.120 ;
      LAYER via ;
        RECT 486.320 1591.580 486.580 1591.840 ;
        RECT 234.240 1589.200 234.500 1589.460 ;
        RECT 228.720 18.060 228.980 18.320 ;
        RECT 234.240 18.060 234.500 18.320 ;
      LAYER met2 ;
        RECT 486.320 1600.000 486.600 1604.000 ;
        RECT 486.380 1591.870 486.520 1600.000 ;
        RECT 486.320 1591.550 486.580 1591.870 ;
        RECT 234.240 1589.170 234.500 1589.490 ;
        RECT 234.300 18.350 234.440 1589.170 ;
        RECT 228.720 18.030 228.980 18.350 ;
        RECT 234.240 18.030 234.500 18.350 ;
        RECT 228.780 2.400 228.920 18.030 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 179.545 15.725 179.715 17.595 ;
        RECT 295.005 16.745 295.175 17.595 ;
      LAYER mcon ;
        RECT 179.545 17.425 179.715 17.595 ;
        RECT 295.005 17.425 295.175 17.595 ;
      LAYER met1 ;
        RECT 313.790 1589.060 314.110 1589.120 ;
        RECT 340.930 1589.060 341.250 1589.120 ;
        RECT 313.790 1588.920 341.250 1589.060 ;
        RECT 313.790 1588.860 314.110 1588.920 ;
        RECT 340.930 1588.860 341.250 1588.920 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 179.485 17.580 179.775 17.625 ;
        RECT 50.210 17.440 179.775 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 179.485 17.395 179.775 17.440 ;
        RECT 227.310 17.580 227.630 17.640 ;
        RECT 294.945 17.580 295.235 17.625 ;
        RECT 227.310 17.440 295.235 17.580 ;
        RECT 227.310 17.380 227.630 17.440 ;
        RECT 294.945 17.395 295.235 17.440 ;
        RECT 294.945 16.900 295.235 16.945 ;
        RECT 313.790 16.900 314.110 16.960 ;
        RECT 294.945 16.760 314.110 16.900 ;
        RECT 294.945 16.715 295.235 16.760 ;
        RECT 313.790 16.700 314.110 16.760 ;
        RECT 179.485 15.880 179.775 15.925 ;
        RECT 226.850 15.880 227.170 15.940 ;
        RECT 179.485 15.740 227.170 15.880 ;
        RECT 179.485 15.695 179.775 15.740 ;
        RECT 226.850 15.680 227.170 15.740 ;
      LAYER via ;
        RECT 313.820 1588.860 314.080 1589.120 ;
        RECT 340.960 1588.860 341.220 1589.120 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 227.340 17.380 227.600 17.640 ;
        RECT 313.820 16.700 314.080 16.960 ;
        RECT 226.880 15.680 227.140 15.940 ;
      LAYER met2 ;
        RECT 340.960 1600.000 341.240 1604.000 ;
        RECT 341.020 1589.150 341.160 1600.000 ;
        RECT 313.820 1588.830 314.080 1589.150 ;
        RECT 340.960 1588.830 341.220 1589.150 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 227.340 17.350 227.600 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 227.400 16.730 227.540 17.350 ;
        RECT 313.880 16.990 314.020 1588.830 ;
        RECT 226.940 16.590 227.540 16.730 ;
        RECT 313.820 16.670 314.080 16.990 ;
        RECT 226.940 15.970 227.080 16.590 ;
        RECT 226.880 15.650 227.140 15.970 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 276.145 1587.205 276.315 1589.755 ;
        RECT 299.605 1587.205 299.775 1588.055 ;
        RECT 327.665 1587.885 327.835 1589.755 ;
        RECT 372.745 1586.865 372.915 1589.755 ;
        RECT 414.145 1587.205 414.315 1590.095 ;
        RECT 423.805 1587.205 423.975 1590.095 ;
        RECT 481.765 1587.205 481.935 1590.095 ;
        RECT 488.205 1589.925 488.375 1593.155 ;
      LAYER mcon ;
        RECT 488.205 1592.985 488.375 1593.155 ;
        RECT 414.145 1589.925 414.315 1590.095 ;
        RECT 276.145 1589.585 276.315 1589.755 ;
        RECT 327.665 1589.585 327.835 1589.755 ;
        RECT 299.605 1587.885 299.775 1588.055 ;
        RECT 372.745 1589.585 372.915 1589.755 ;
        RECT 423.805 1589.925 423.975 1590.095 ;
        RECT 481.765 1589.925 481.935 1590.095 ;
      LAYER met1 ;
        RECT 488.145 1593.140 488.435 1593.185 ;
        RECT 505.610 1593.140 505.930 1593.200 ;
        RECT 488.145 1593.000 505.930 1593.140 ;
        RECT 488.145 1592.955 488.435 1593.000 ;
        RECT 505.610 1592.940 505.930 1593.000 ;
        RECT 414.085 1590.080 414.375 1590.125 ;
        RECT 423.745 1590.080 424.035 1590.125 ;
        RECT 414.085 1589.940 424.035 1590.080 ;
        RECT 414.085 1589.895 414.375 1589.940 ;
        RECT 423.745 1589.895 424.035 1589.940 ;
        RECT 481.705 1590.080 481.995 1590.125 ;
        RECT 488.145 1590.080 488.435 1590.125 ;
        RECT 481.705 1589.940 488.435 1590.080 ;
        RECT 481.705 1589.895 481.995 1589.940 ;
        RECT 488.145 1589.895 488.435 1589.940 ;
        RECT 254.910 1589.740 255.230 1589.800 ;
        RECT 276.085 1589.740 276.375 1589.785 ;
        RECT 254.910 1589.600 276.375 1589.740 ;
        RECT 254.910 1589.540 255.230 1589.600 ;
        RECT 276.085 1589.555 276.375 1589.600 ;
        RECT 327.605 1589.740 327.895 1589.785 ;
        RECT 372.685 1589.740 372.975 1589.785 ;
        RECT 327.605 1589.600 372.975 1589.740 ;
        RECT 327.605 1589.555 327.895 1589.600 ;
        RECT 372.685 1589.555 372.975 1589.600 ;
        RECT 299.545 1588.040 299.835 1588.085 ;
        RECT 327.605 1588.040 327.895 1588.085 ;
        RECT 299.545 1587.900 327.895 1588.040 ;
        RECT 299.545 1587.855 299.835 1587.900 ;
        RECT 327.605 1587.855 327.895 1587.900 ;
        RECT 276.085 1587.360 276.375 1587.405 ;
        RECT 299.545 1587.360 299.835 1587.405 ;
        RECT 414.085 1587.360 414.375 1587.405 ;
        RECT 276.085 1587.220 299.835 1587.360 ;
        RECT 276.085 1587.175 276.375 1587.220 ;
        RECT 299.545 1587.175 299.835 1587.220 ;
        RECT 375.060 1587.220 414.375 1587.360 ;
        RECT 372.685 1587.020 372.975 1587.065 ;
        RECT 375.060 1587.020 375.200 1587.220 ;
        RECT 414.085 1587.175 414.375 1587.220 ;
        RECT 423.745 1587.360 424.035 1587.405 ;
        RECT 481.705 1587.360 481.995 1587.405 ;
        RECT 423.745 1587.220 444.660 1587.360 ;
        RECT 423.745 1587.175 424.035 1587.220 ;
        RECT 372.685 1586.880 375.200 1587.020 ;
        RECT 444.520 1587.020 444.660 1587.220 ;
        RECT 472.120 1587.220 481.995 1587.360 ;
        RECT 472.120 1587.020 472.260 1587.220 ;
        RECT 481.705 1587.175 481.995 1587.220 ;
        RECT 444.520 1586.880 472.260 1587.020 ;
        RECT 372.685 1586.835 372.975 1586.880 ;
        RECT 252.610 18.260 252.930 18.320 ;
        RECT 254.910 18.260 255.230 18.320 ;
        RECT 252.610 18.120 255.230 18.260 ;
        RECT 252.610 18.060 252.930 18.120 ;
        RECT 254.910 18.060 255.230 18.120 ;
      LAYER via ;
        RECT 505.640 1592.940 505.900 1593.200 ;
        RECT 254.940 1589.540 255.200 1589.800 ;
        RECT 252.640 18.060 252.900 18.320 ;
        RECT 254.940 18.060 255.200 18.320 ;
      LAYER met2 ;
        RECT 505.640 1600.000 505.920 1604.000 ;
        RECT 505.700 1593.230 505.840 1600.000 ;
        RECT 505.640 1592.910 505.900 1593.230 ;
        RECT 254.940 1589.510 255.200 1589.830 ;
        RECT 255.000 18.350 255.140 1589.510 ;
        RECT 252.640 18.030 252.900 18.350 ;
        RECT 254.940 18.030 255.200 18.350 ;
        RECT 252.700 2.400 252.840 18.030 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 513.890 1587.360 514.210 1587.420 ;
        RECT 519.870 1587.360 520.190 1587.420 ;
        RECT 513.890 1587.220 520.190 1587.360 ;
        RECT 513.890 1587.160 514.210 1587.220 ;
        RECT 519.870 1587.160 520.190 1587.220 ;
        RECT 270.090 18.260 270.410 18.320 ;
        RECT 513.890 18.260 514.210 18.320 ;
        RECT 270.090 18.120 514.210 18.260 ;
        RECT 270.090 18.060 270.410 18.120 ;
        RECT 513.890 18.060 514.210 18.120 ;
      LAYER via ;
        RECT 513.920 1587.160 514.180 1587.420 ;
        RECT 519.900 1587.160 520.160 1587.420 ;
        RECT 270.120 18.060 270.380 18.320 ;
        RECT 513.920 18.060 514.180 18.320 ;
      LAYER met2 ;
        RECT 519.900 1600.000 520.180 1604.000 ;
        RECT 519.960 1587.450 520.100 1600.000 ;
        RECT 513.920 1587.130 514.180 1587.450 ;
        RECT 519.900 1587.130 520.160 1587.450 ;
        RECT 513.980 18.350 514.120 1587.130 ;
        RECT 270.120 18.030 270.380 18.350 ;
        RECT 513.920 18.030 514.180 18.350 ;
        RECT 270.180 2.400 270.320 18.030 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 1588.720 289.730 1588.780 ;
        RECT 534.590 1588.720 534.910 1588.780 ;
        RECT 289.410 1588.580 463.060 1588.720 ;
        RECT 289.410 1588.520 289.730 1588.580 ;
        RECT 462.920 1588.380 463.060 1588.580 ;
        RECT 472.120 1588.580 534.910 1588.720 ;
        RECT 472.120 1588.380 472.260 1588.580 ;
        RECT 534.590 1588.520 534.910 1588.580 ;
        RECT 462.920 1588.240 472.260 1588.380 ;
      LAYER via ;
        RECT 289.440 1588.520 289.700 1588.780 ;
        RECT 534.620 1588.520 534.880 1588.780 ;
      LAYER met2 ;
        RECT 534.620 1600.000 534.900 1604.000 ;
        RECT 534.680 1588.810 534.820 1600.000 ;
        RECT 289.440 1588.490 289.700 1588.810 ;
        RECT 534.620 1588.490 534.880 1588.810 ;
        RECT 289.500 3.130 289.640 1588.490 ;
        RECT 288.120 2.990 289.640 3.130 ;
        RECT 288.120 2.400 288.260 2.990 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 20.640 306.290 20.700 ;
        RECT 310.110 20.640 310.430 20.700 ;
        RECT 305.970 20.500 310.430 20.640 ;
        RECT 305.970 20.440 306.290 20.500 ;
        RECT 310.110 20.440 310.430 20.500 ;
      LAYER via ;
        RECT 306.000 20.440 306.260 20.700 ;
        RECT 310.140 20.440 310.400 20.700 ;
      LAYER met2 ;
        RECT 549.340 1600.450 549.620 1604.000 ;
        RECT 547.560 1600.310 549.620 1600.450 ;
        RECT 547.560 1590.365 547.700 1600.310 ;
        RECT 549.340 1600.000 549.620 1600.310 ;
        RECT 310.130 1589.995 310.410 1590.365 ;
        RECT 547.490 1589.995 547.770 1590.365 ;
        RECT 310.200 20.730 310.340 1589.995 ;
        RECT 306.000 20.410 306.260 20.730 ;
        RECT 310.140 20.410 310.400 20.730 ;
        RECT 306.060 2.400 306.200 20.410 ;
        RECT 305.850 -4.800 306.410 2.400 ;
      LAYER via2 ;
        RECT 310.130 1590.040 310.410 1590.320 ;
        RECT 547.490 1590.040 547.770 1590.320 ;
      LAYER met3 ;
        RECT 310.105 1590.330 310.435 1590.345 ;
        RECT 547.465 1590.330 547.795 1590.345 ;
        RECT 310.105 1590.030 547.795 1590.330 ;
        RECT 310.105 1590.015 310.435 1590.030 ;
        RECT 547.465 1590.015 547.795 1590.030 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 17.580 324.230 17.640 ;
        RECT 548.390 17.580 548.710 17.640 ;
        RECT 323.910 17.440 548.710 17.580 ;
        RECT 323.910 17.380 324.230 17.440 ;
        RECT 548.390 17.380 548.710 17.440 ;
      LAYER via ;
        RECT 323.940 17.380 324.200 17.640 ;
        RECT 548.420 17.380 548.680 17.640 ;
      LAYER met2 ;
        RECT 563.600 1600.000 563.880 1604.000 ;
        RECT 563.660 1590.365 563.800 1600.000 ;
        RECT 548.410 1589.995 548.690 1590.365 ;
        RECT 563.590 1589.995 563.870 1590.365 ;
        RECT 548.480 17.670 548.620 1589.995 ;
        RECT 323.940 17.350 324.200 17.670 ;
        RECT 548.420 17.350 548.680 17.670 ;
        RECT 324.000 2.400 324.140 17.350 ;
        RECT 323.790 -4.800 324.350 2.400 ;
      LAYER via2 ;
        RECT 548.410 1590.040 548.690 1590.320 ;
        RECT 563.590 1590.040 563.870 1590.320 ;
      LAYER met3 ;
        RECT 548.385 1590.330 548.715 1590.345 ;
        RECT 563.565 1590.330 563.895 1590.345 ;
        RECT 548.385 1590.030 563.895 1590.330 ;
        RECT 548.385 1590.015 548.715 1590.030 ;
        RECT 563.565 1590.015 563.895 1590.030 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 344.610 1588.040 344.930 1588.100 ;
        RECT 578.290 1588.040 578.610 1588.100 ;
        RECT 344.610 1587.900 578.610 1588.040 ;
        RECT 344.610 1587.840 344.930 1587.900 ;
        RECT 578.290 1587.840 578.610 1587.900 ;
        RECT 341.390 20.640 341.710 20.700 ;
        RECT 344.610 20.640 344.930 20.700 ;
        RECT 341.390 20.500 344.930 20.640 ;
        RECT 341.390 20.440 341.710 20.500 ;
        RECT 344.610 20.440 344.930 20.500 ;
      LAYER via ;
        RECT 344.640 1587.840 344.900 1588.100 ;
        RECT 578.320 1587.840 578.580 1588.100 ;
        RECT 341.420 20.440 341.680 20.700 ;
        RECT 344.640 20.440 344.900 20.700 ;
      LAYER met2 ;
        RECT 578.320 1600.000 578.600 1604.000 ;
        RECT 578.380 1588.130 578.520 1600.000 ;
        RECT 344.640 1587.810 344.900 1588.130 ;
        RECT 578.320 1587.810 578.580 1588.130 ;
        RECT 344.700 20.730 344.840 1587.810 ;
        RECT 341.420 20.410 341.680 20.730 ;
        RECT 344.640 20.410 344.900 20.730 ;
        RECT 341.480 2.400 341.620 20.410 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 562.190 1591.100 562.510 1591.160 ;
        RECT 592.550 1591.100 592.870 1591.160 ;
        RECT 562.190 1590.960 592.870 1591.100 ;
        RECT 562.190 1590.900 562.510 1590.960 ;
        RECT 592.550 1590.900 592.870 1590.960 ;
        RECT 359.330 16.900 359.650 16.960 ;
        RECT 562.190 16.900 562.510 16.960 ;
        RECT 359.330 16.760 562.510 16.900 ;
        RECT 359.330 16.700 359.650 16.760 ;
        RECT 562.190 16.700 562.510 16.760 ;
      LAYER via ;
        RECT 562.220 1590.900 562.480 1591.160 ;
        RECT 592.580 1590.900 592.840 1591.160 ;
        RECT 359.360 16.700 359.620 16.960 ;
        RECT 562.220 16.700 562.480 16.960 ;
      LAYER met2 ;
        RECT 592.580 1600.000 592.860 1604.000 ;
        RECT 592.640 1591.190 592.780 1600.000 ;
        RECT 562.220 1590.870 562.480 1591.190 ;
        RECT 592.580 1590.870 592.840 1591.190 ;
        RECT 562.280 16.990 562.420 1590.870 ;
        RECT 359.360 16.670 359.620 16.990 ;
        RECT 562.220 16.670 562.480 16.990 ;
        RECT 359.420 2.400 359.560 16.670 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 379.110 1591.440 379.430 1591.500 ;
        RECT 607.270 1591.440 607.590 1591.500 ;
        RECT 379.110 1591.300 607.590 1591.440 ;
        RECT 379.110 1591.240 379.430 1591.300 ;
        RECT 607.270 1591.240 607.590 1591.300 ;
      LAYER via ;
        RECT 379.140 1591.240 379.400 1591.500 ;
        RECT 607.300 1591.240 607.560 1591.500 ;
      LAYER met2 ;
        RECT 607.300 1600.000 607.580 1604.000 ;
        RECT 607.360 1591.530 607.500 1600.000 ;
        RECT 379.140 1591.210 379.400 1591.530 ;
        RECT 607.300 1591.210 607.560 1591.530 ;
        RECT 379.200 3.130 379.340 1591.210 ;
        RECT 377.360 2.990 379.340 3.130 ;
        RECT 377.360 2.400 377.500 2.990 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 574.225 18.785 574.395 19.975 ;
      LAYER mcon ;
        RECT 574.225 19.805 574.395 19.975 ;
      LAYER met1 ;
        RECT 582.890 1588.040 583.210 1588.100 ;
        RECT 621.990 1588.040 622.310 1588.100 ;
        RECT 582.890 1587.900 622.310 1588.040 ;
        RECT 582.890 1587.840 583.210 1587.900 ;
        RECT 621.990 1587.840 622.310 1587.900 ;
        RECT 574.165 19.960 574.455 20.005 ;
        RECT 582.890 19.960 583.210 20.020 ;
        RECT 574.165 19.820 583.210 19.960 ;
        RECT 574.165 19.775 574.455 19.820 ;
        RECT 582.890 19.760 583.210 19.820 ;
        RECT 395.210 18.940 395.530 19.000 ;
        RECT 574.165 18.940 574.455 18.985 ;
        RECT 395.210 18.800 574.455 18.940 ;
        RECT 395.210 18.740 395.530 18.800 ;
        RECT 574.165 18.755 574.455 18.800 ;
      LAYER via ;
        RECT 582.920 1587.840 583.180 1588.100 ;
        RECT 622.020 1587.840 622.280 1588.100 ;
        RECT 582.920 19.760 583.180 20.020 ;
        RECT 395.240 18.740 395.500 19.000 ;
      LAYER met2 ;
        RECT 622.020 1600.000 622.300 1604.000 ;
        RECT 622.080 1588.130 622.220 1600.000 ;
        RECT 582.920 1587.810 583.180 1588.130 ;
        RECT 622.020 1587.810 622.280 1588.130 ;
        RECT 582.980 20.050 583.120 1587.810 ;
        RECT 582.920 19.730 583.180 20.050 ;
        RECT 395.240 18.710 395.500 19.030 ;
        RECT 395.300 2.400 395.440 18.710 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.150 1592.120 413.470 1592.180 ;
        RECT 636.250 1592.120 636.570 1592.180 ;
        RECT 413.150 1591.980 636.570 1592.120 ;
        RECT 413.150 1591.920 413.470 1591.980 ;
        RECT 636.250 1591.920 636.570 1591.980 ;
      LAYER via ;
        RECT 413.180 1591.920 413.440 1592.180 ;
        RECT 636.280 1591.920 636.540 1592.180 ;
      LAYER met2 ;
        RECT 636.280 1600.000 636.560 1604.000 ;
        RECT 636.340 1592.210 636.480 1600.000 ;
        RECT 413.180 1591.890 413.440 1592.210 ;
        RECT 636.280 1591.890 636.540 1592.210 ;
        RECT 413.240 1586.170 413.380 1591.890 ;
        RECT 413.240 1586.030 413.840 1586.170 ;
        RECT 413.700 3.130 413.840 1586.030 ;
        RECT 413.240 2.990 413.840 3.130 ;
        RECT 413.240 2.400 413.380 2.990 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 75.510 1591.440 75.830 1591.500 ;
        RECT 360.250 1591.440 360.570 1591.500 ;
        RECT 75.510 1591.300 360.570 1591.440 ;
        RECT 75.510 1591.240 75.830 1591.300 ;
        RECT 360.250 1591.240 360.570 1591.300 ;
        RECT 74.130 14.180 74.450 14.240 ;
        RECT 75.510 14.180 75.830 14.240 ;
        RECT 74.130 14.040 75.830 14.180 ;
        RECT 74.130 13.980 74.450 14.040 ;
        RECT 75.510 13.980 75.830 14.040 ;
      LAYER via ;
        RECT 75.540 1591.240 75.800 1591.500 ;
        RECT 360.280 1591.240 360.540 1591.500 ;
        RECT 74.160 13.980 74.420 14.240 ;
        RECT 75.540 13.980 75.800 14.240 ;
      LAYER met2 ;
        RECT 360.280 1600.000 360.560 1604.000 ;
        RECT 360.340 1591.530 360.480 1600.000 ;
        RECT 75.540 1591.210 75.800 1591.530 ;
        RECT 360.280 1591.210 360.540 1591.530 ;
        RECT 75.600 14.270 75.740 1591.210 ;
        RECT 74.160 13.950 74.420 14.270 ;
        RECT 75.540 13.950 75.800 14.270 ;
        RECT 74.220 2.400 74.360 13.950 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 573.765 19.805 573.935 20.655 ;
      LAYER mcon ;
        RECT 573.765 20.485 573.935 20.655 ;
      LAYER met1 ;
        RECT 573.705 20.640 573.995 20.685 ;
        RECT 573.705 20.500 601.980 20.640 ;
        RECT 573.705 20.455 573.995 20.500 ;
        RECT 601.840 20.300 601.980 20.500 ;
        RECT 610.490 20.300 610.810 20.360 ;
        RECT 601.840 20.160 610.810 20.300 ;
        RECT 610.490 20.100 610.810 20.160 ;
        RECT 573.705 19.960 573.995 20.005 ;
        RECT 445.440 19.820 573.995 19.960 ;
        RECT 432.010 19.620 432.330 19.680 ;
        RECT 445.440 19.620 445.580 19.820 ;
        RECT 573.705 19.775 573.995 19.820 ;
        RECT 432.010 19.480 445.580 19.620 ;
        RECT 432.010 19.420 432.330 19.480 ;
      LAYER via ;
        RECT 610.520 20.100 610.780 20.360 ;
        RECT 432.040 19.420 432.300 19.680 ;
      LAYER met2 ;
        RECT 651.000 1600.000 651.280 1604.000 ;
        RECT 651.060 1590.365 651.200 1600.000 ;
        RECT 610.510 1589.995 610.790 1590.365 ;
        RECT 650.990 1589.995 651.270 1590.365 ;
        RECT 610.580 20.390 610.720 1589.995 ;
        RECT 610.520 20.070 610.780 20.390 ;
        RECT 432.040 19.390 432.300 19.710 ;
        RECT 432.100 9.930 432.240 19.390 ;
        RECT 430.720 9.790 432.240 9.930 ;
        RECT 430.720 2.400 430.860 9.790 ;
        RECT 430.510 -4.800 431.070 2.400 ;
      LAYER via2 ;
        RECT 610.510 1590.040 610.790 1590.320 ;
        RECT 650.990 1590.040 651.270 1590.320 ;
      LAYER met3 ;
        RECT 610.485 1590.330 610.815 1590.345 ;
        RECT 650.965 1590.330 651.295 1590.345 ;
        RECT 610.485 1590.030 651.295 1590.330 ;
        RECT 610.485 1590.015 610.815 1590.030 ;
        RECT 650.965 1590.015 651.295 1590.030 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 454.550 1592.460 454.870 1592.520 ;
        RECT 665.230 1592.460 665.550 1592.520 ;
        RECT 454.550 1592.320 665.550 1592.460 ;
        RECT 454.550 1592.260 454.870 1592.320 ;
        RECT 665.230 1592.260 665.550 1592.320 ;
        RECT 448.570 20.640 448.890 20.700 ;
        RECT 454.550 20.640 454.870 20.700 ;
        RECT 448.570 20.500 454.870 20.640 ;
        RECT 448.570 20.440 448.890 20.500 ;
        RECT 454.550 20.440 454.870 20.500 ;
      LAYER via ;
        RECT 454.580 1592.260 454.840 1592.520 ;
        RECT 665.260 1592.260 665.520 1592.520 ;
        RECT 448.600 20.440 448.860 20.700 ;
        RECT 454.580 20.440 454.840 20.700 ;
      LAYER met2 ;
        RECT 665.260 1600.000 665.540 1604.000 ;
        RECT 665.320 1592.550 665.460 1600.000 ;
        RECT 454.580 1592.230 454.840 1592.550 ;
        RECT 665.260 1592.230 665.520 1592.550 ;
        RECT 454.640 20.730 454.780 1592.230 ;
        RECT 448.600 20.410 448.860 20.730 ;
        RECT 454.580 20.410 454.840 20.730 ;
        RECT 448.660 2.400 448.800 20.410 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 1592.800 469.130 1592.860 ;
        RECT 679.950 1592.800 680.270 1592.860 ;
        RECT 468.810 1592.660 680.270 1592.800 ;
        RECT 468.810 1592.600 469.130 1592.660 ;
        RECT 679.950 1592.600 680.270 1592.660 ;
        RECT 466.510 20.640 466.830 20.700 ;
        RECT 468.810 20.640 469.130 20.700 ;
        RECT 466.510 20.500 469.130 20.640 ;
        RECT 466.510 20.440 466.830 20.500 ;
        RECT 468.810 20.440 469.130 20.500 ;
      LAYER via ;
        RECT 468.840 1592.600 469.100 1592.860 ;
        RECT 679.980 1592.600 680.240 1592.860 ;
        RECT 466.540 20.440 466.800 20.700 ;
        RECT 468.840 20.440 469.100 20.700 ;
      LAYER met2 ;
        RECT 679.980 1600.000 680.260 1604.000 ;
        RECT 680.040 1592.890 680.180 1600.000 ;
        RECT 468.840 1592.570 469.100 1592.890 ;
        RECT 679.980 1592.570 680.240 1592.890 ;
        RECT 468.900 20.730 469.040 1592.570 ;
        RECT 466.540 20.410 466.800 20.730 ;
        RECT 468.840 20.410 469.100 20.730 ;
        RECT 466.600 2.400 466.740 20.410 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 578.365 18.785 578.535 20.315 ;
      LAYER mcon ;
        RECT 578.365 20.145 578.535 20.315 ;
      LAYER met1 ;
        RECT 624.290 1587.700 624.610 1587.760 ;
        RECT 694.670 1587.700 694.990 1587.760 ;
        RECT 624.290 1587.560 694.990 1587.700 ;
        RECT 624.290 1587.500 624.610 1587.560 ;
        RECT 694.670 1587.500 694.990 1587.560 ;
        RECT 484.450 20.300 484.770 20.360 ;
        RECT 578.305 20.300 578.595 20.345 ;
        RECT 484.450 20.160 578.595 20.300 ;
        RECT 484.450 20.100 484.770 20.160 ;
        RECT 578.305 20.115 578.595 20.160 ;
        RECT 578.305 18.940 578.595 18.985 ;
        RECT 624.290 18.940 624.610 19.000 ;
        RECT 578.305 18.800 624.610 18.940 ;
        RECT 578.305 18.755 578.595 18.800 ;
        RECT 624.290 18.740 624.610 18.800 ;
      LAYER via ;
        RECT 624.320 1587.500 624.580 1587.760 ;
        RECT 694.700 1587.500 694.960 1587.760 ;
        RECT 484.480 20.100 484.740 20.360 ;
        RECT 624.320 18.740 624.580 19.000 ;
      LAYER met2 ;
        RECT 694.700 1600.000 694.980 1604.000 ;
        RECT 694.760 1587.790 694.900 1600.000 ;
        RECT 624.320 1587.470 624.580 1587.790 ;
        RECT 694.700 1587.470 694.960 1587.790 ;
        RECT 484.480 20.070 484.740 20.390 ;
        RECT 484.540 2.400 484.680 20.070 ;
        RECT 624.380 19.030 624.520 1587.470 ;
        RECT 624.320 18.710 624.580 19.030 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 1593.480 503.630 1593.540 ;
        RECT 708.930 1593.480 709.250 1593.540 ;
        RECT 503.310 1593.340 506.760 1593.480 ;
        RECT 503.310 1593.280 503.630 1593.340 ;
        RECT 506.620 1593.140 506.760 1593.340 ;
        RECT 543.880 1593.340 709.250 1593.480 ;
        RECT 543.880 1593.140 544.020 1593.340 ;
        RECT 708.930 1593.280 709.250 1593.340 ;
        RECT 506.620 1593.000 544.020 1593.140 ;
      LAYER via ;
        RECT 503.340 1593.280 503.600 1593.540 ;
        RECT 708.960 1593.280 709.220 1593.540 ;
      LAYER met2 ;
        RECT 708.960 1600.000 709.240 1604.000 ;
        RECT 709.020 1593.570 709.160 1600.000 ;
        RECT 503.340 1593.250 503.600 1593.570 ;
        RECT 708.960 1593.250 709.220 1593.570 ;
        RECT 503.400 3.130 503.540 1593.250 ;
        RECT 502.480 2.990 503.540 3.130 ;
        RECT 502.480 2.400 502.620 2.990 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 638.550 1588.040 638.870 1588.100 ;
        RECT 723.650 1588.040 723.970 1588.100 ;
        RECT 638.550 1587.900 723.970 1588.040 ;
        RECT 638.550 1587.840 638.870 1587.900 ;
        RECT 723.650 1587.840 723.970 1587.900 ;
        RECT 519.870 15.540 520.190 15.600 ;
        RECT 638.550 15.540 638.870 15.600 ;
        RECT 519.870 15.400 638.870 15.540 ;
        RECT 519.870 15.340 520.190 15.400 ;
        RECT 638.550 15.340 638.870 15.400 ;
      LAYER via ;
        RECT 638.580 1587.840 638.840 1588.100 ;
        RECT 723.680 1587.840 723.940 1588.100 ;
        RECT 519.900 15.340 520.160 15.600 ;
        RECT 638.580 15.340 638.840 15.600 ;
      LAYER met2 ;
        RECT 723.680 1600.000 723.960 1604.000 ;
        RECT 723.740 1588.130 723.880 1600.000 ;
        RECT 638.580 1587.810 638.840 1588.130 ;
        RECT 723.680 1587.810 723.940 1588.130 ;
        RECT 638.640 15.630 638.780 1587.810 ;
        RECT 519.900 15.310 520.160 15.630 ;
        RECT 638.580 15.310 638.840 15.630 ;
        RECT 519.960 2.400 520.100 15.310 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 575.605 1588.565 575.775 1593.835 ;
      LAYER mcon ;
        RECT 575.605 1593.665 575.775 1593.835 ;
      LAYER met1 ;
        RECT 575.545 1593.820 575.835 1593.865 ;
        RECT 737.910 1593.820 738.230 1593.880 ;
        RECT 575.545 1593.680 738.230 1593.820 ;
        RECT 575.545 1593.635 575.835 1593.680 ;
        RECT 737.910 1593.620 738.230 1593.680 ;
        RECT 537.810 1588.720 538.130 1588.780 ;
        RECT 575.545 1588.720 575.835 1588.765 ;
        RECT 537.810 1588.580 575.835 1588.720 ;
        RECT 537.810 1588.520 538.130 1588.580 ;
        RECT 575.545 1588.535 575.835 1588.580 ;
      LAYER via ;
        RECT 737.940 1593.620 738.200 1593.880 ;
        RECT 537.840 1588.520 538.100 1588.780 ;
      LAYER met2 ;
        RECT 737.940 1600.000 738.220 1604.000 ;
        RECT 738.000 1593.910 738.140 1600.000 ;
        RECT 737.940 1593.590 738.200 1593.910 ;
        RECT 537.840 1588.490 538.100 1588.810 ;
        RECT 537.900 2.400 538.040 1588.490 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 638.090 1592.120 638.410 1592.180 ;
        RECT 752.630 1592.120 752.950 1592.180 ;
        RECT 638.090 1591.980 752.950 1592.120 ;
        RECT 638.090 1591.920 638.410 1591.980 ;
        RECT 752.630 1591.920 752.950 1591.980 ;
        RECT 555.750 14.860 556.070 14.920 ;
        RECT 638.090 14.860 638.410 14.920 ;
        RECT 555.750 14.720 638.410 14.860 ;
        RECT 555.750 14.660 556.070 14.720 ;
        RECT 638.090 14.660 638.410 14.720 ;
      LAYER via ;
        RECT 638.120 1591.920 638.380 1592.180 ;
        RECT 752.660 1591.920 752.920 1592.180 ;
        RECT 555.780 14.660 556.040 14.920 ;
        RECT 638.120 14.660 638.380 14.920 ;
      LAYER met2 ;
        RECT 752.660 1600.000 752.940 1604.000 ;
        RECT 752.720 1592.210 752.860 1600.000 ;
        RECT 638.120 1591.890 638.380 1592.210 ;
        RECT 752.660 1591.890 752.920 1592.210 ;
        RECT 638.180 14.950 638.320 1591.890 ;
        RECT 555.780 14.630 556.040 14.950 ;
        RECT 638.120 14.630 638.380 14.950 ;
        RECT 555.840 2.400 555.980 14.630 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 720.890 1592.460 721.210 1592.520 ;
        RECT 767.350 1592.460 767.670 1592.520 ;
        RECT 720.890 1592.320 767.670 1592.460 ;
        RECT 720.890 1592.260 721.210 1592.320 ;
        RECT 767.350 1592.260 767.670 1592.320 ;
        RECT 573.690 15.880 574.010 15.940 ;
        RECT 720.890 15.880 721.210 15.940 ;
        RECT 573.690 15.740 721.210 15.880 ;
        RECT 573.690 15.680 574.010 15.740 ;
        RECT 720.890 15.680 721.210 15.740 ;
      LAYER via ;
        RECT 720.920 1592.260 721.180 1592.520 ;
        RECT 767.380 1592.260 767.640 1592.520 ;
        RECT 573.720 15.680 573.980 15.940 ;
        RECT 720.920 15.680 721.180 15.940 ;
      LAYER met2 ;
        RECT 767.380 1600.000 767.660 1604.000 ;
        RECT 767.440 1592.550 767.580 1600.000 ;
        RECT 720.920 1592.230 721.180 1592.550 ;
        RECT 767.380 1592.230 767.640 1592.550 ;
        RECT 720.980 15.970 721.120 1592.230 ;
        RECT 573.720 15.650 573.980 15.970 ;
        RECT 720.920 15.650 721.180 15.970 ;
        RECT 573.780 2.400 573.920 15.650 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 621.605 15.045 621.775 16.575 ;
        RECT 675.885 14.705 676.055 16.915 ;
      LAYER mcon ;
        RECT 675.885 16.745 676.055 16.915 ;
        RECT 621.605 16.405 621.775 16.575 ;
      LAYER met1 ;
        RECT 755.390 1587.360 755.710 1587.420 ;
        RECT 781.610 1587.360 781.930 1587.420 ;
        RECT 755.390 1587.220 781.930 1587.360 ;
        RECT 755.390 1587.160 755.710 1587.220 ;
        RECT 781.610 1587.160 781.930 1587.220 ;
        RECT 675.825 16.900 676.115 16.945 ;
        RECT 676.730 16.900 677.050 16.960 ;
        RECT 675.825 16.760 677.050 16.900 ;
        RECT 675.825 16.715 676.115 16.760 ;
        RECT 676.730 16.700 677.050 16.760 ;
        RECT 677.650 16.900 677.970 16.960 ;
        RECT 755.390 16.900 755.710 16.960 ;
        RECT 677.650 16.760 755.710 16.900 ;
        RECT 677.650 16.700 677.970 16.760 ;
        RECT 755.390 16.700 755.710 16.760 ;
        RECT 591.170 16.560 591.490 16.620 ;
        RECT 621.545 16.560 621.835 16.605 ;
        RECT 591.170 16.420 621.835 16.560 ;
        RECT 591.170 16.360 591.490 16.420 ;
        RECT 621.545 16.375 621.835 16.420 ;
        RECT 621.545 15.200 621.835 15.245 ;
        RECT 621.545 15.060 638.780 15.200 ;
        RECT 621.545 15.015 621.835 15.060 ;
        RECT 638.640 14.860 638.780 15.060 ;
        RECT 675.825 14.860 676.115 14.905 ;
        RECT 638.640 14.720 676.115 14.860 ;
        RECT 675.825 14.675 676.115 14.720 ;
      LAYER via ;
        RECT 755.420 1587.160 755.680 1587.420 ;
        RECT 781.640 1587.160 781.900 1587.420 ;
        RECT 676.760 16.700 677.020 16.960 ;
        RECT 677.680 16.700 677.940 16.960 ;
        RECT 755.420 16.700 755.680 16.960 ;
        RECT 591.200 16.360 591.460 16.620 ;
      LAYER met2 ;
        RECT 781.640 1600.000 781.920 1604.000 ;
        RECT 781.700 1587.450 781.840 1600.000 ;
        RECT 755.420 1587.130 755.680 1587.450 ;
        RECT 781.640 1587.130 781.900 1587.450 ;
        RECT 755.480 16.990 755.620 1587.130 ;
        RECT 676.760 16.730 677.020 16.990 ;
        RECT 677.680 16.730 677.940 16.990 ;
        RECT 676.760 16.670 677.940 16.730 ;
        RECT 755.420 16.670 755.680 16.990 ;
        RECT 591.200 16.330 591.460 16.650 ;
        RECT 676.820 16.590 677.880 16.670 ;
        RECT 591.260 2.400 591.400 16.330 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 226.925 15.045 227.095 16.915 ;
        RECT 278.905 14.365 279.075 16.915 ;
      LAYER mcon ;
        RECT 226.925 16.745 227.095 16.915 ;
        RECT 278.905 16.745 279.075 16.915 ;
      LAYER met1 ;
        RECT 334.490 1587.700 334.810 1587.760 ;
        RECT 379.570 1587.700 379.890 1587.760 ;
        RECT 334.490 1587.560 379.890 1587.700 ;
        RECT 334.490 1587.500 334.810 1587.560 ;
        RECT 379.570 1587.500 379.890 1587.560 ;
        RECT 97.590 16.900 97.910 16.960 ;
        RECT 179.470 16.900 179.790 16.960 ;
        RECT 97.590 16.760 179.790 16.900 ;
        RECT 97.590 16.700 97.910 16.760 ;
        RECT 179.470 16.700 179.790 16.760 ;
        RECT 226.865 16.900 227.155 16.945 ;
        RECT 278.845 16.900 279.135 16.945 ;
        RECT 226.865 16.760 279.135 16.900 ;
        RECT 226.865 16.715 227.155 16.760 ;
        RECT 278.845 16.715 279.135 16.760 ;
        RECT 179.470 15.200 179.790 15.260 ;
        RECT 226.865 15.200 227.155 15.245 ;
        RECT 179.470 15.060 227.155 15.200 ;
        RECT 179.470 15.000 179.790 15.060 ;
        RECT 226.865 15.015 227.155 15.060 ;
        RECT 278.845 14.520 279.135 14.565 ;
        RECT 334.490 14.520 334.810 14.580 ;
        RECT 278.845 14.380 334.810 14.520 ;
        RECT 278.845 14.335 279.135 14.380 ;
        RECT 334.490 14.320 334.810 14.380 ;
      LAYER via ;
        RECT 334.520 1587.500 334.780 1587.760 ;
        RECT 379.600 1587.500 379.860 1587.760 ;
        RECT 97.620 16.700 97.880 16.960 ;
        RECT 179.500 16.700 179.760 16.960 ;
        RECT 179.500 15.000 179.760 15.260 ;
        RECT 334.520 14.320 334.780 14.580 ;
      LAYER met2 ;
        RECT 379.600 1600.000 379.880 1604.000 ;
        RECT 379.660 1587.790 379.800 1600.000 ;
        RECT 334.520 1587.470 334.780 1587.790 ;
        RECT 379.600 1587.470 379.860 1587.790 ;
        RECT 97.620 16.670 97.880 16.990 ;
        RECT 179.500 16.670 179.760 16.990 ;
        RECT 97.680 2.400 97.820 16.670 ;
        RECT 179.560 15.290 179.700 16.670 ;
        RECT 179.500 14.970 179.760 15.290 ;
        RECT 334.580 14.610 334.720 1587.470 ;
        RECT 334.520 14.290 334.780 14.610 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 613.710 1590.760 614.030 1590.820 ;
        RECT 796.330 1590.760 796.650 1590.820 ;
        RECT 613.710 1590.620 796.650 1590.760 ;
        RECT 613.710 1590.560 614.030 1590.620 ;
        RECT 796.330 1590.560 796.650 1590.620 ;
        RECT 609.110 20.640 609.430 20.700 ;
        RECT 613.710 20.640 614.030 20.700 ;
        RECT 609.110 20.500 614.030 20.640 ;
        RECT 609.110 20.440 609.430 20.500 ;
        RECT 613.710 20.440 614.030 20.500 ;
      LAYER via ;
        RECT 613.740 1590.560 614.000 1590.820 ;
        RECT 796.360 1590.560 796.620 1590.820 ;
        RECT 609.140 20.440 609.400 20.700 ;
        RECT 613.740 20.440 614.000 20.700 ;
      LAYER met2 ;
        RECT 796.360 1600.000 796.640 1604.000 ;
        RECT 796.420 1590.850 796.560 1600.000 ;
        RECT 613.740 1590.530 614.000 1590.850 ;
        RECT 796.360 1590.530 796.620 1590.850 ;
        RECT 613.800 20.730 613.940 1590.530 ;
        RECT 609.140 20.410 609.400 20.730 ;
        RECT 613.740 20.410 614.000 20.730 ;
        RECT 609.200 2.400 609.340 20.410 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 676.345 16.405 677.435 16.575 ;
      LAYER mcon ;
        RECT 677.265 16.405 677.435 16.575 ;
      LAYER met1 ;
        RECT 789.890 1587.360 790.210 1587.420 ;
        RECT 810.590 1587.360 810.910 1587.420 ;
        RECT 789.890 1587.220 810.910 1587.360 ;
        RECT 789.890 1587.160 790.210 1587.220 ;
        RECT 810.590 1587.160 810.910 1587.220 ;
        RECT 627.050 16.560 627.370 16.620 ;
        RECT 676.285 16.560 676.575 16.605 ;
        RECT 627.050 16.420 676.575 16.560 ;
        RECT 627.050 16.360 627.370 16.420 ;
        RECT 676.285 16.375 676.575 16.420 ;
        RECT 677.205 16.560 677.495 16.605 ;
        RECT 789.890 16.560 790.210 16.620 ;
        RECT 677.205 16.420 790.210 16.560 ;
        RECT 677.205 16.375 677.495 16.420 ;
        RECT 789.890 16.360 790.210 16.420 ;
      LAYER via ;
        RECT 789.920 1587.160 790.180 1587.420 ;
        RECT 810.620 1587.160 810.880 1587.420 ;
        RECT 627.080 16.360 627.340 16.620 ;
        RECT 789.920 16.360 790.180 16.620 ;
      LAYER met2 ;
        RECT 810.620 1600.000 810.900 1604.000 ;
        RECT 810.680 1587.450 810.820 1600.000 ;
        RECT 789.920 1587.130 790.180 1587.450 ;
        RECT 810.620 1587.130 810.880 1587.450 ;
        RECT 789.980 16.650 790.120 1587.130 ;
        RECT 627.080 16.330 627.340 16.650 ;
        RECT 789.920 16.330 790.180 16.650 ;
        RECT 627.140 2.400 627.280 16.330 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 362.090 1589.060 362.410 1589.120 ;
        RECT 396.130 1589.060 396.450 1589.120 ;
        RECT 362.090 1588.920 396.450 1589.060 ;
        RECT 362.090 1588.860 362.410 1588.920 ;
        RECT 396.130 1588.860 396.450 1588.920 ;
        RECT 121.510 18.940 121.830 19.000 ;
        RECT 362.090 18.940 362.410 19.000 ;
        RECT 121.510 18.800 362.410 18.940 ;
        RECT 121.510 18.740 121.830 18.800 ;
        RECT 362.090 18.740 362.410 18.800 ;
      LAYER via ;
        RECT 362.120 1588.860 362.380 1589.120 ;
        RECT 396.160 1588.860 396.420 1589.120 ;
        RECT 121.540 18.740 121.800 19.000 ;
        RECT 362.120 18.740 362.380 19.000 ;
      LAYER met2 ;
        RECT 398.920 1600.450 399.200 1604.000 ;
        RECT 396.220 1600.310 399.200 1600.450 ;
        RECT 396.220 1589.150 396.360 1600.310 ;
        RECT 398.920 1600.000 399.200 1600.310 ;
        RECT 362.120 1588.830 362.380 1589.150 ;
        RECT 396.160 1588.830 396.420 1589.150 ;
        RECT 362.180 19.030 362.320 1588.830 ;
        RECT 121.540 18.710 121.800 19.030 ;
        RECT 362.120 18.710 362.380 19.030 ;
        RECT 121.600 2.400 121.740 18.710 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 395.285 1589.925 395.455 1593.495 ;
      LAYER mcon ;
        RECT 395.285 1593.325 395.455 1593.495 ;
      LAYER met1 ;
        RECT 395.225 1593.480 395.515 1593.525 ;
        RECT 416.830 1593.480 417.150 1593.540 ;
        RECT 395.225 1593.340 417.150 1593.480 ;
        RECT 395.225 1593.295 395.515 1593.340 ;
        RECT 416.830 1593.280 417.150 1593.340 ;
        RECT 161.990 1590.080 162.310 1590.140 ;
        RECT 395.225 1590.080 395.515 1590.125 ;
        RECT 161.990 1589.940 395.515 1590.080 ;
        RECT 161.990 1589.880 162.310 1589.940 ;
        RECT 395.225 1589.895 395.515 1589.940 ;
        RECT 145.430 17.920 145.750 17.980 ;
        RECT 161.990 17.920 162.310 17.980 ;
        RECT 145.430 17.780 162.310 17.920 ;
        RECT 145.430 17.720 145.750 17.780 ;
        RECT 161.990 17.720 162.310 17.780 ;
      LAYER via ;
        RECT 416.860 1593.280 417.120 1593.540 ;
        RECT 162.020 1589.880 162.280 1590.140 ;
        RECT 145.460 17.720 145.720 17.980 ;
        RECT 162.020 17.720 162.280 17.980 ;
      LAYER met2 ;
        RECT 418.240 1600.450 418.520 1604.000 ;
        RECT 416.920 1600.310 418.520 1600.450 ;
        RECT 416.920 1593.570 417.060 1600.310 ;
        RECT 418.240 1600.000 418.520 1600.310 ;
        RECT 416.860 1593.250 417.120 1593.570 ;
        RECT 162.020 1589.850 162.280 1590.170 ;
        RECT 162.080 18.010 162.220 1589.850 ;
        RECT 145.460 17.690 145.720 18.010 ;
        RECT 162.020 17.690 162.280 18.010 ;
        RECT 145.520 2.400 145.660 17.690 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 397.050 1589.060 397.370 1589.120 ;
        RECT 430.630 1589.060 430.950 1589.120 ;
        RECT 397.050 1588.920 430.950 1589.060 ;
        RECT 397.050 1588.860 397.370 1588.920 ;
        RECT 430.630 1588.860 430.950 1588.920 ;
        RECT 163.370 19.280 163.690 19.340 ;
        RECT 397.050 19.280 397.370 19.340 ;
        RECT 163.370 19.140 397.370 19.280 ;
        RECT 163.370 19.080 163.690 19.140 ;
        RECT 397.050 19.080 397.370 19.140 ;
      LAYER via ;
        RECT 397.080 1588.860 397.340 1589.120 ;
        RECT 430.660 1588.860 430.920 1589.120 ;
        RECT 163.400 19.080 163.660 19.340 ;
        RECT 397.080 19.080 397.340 19.340 ;
      LAYER met2 ;
        RECT 432.960 1600.450 433.240 1604.000 ;
        RECT 430.720 1600.310 433.240 1600.450 ;
        RECT 430.720 1589.150 430.860 1600.310 ;
        RECT 432.960 1600.000 433.240 1600.310 ;
        RECT 397.080 1588.830 397.340 1589.150 ;
        RECT 430.660 1588.830 430.920 1589.150 ;
        RECT 397.140 19.370 397.280 1588.830 ;
        RECT 163.400 19.050 163.660 19.370 ;
        RECT 397.080 19.050 397.340 19.370 ;
        RECT 163.460 2.400 163.600 19.050 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 424.190 1590.080 424.510 1590.140 ;
        RECT 447.190 1590.080 447.510 1590.140 ;
        RECT 424.190 1589.940 447.510 1590.080 ;
        RECT 424.190 1589.880 424.510 1589.940 ;
        RECT 447.190 1589.880 447.510 1589.940 ;
        RECT 180.850 18.600 181.170 18.660 ;
        RECT 424.190 18.600 424.510 18.660 ;
        RECT 180.850 18.460 424.510 18.600 ;
        RECT 180.850 18.400 181.170 18.460 ;
        RECT 424.190 18.400 424.510 18.460 ;
      LAYER via ;
        RECT 424.220 1589.880 424.480 1590.140 ;
        RECT 447.220 1589.880 447.480 1590.140 ;
        RECT 180.880 18.400 181.140 18.660 ;
        RECT 424.220 18.400 424.480 18.660 ;
      LAYER met2 ;
        RECT 447.220 1600.000 447.500 1604.000 ;
        RECT 447.280 1590.170 447.420 1600.000 ;
        RECT 424.220 1589.850 424.480 1590.170 ;
        RECT 447.220 1589.850 447.480 1590.170 ;
        RECT 424.280 18.690 424.420 1589.850 ;
        RECT 180.880 18.370 181.140 18.690 ;
        RECT 424.220 18.370 424.480 18.690 ;
        RECT 180.940 2.400 181.080 18.370 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 431.550 1589.060 431.870 1589.120 ;
        RECT 461.910 1589.060 462.230 1589.120 ;
        RECT 431.550 1588.920 462.230 1589.060 ;
        RECT 431.550 1588.860 431.870 1588.920 ;
        RECT 461.910 1588.860 462.230 1588.920 ;
        RECT 198.790 19.620 199.110 19.680 ;
        RECT 431.550 19.620 431.870 19.680 ;
        RECT 198.790 19.480 431.870 19.620 ;
        RECT 198.790 19.420 199.110 19.480 ;
        RECT 431.550 19.420 431.870 19.480 ;
      LAYER via ;
        RECT 431.580 1588.860 431.840 1589.120 ;
        RECT 461.940 1588.860 462.200 1589.120 ;
        RECT 198.820 19.420 199.080 19.680 ;
        RECT 431.580 19.420 431.840 19.680 ;
      LAYER met2 ;
        RECT 461.940 1600.000 462.220 1604.000 ;
        RECT 462.000 1589.150 462.140 1600.000 ;
        RECT 431.580 1588.830 431.840 1589.150 ;
        RECT 461.940 1588.830 462.200 1589.150 ;
        RECT 431.640 19.710 431.780 1588.830 ;
        RECT 198.820 19.390 199.080 19.710 ;
        RECT 431.580 19.390 431.840 19.710 ;
        RECT 198.880 2.400 199.020 19.390 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 220.410 1593.140 220.730 1593.200 ;
        RECT 476.630 1593.140 476.950 1593.200 ;
        RECT 220.410 1593.000 476.950 1593.140 ;
        RECT 220.410 1592.940 220.730 1593.000 ;
        RECT 476.630 1592.940 476.950 1593.000 ;
        RECT 216.730 18.260 217.050 18.320 ;
        RECT 220.410 18.260 220.730 18.320 ;
        RECT 216.730 18.120 220.730 18.260 ;
        RECT 216.730 18.060 217.050 18.120 ;
        RECT 220.410 18.060 220.730 18.120 ;
      LAYER via ;
        RECT 220.440 1592.940 220.700 1593.200 ;
        RECT 476.660 1592.940 476.920 1593.200 ;
        RECT 216.760 18.060 217.020 18.320 ;
        RECT 220.440 18.060 220.700 18.320 ;
      LAYER met2 ;
        RECT 476.660 1600.000 476.940 1604.000 ;
        RECT 476.720 1593.230 476.860 1600.000 ;
        RECT 220.440 1592.910 220.700 1593.230 ;
        RECT 476.660 1592.910 476.920 1593.230 ;
        RECT 220.500 18.350 220.640 1592.910 ;
        RECT 216.760 18.030 217.020 18.350 ;
        RECT 220.440 18.030 220.700 18.350 ;
        RECT 216.820 2.400 216.960 18.030 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 459.150 1587.700 459.470 1587.760 ;
        RECT 490.890 1587.700 491.210 1587.760 ;
        RECT 459.150 1587.560 491.210 1587.700 ;
        RECT 459.150 1587.500 459.470 1587.560 ;
        RECT 490.890 1587.500 491.210 1587.560 ;
        RECT 234.670 16.220 234.990 16.280 ;
        RECT 459.150 16.220 459.470 16.280 ;
        RECT 234.670 16.080 459.470 16.220 ;
        RECT 234.670 16.020 234.990 16.080 ;
        RECT 459.150 16.020 459.470 16.080 ;
      LAYER via ;
        RECT 459.180 1587.500 459.440 1587.760 ;
        RECT 490.920 1587.500 491.180 1587.760 ;
        RECT 234.700 16.020 234.960 16.280 ;
        RECT 459.180 16.020 459.440 16.280 ;
      LAYER met2 ;
        RECT 490.920 1600.000 491.200 1604.000 ;
        RECT 490.980 1587.790 491.120 1600.000 ;
        RECT 459.180 1587.470 459.440 1587.790 ;
        RECT 490.920 1587.470 491.180 1587.790 ;
        RECT 459.240 16.310 459.380 1587.470 ;
        RECT 234.700 15.990 234.960 16.310 ;
        RECT 459.180 15.990 459.440 16.310 ;
        RECT 234.760 2.400 234.900 15.990 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 313.405 1586.865 313.575 1589.075 ;
      LAYER mcon ;
        RECT 313.405 1588.905 313.575 1589.075 ;
      LAYER met1 ;
        RECT 99.890 1589.060 100.210 1589.120 ;
        RECT 313.345 1589.060 313.635 1589.105 ;
        RECT 99.890 1588.920 313.635 1589.060 ;
        RECT 99.890 1588.860 100.210 1588.920 ;
        RECT 313.345 1588.875 313.635 1588.920 ;
        RECT 344.150 1588.040 344.470 1588.100 ;
        RECT 328.140 1587.900 344.470 1588.040 ;
        RECT 313.345 1587.020 313.635 1587.065 ;
        RECT 328.140 1587.020 328.280 1587.900 ;
        RECT 344.150 1587.840 344.470 1587.900 ;
        RECT 313.345 1586.880 328.280 1587.020 ;
        RECT 313.345 1586.835 313.635 1586.880 ;
        RECT 56.190 18.600 56.510 18.660 ;
        RECT 99.890 18.600 100.210 18.660 ;
        RECT 56.190 18.460 100.210 18.600 ;
        RECT 56.190 18.400 56.510 18.460 ;
        RECT 99.890 18.400 100.210 18.460 ;
      LAYER via ;
        RECT 99.920 1588.860 100.180 1589.120 ;
        RECT 344.180 1587.840 344.440 1588.100 ;
        RECT 56.220 18.400 56.480 18.660 ;
        RECT 99.920 18.400 100.180 18.660 ;
      LAYER met2 ;
        RECT 345.560 1600.450 345.840 1604.000 ;
        RECT 345.160 1600.310 345.840 1600.450 ;
        RECT 99.920 1588.830 100.180 1589.150 ;
        RECT 345.160 1588.890 345.300 1600.310 ;
        RECT 345.560 1600.000 345.840 1600.310 ;
        RECT 99.980 18.690 100.120 1588.830 ;
        RECT 344.240 1588.750 345.300 1588.890 ;
        RECT 344.240 1588.130 344.380 1588.750 ;
        RECT 344.180 1587.810 344.440 1588.130 ;
        RECT 56.220 18.370 56.480 18.690 ;
        RECT 99.920 18.370 100.180 18.690 ;
        RECT 56.280 2.400 56.420 18.370 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 1592.120 82.730 1592.180 ;
        RECT 364.850 1592.120 365.170 1592.180 ;
        RECT 82.410 1591.980 365.170 1592.120 ;
        RECT 82.410 1591.920 82.730 1591.980 ;
        RECT 364.850 1591.920 365.170 1591.980 ;
        RECT 80.110 20.640 80.430 20.700 ;
        RECT 82.410 20.640 82.730 20.700 ;
        RECT 80.110 20.500 82.730 20.640 ;
        RECT 80.110 20.440 80.430 20.500 ;
        RECT 82.410 20.440 82.730 20.500 ;
      LAYER via ;
        RECT 82.440 1591.920 82.700 1592.180 ;
        RECT 364.880 1591.920 365.140 1592.180 ;
        RECT 80.140 20.440 80.400 20.700 ;
        RECT 82.440 20.440 82.700 20.700 ;
      LAYER met2 ;
        RECT 364.880 1600.000 365.160 1604.000 ;
        RECT 364.940 1592.210 365.080 1600.000 ;
        RECT 82.440 1591.890 82.700 1592.210 ;
        RECT 364.880 1591.890 365.140 1592.210 ;
        RECT 82.500 20.730 82.640 1591.890 ;
        RECT 80.140 20.410 80.400 20.730 ;
        RECT 82.440 20.410 82.700 20.730 ;
        RECT 80.200 2.400 80.340 20.410 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 1592.460 109.870 1592.520 ;
        RECT 384.630 1592.460 384.950 1592.520 ;
        RECT 109.550 1592.320 384.950 1592.460 ;
        RECT 109.550 1592.260 109.870 1592.320 ;
        RECT 384.630 1592.260 384.950 1592.320 ;
        RECT 103.570 20.640 103.890 20.700 ;
        RECT 109.550 20.640 109.870 20.700 ;
        RECT 103.570 20.500 109.870 20.640 ;
        RECT 103.570 20.440 103.890 20.500 ;
        RECT 109.550 20.440 109.870 20.500 ;
      LAYER via ;
        RECT 109.580 1592.260 109.840 1592.520 ;
        RECT 384.660 1592.260 384.920 1592.520 ;
        RECT 103.600 20.440 103.860 20.700 ;
        RECT 109.580 20.440 109.840 20.700 ;
      LAYER met2 ;
        RECT 384.660 1600.000 384.940 1604.000 ;
        RECT 384.720 1592.550 384.860 1600.000 ;
        RECT 109.580 1592.230 109.840 1592.550 ;
        RECT 384.660 1592.230 384.920 1592.550 ;
        RECT 109.640 20.730 109.780 1592.230 ;
        RECT 103.600 20.410 103.860 20.730 ;
        RECT 109.580 20.410 109.840 20.730 ;
        RECT 103.660 2.400 103.800 20.410 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 1592.120 365.630 1592.180 ;
        RECT 403.950 1592.120 404.270 1592.180 ;
        RECT 365.310 1591.980 404.270 1592.120 ;
        RECT 365.310 1591.920 365.630 1591.980 ;
        RECT 403.950 1591.920 404.270 1591.980 ;
        RECT 362.550 1590.760 362.870 1590.820 ;
        RECT 365.310 1590.760 365.630 1590.820 ;
        RECT 362.550 1590.620 365.630 1590.760 ;
        RECT 362.550 1590.560 362.870 1590.620 ;
        RECT 365.310 1590.560 365.630 1590.620 ;
        RECT 127.490 19.960 127.810 20.020 ;
        RECT 362.550 19.960 362.870 20.020 ;
        RECT 127.490 19.820 362.870 19.960 ;
        RECT 127.490 19.760 127.810 19.820 ;
        RECT 362.550 19.760 362.870 19.820 ;
      LAYER via ;
        RECT 365.340 1591.920 365.600 1592.180 ;
        RECT 403.980 1591.920 404.240 1592.180 ;
        RECT 362.580 1590.560 362.840 1590.820 ;
        RECT 365.340 1590.560 365.600 1590.820 ;
        RECT 127.520 19.760 127.780 20.020 ;
        RECT 362.580 19.760 362.840 20.020 ;
      LAYER met2 ;
        RECT 403.980 1600.000 404.260 1604.000 ;
        RECT 404.040 1592.210 404.180 1600.000 ;
        RECT 365.340 1591.890 365.600 1592.210 ;
        RECT 403.980 1591.890 404.240 1592.210 ;
        RECT 365.400 1590.850 365.540 1591.890 ;
        RECT 362.580 1590.530 362.840 1590.850 ;
        RECT 365.340 1590.530 365.600 1590.850 ;
        RECT 362.640 20.050 362.780 1590.530 ;
        RECT 127.520 19.730 127.780 20.050 ;
        RECT 362.580 19.730 362.840 20.050 ;
        RECT 127.580 2.400 127.720 19.730 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 295.925 1587.545 296.095 1590.435 ;
      LAYER mcon ;
        RECT 295.925 1590.265 296.095 1590.435 ;
      LAYER met1 ;
        RECT 295.865 1590.420 296.155 1590.465 ;
        RECT 321.610 1590.420 321.930 1590.480 ;
        RECT 295.865 1590.280 321.930 1590.420 ;
        RECT 295.865 1590.235 296.155 1590.280 ;
        RECT 321.610 1590.220 321.930 1590.280 ;
        RECT 168.890 1587.700 169.210 1587.760 ;
        RECT 295.865 1587.700 296.155 1587.745 ;
        RECT 168.890 1587.560 296.155 1587.700 ;
        RECT 168.890 1587.500 169.210 1587.560 ;
        RECT 295.865 1587.515 296.155 1587.560 ;
        RECT 168.890 18.600 169.210 18.660 ;
        RECT 139.080 18.460 169.210 18.600 ;
        RECT 26.290 18.260 26.610 18.320 ;
        RECT 139.080 18.260 139.220 18.460 ;
        RECT 168.890 18.400 169.210 18.460 ;
        RECT 26.290 18.120 139.220 18.260 ;
        RECT 26.290 18.060 26.610 18.120 ;
      LAYER via ;
        RECT 321.640 1590.220 321.900 1590.480 ;
        RECT 168.920 1587.500 169.180 1587.760 ;
        RECT 26.320 18.060 26.580 18.320 ;
        RECT 168.920 18.400 169.180 18.660 ;
      LAYER met2 ;
        RECT 321.640 1600.000 321.920 1604.000 ;
        RECT 321.700 1590.510 321.840 1600.000 ;
        RECT 321.640 1590.190 321.900 1590.510 ;
        RECT 168.920 1587.470 169.180 1587.790 ;
        RECT 168.980 18.690 169.120 1587.470 ;
        RECT 168.920 18.370 169.180 18.690 ;
        RECT 26.320 18.030 26.580 18.350 ;
        RECT 26.380 2.400 26.520 18.030 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 131.245 16.065 131.415 17.255 ;
        RECT 179.085 16.065 179.255 17.255 ;
        RECT 180.005 14.705 180.175 17.255 ;
        RECT 226.465 14.705 226.635 17.255 ;
        RECT 276.605 15.045 276.775 17.255 ;
        RECT 299.605 15.045 299.775 17.595 ;
      LAYER mcon ;
        RECT 299.605 17.425 299.775 17.595 ;
        RECT 131.245 17.085 131.415 17.255 ;
        RECT 179.085 17.085 179.255 17.255 ;
        RECT 180.005 17.085 180.175 17.255 ;
        RECT 226.465 17.085 226.635 17.255 ;
        RECT 276.605 17.085 276.775 17.255 ;
      LAYER met1 ;
        RECT 32.270 17.580 32.590 17.640 ;
        RECT 299.545 17.580 299.835 17.625 ;
        RECT 32.270 17.440 44.000 17.580 ;
        RECT 32.270 17.380 32.590 17.440 ;
        RECT 43.860 17.240 44.000 17.440 ;
        RECT 299.545 17.440 314.480 17.580 ;
        RECT 299.545 17.395 299.835 17.440 ;
        RECT 131.185 17.240 131.475 17.285 ;
        RECT 43.860 17.100 131.475 17.240 ;
        RECT 131.185 17.055 131.475 17.100 ;
        RECT 179.025 17.240 179.315 17.285 ;
        RECT 179.945 17.240 180.235 17.285 ;
        RECT 179.025 17.100 180.235 17.240 ;
        RECT 179.025 17.055 179.315 17.100 ;
        RECT 179.945 17.055 180.235 17.100 ;
        RECT 226.405 17.240 226.695 17.285 ;
        RECT 276.545 17.240 276.835 17.285 ;
        RECT 226.405 17.100 276.835 17.240 ;
        RECT 226.405 17.055 226.695 17.100 ;
        RECT 276.545 17.055 276.835 17.100 ;
        RECT 314.340 16.900 314.480 17.440 ;
        RECT 324.830 16.900 325.150 16.960 ;
        RECT 314.340 16.760 325.150 16.900 ;
        RECT 324.830 16.700 325.150 16.760 ;
        RECT 131.185 16.220 131.475 16.265 ;
        RECT 179.025 16.220 179.315 16.265 ;
        RECT 131.185 16.080 179.315 16.220 ;
        RECT 131.185 16.035 131.475 16.080 ;
        RECT 179.025 16.035 179.315 16.080 ;
        RECT 276.545 15.200 276.835 15.245 ;
        RECT 299.545 15.200 299.835 15.245 ;
        RECT 276.545 15.060 299.835 15.200 ;
        RECT 276.545 15.015 276.835 15.060 ;
        RECT 299.545 15.015 299.835 15.060 ;
        RECT 179.945 14.860 180.235 14.905 ;
        RECT 226.405 14.860 226.695 14.905 ;
        RECT 179.945 14.720 226.695 14.860 ;
        RECT 179.945 14.675 180.235 14.720 ;
        RECT 226.405 14.675 226.695 14.720 ;
      LAYER via ;
        RECT 32.300 17.380 32.560 17.640 ;
        RECT 324.860 16.700 325.120 16.960 ;
      LAYER met2 ;
        RECT 326.240 1600.450 326.520 1604.000 ;
        RECT 324.920 1600.310 326.520 1600.450 ;
        RECT 32.300 17.350 32.560 17.670 ;
        RECT 32.360 2.400 32.500 17.350 ;
        RECT 324.920 16.990 325.060 1600.310 ;
        RECT 326.240 1600.000 326.520 1600.310 ;
        RECT 324.860 16.670 325.120 16.990 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.480 3243.600 684.050 3244.660 ;
        RECT 1331.480 3243.600 1334.050 3244.660 ;
        RECT 1931.480 3243.600 1934.050 3244.660 ;
        RECT 2581.480 3243.600 2584.050 3244.660 ;
        RECT 2581.480 2043.600 2584.050 2044.660 ;
        RECT 1552.430 1611.575 1555.000 1612.635 ;
      LAYER via3 ;
        RECT 682.500 3243.620 684.020 3244.630 ;
        RECT 1332.500 3243.620 1334.020 3244.630 ;
        RECT 1932.500 3243.620 1934.020 3244.630 ;
        RECT 2582.500 3243.620 2584.020 3244.630 ;
        RECT 2582.500 2043.620 2584.020 2044.630 ;
        RECT 1552.460 1611.605 1553.980 1612.615 ;
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 364.020 3271.235 367.020 3529.000 ;
        RECT 382.020 3271.235 385.020 3538.400 ;
        RECT 400.020 3271.235 403.020 3547.800 ;
        RECT 418.020 3271.235 421.020 3557.200 ;
        RECT 544.020 3271.235 547.020 3529.000 ;
        RECT 562.020 3271.235 565.020 3538.400 ;
        RECT 580.020 3271.235 583.020 3547.800 ;
        RECT 598.020 3271.235 601.020 3557.200 ;
        RECT 682.470 2803.670 684.070 3244.680 ;
        RECT 382.020 2715.000 385.020 2785.000 ;
        RECT 400.020 2715.000 403.020 2785.000 ;
        RECT 418.020 2715.000 421.020 2785.000 ;
        RECT 562.020 2715.000 565.020 2785.000 ;
        RECT 580.020 2715.000 583.020 2785.000 ;
        RECT 598.020 2715.000 601.020 2785.000 ;
        RECT 724.020 2715.000 727.020 3529.000 ;
        RECT 742.020 2715.000 745.020 3538.400 ;
        RECT 760.020 2715.000 763.020 3547.800 ;
        RECT 778.020 2715.000 781.020 3557.200 ;
        RECT 904.020 2715.000 907.020 3529.000 ;
        RECT 922.020 2715.000 925.020 3538.400 ;
        RECT 940.020 3271.235 943.020 3547.800 ;
        RECT 958.020 3271.235 961.020 3557.200 ;
        RECT 1084.020 3271.235 1087.020 3529.000 ;
        RECT 1102.020 3271.235 1105.020 3538.400 ;
        RECT 1120.020 3271.235 1123.020 3547.800 ;
        RECT 1138.020 3271.235 1141.020 3557.200 ;
        RECT 1264.020 3271.235 1267.020 3529.000 ;
        RECT 1282.020 3271.235 1285.020 3538.400 ;
        RECT 1300.020 3271.235 1303.020 3547.800 ;
        RECT 1318.020 3271.235 1321.020 3557.200 ;
        RECT 1332.470 2803.670 1334.070 3244.680 ;
        RECT 940.020 2715.000 943.020 2785.000 ;
        RECT 958.020 2715.000 961.020 2785.000 ;
        RECT 1102.020 2715.000 1105.020 2785.000 ;
        RECT 1120.020 2715.000 1123.020 2785.000 ;
        RECT 1138.020 2715.000 1141.020 2785.000 ;
        RECT 1282.020 2715.000 1285.020 2785.000 ;
        RECT 1300.020 2715.000 1303.020 2785.000 ;
        RECT 1318.020 2715.000 1321.020 2785.000 ;
        RECT 320.970 1610.640 322.570 2688.240 ;
        RECT 364.020 -9.320 367.020 1585.000 ;
        RECT 382.020 -18.720 385.020 1585.000 ;
        RECT 400.020 -28.120 403.020 1585.000 ;
        RECT 418.020 -37.520 421.020 1585.000 ;
        RECT 544.020 -9.320 547.020 1585.000 ;
        RECT 562.020 -18.720 565.020 1585.000 ;
        RECT 580.020 -28.120 583.020 1585.000 ;
        RECT 598.020 -37.520 601.020 1585.000 ;
        RECT 724.020 -9.320 727.020 1585.000 ;
        RECT 742.020 -18.720 745.020 1585.000 ;
        RECT 760.020 -28.120 763.020 1585.000 ;
        RECT 778.020 -37.520 781.020 1585.000 ;
        RECT 904.020 -9.320 907.020 1585.000 ;
        RECT 922.020 -18.720 925.020 1585.000 ;
        RECT 940.020 -28.120 943.020 1585.000 ;
        RECT 958.020 -37.520 961.020 1585.000 ;
        RECT 1084.020 -9.320 1087.020 1585.000 ;
        RECT 1102.020 -18.720 1105.020 1585.000 ;
        RECT 1120.020 -28.120 1123.020 1585.000 ;
        RECT 1138.020 -37.520 1141.020 1585.000 ;
        RECT 1264.020 -9.320 1267.020 1585.000 ;
        RECT 1282.020 -18.720 1285.020 1585.000 ;
        RECT 1300.020 -28.120 1303.020 1585.000 ;
        RECT 1318.020 -37.520 1321.020 1585.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1462.020 -18.720 1465.020 3538.400 ;
        RECT 1480.020 -28.120 1483.020 3547.800 ;
        RECT 1498.020 -37.520 1501.020 3557.200 ;
        RECT 1624.020 3271.235 1627.020 3529.000 ;
        RECT 1642.020 3271.235 1645.020 3538.400 ;
        RECT 1660.020 3271.235 1663.020 3547.800 ;
        RECT 1678.020 3271.235 1681.020 3557.200 ;
        RECT 1804.020 3271.235 1807.020 3529.000 ;
        RECT 1822.020 3271.235 1825.020 3538.400 ;
        RECT 1840.020 3271.235 1843.020 3547.800 ;
        RECT 1858.020 3271.235 1861.020 3557.200 ;
        RECT 1932.470 2803.670 1934.070 3244.680 ;
        RECT 1624.020 2071.235 1627.020 2785.000 ;
        RECT 1642.020 2071.235 1645.020 2785.000 ;
        RECT 1660.020 2071.235 1663.020 2785.000 ;
        RECT 1678.020 2071.235 1681.020 2785.000 ;
        RECT 1804.020 2071.235 1807.020 2785.000 ;
        RECT 1822.020 2071.235 1825.020 2785.000 ;
        RECT 1840.020 2071.235 1843.020 2785.000 ;
        RECT 1858.020 2071.235 1861.020 2785.000 ;
        RECT 1552.410 1611.555 1554.010 2052.565 ;
        RECT 1984.020 1515.000 1987.020 3529.000 ;
        RECT 2002.020 1515.000 2005.020 3538.400 ;
        RECT 2020.020 1515.000 2023.020 3547.800 ;
        RECT 2038.020 1515.000 2041.020 3557.200 ;
        RECT 2164.020 1515.000 2167.020 3529.000 ;
        RECT 2182.020 3271.235 2185.020 3538.400 ;
        RECT 2200.020 3271.235 2203.020 3547.800 ;
        RECT 2218.020 3271.235 2221.020 3557.200 ;
        RECT 2344.020 3271.235 2347.020 3529.000 ;
        RECT 2362.020 3271.235 2365.020 3538.400 ;
        RECT 2380.020 3271.235 2383.020 3547.800 ;
        RECT 2398.020 3271.235 2401.020 3557.200 ;
        RECT 2524.020 3271.235 2527.020 3529.000 ;
        RECT 2542.020 3271.235 2545.020 3538.400 ;
        RECT 2560.020 3271.235 2563.020 3547.800 ;
        RECT 2578.020 3271.235 2581.020 3557.200 ;
        RECT 2582.470 2803.670 2584.070 3244.680 ;
        RECT 2182.020 2071.235 2185.020 2785.000 ;
        RECT 2200.020 2071.235 2203.020 2785.000 ;
        RECT 2218.020 2071.235 2221.020 2785.000 ;
        RECT 2344.020 2071.235 2347.020 2785.000 ;
        RECT 2362.020 2071.235 2365.020 2785.000 ;
        RECT 2380.020 2071.235 2383.020 2785.000 ;
        RECT 2398.020 2071.235 2401.020 2785.000 ;
        RECT 2524.020 2071.235 2527.020 2785.000 ;
        RECT 2542.020 2071.235 2545.020 2785.000 ;
        RECT 2560.020 2071.235 2563.020 2785.000 ;
        RECT 2578.020 2071.235 2581.020 2785.000 ;
        RECT 2582.470 1603.670 2584.070 2044.680 ;
        RECT 1570.970 410.640 1572.570 1488.240 ;
        RECT 1624.020 -9.320 1627.020 385.000 ;
        RECT 1642.020 -18.720 1645.020 385.000 ;
        RECT 1660.020 -28.120 1663.020 385.000 ;
        RECT 1678.020 -37.520 1681.020 385.000 ;
        RECT 1804.020 -9.320 1807.020 385.000 ;
        RECT 1822.020 -18.720 1825.020 385.000 ;
        RECT 1840.020 -28.120 1843.020 385.000 ;
        RECT 1858.020 -37.520 1861.020 385.000 ;
        RECT 1984.020 -9.320 1987.020 385.000 ;
        RECT 2002.020 -18.720 2005.020 385.000 ;
        RECT 2020.020 -28.120 2023.020 385.000 ;
        RECT 2038.020 -37.520 2041.020 385.000 ;
        RECT 2164.020 -9.320 2167.020 385.000 ;
        RECT 2182.020 -18.720 2185.020 385.000 ;
        RECT 2200.020 -28.120 2203.020 385.000 ;
        RECT 2218.020 -37.520 2221.020 385.000 ;
        RECT 2344.020 -9.320 2347.020 385.000 ;
        RECT 2362.020 -18.720 2365.020 385.000 ;
        RECT 2380.020 -28.120 2383.020 385.000 ;
        RECT 2398.020 -37.520 2401.020 385.000 ;
        RECT 2524.020 -9.320 2527.020 385.000 ;
        RECT 2542.020 -18.720 2545.020 385.000 ;
        RECT 2560.020 -28.120 2563.020 385.000 ;
        RECT 2578.020 -37.520 2581.020 385.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 682.680 3125.090 683.860 3126.270 ;
        RECT 682.680 3123.490 683.860 3124.670 ;
        RECT 682.680 3107.090 683.860 3108.270 ;
        RECT 682.680 3105.490 683.860 3106.670 ;
        RECT 682.680 3089.090 683.860 3090.270 ;
        RECT 682.680 3087.490 683.860 3088.670 ;
        RECT 682.680 3071.090 683.860 3072.270 ;
        RECT 682.680 3069.490 683.860 3070.670 ;
        RECT 682.680 2945.090 683.860 2946.270 ;
        RECT 682.680 2943.490 683.860 2944.670 ;
        RECT 682.680 2927.090 683.860 2928.270 ;
        RECT 682.680 2925.490 683.860 2926.670 ;
        RECT 682.680 2909.090 683.860 2910.270 ;
        RECT 682.680 2907.490 683.860 2908.670 ;
        RECT 682.680 2891.090 683.860 2892.270 ;
        RECT 682.680 2889.490 683.860 2890.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 1332.680 3125.090 1333.860 3126.270 ;
        RECT 1332.680 3123.490 1333.860 3124.670 ;
        RECT 1332.680 3107.090 1333.860 3108.270 ;
        RECT 1332.680 3105.490 1333.860 3106.670 ;
        RECT 1332.680 3089.090 1333.860 3090.270 ;
        RECT 1332.680 3087.490 1333.860 3088.670 ;
        RECT 1332.680 3071.090 1333.860 3072.270 ;
        RECT 1332.680 3069.490 1333.860 3070.670 ;
        RECT 1332.680 2945.090 1333.860 2946.270 ;
        RECT 1332.680 2943.490 1333.860 2944.670 ;
        RECT 1332.680 2927.090 1333.860 2928.270 ;
        RECT 1332.680 2925.490 1333.860 2926.670 ;
        RECT 1332.680 2909.090 1333.860 2910.270 ;
        RECT 1332.680 2907.490 1333.860 2908.670 ;
        RECT 1332.680 2891.090 1333.860 2892.270 ;
        RECT 1332.680 2889.490 1333.860 2890.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 321.180 2585.090 322.360 2586.270 ;
        RECT 321.180 2583.490 322.360 2584.670 ;
        RECT 321.180 2567.090 322.360 2568.270 ;
        RECT 321.180 2565.490 322.360 2566.670 ;
        RECT 321.180 2549.090 322.360 2550.270 ;
        RECT 321.180 2547.490 322.360 2548.670 ;
        RECT 321.180 2531.090 322.360 2532.270 ;
        RECT 321.180 2529.490 322.360 2530.670 ;
        RECT 321.180 2405.090 322.360 2406.270 ;
        RECT 321.180 2403.490 322.360 2404.670 ;
        RECT 321.180 2387.090 322.360 2388.270 ;
        RECT 321.180 2385.490 322.360 2386.670 ;
        RECT 321.180 2369.090 322.360 2370.270 ;
        RECT 321.180 2367.490 322.360 2368.670 ;
        RECT 321.180 2351.090 322.360 2352.270 ;
        RECT 321.180 2349.490 322.360 2350.670 ;
        RECT 321.180 2225.090 322.360 2226.270 ;
        RECT 321.180 2223.490 322.360 2224.670 ;
        RECT 321.180 2207.090 322.360 2208.270 ;
        RECT 321.180 2205.490 322.360 2206.670 ;
        RECT 321.180 2189.090 322.360 2190.270 ;
        RECT 321.180 2187.490 322.360 2188.670 ;
        RECT 321.180 2171.090 322.360 2172.270 ;
        RECT 321.180 2169.490 322.360 2170.670 ;
        RECT 321.180 2045.090 322.360 2046.270 ;
        RECT 321.180 2043.490 322.360 2044.670 ;
        RECT 321.180 2027.090 322.360 2028.270 ;
        RECT 321.180 2025.490 322.360 2026.670 ;
        RECT 321.180 2009.090 322.360 2010.270 ;
        RECT 321.180 2007.490 322.360 2008.670 ;
        RECT 321.180 1991.090 322.360 1992.270 ;
        RECT 321.180 1989.490 322.360 1990.670 ;
        RECT 321.180 1865.090 322.360 1866.270 ;
        RECT 321.180 1863.490 322.360 1864.670 ;
        RECT 321.180 1847.090 322.360 1848.270 ;
        RECT 321.180 1845.490 322.360 1846.670 ;
        RECT 321.180 1829.090 322.360 1830.270 ;
        RECT 321.180 1827.490 322.360 1828.670 ;
        RECT 321.180 1811.090 322.360 1812.270 ;
        RECT 321.180 1809.490 322.360 1810.670 ;
        RECT 321.180 1685.090 322.360 1686.270 ;
        RECT 321.180 1683.490 322.360 1684.670 ;
        RECT 321.180 1667.090 322.360 1668.270 ;
        RECT 321.180 1665.490 322.360 1666.670 ;
        RECT 321.180 1649.090 322.360 1650.270 ;
        RECT 321.180 1647.490 322.360 1648.670 ;
        RECT 321.180 1631.090 322.360 1632.270 ;
        RECT 321.180 1629.490 322.360 1630.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1932.680 3125.090 1933.860 3126.270 ;
        RECT 1932.680 3123.490 1933.860 3124.670 ;
        RECT 1932.680 3107.090 1933.860 3108.270 ;
        RECT 1932.680 3105.490 1933.860 3106.670 ;
        RECT 1932.680 3089.090 1933.860 3090.270 ;
        RECT 1932.680 3087.490 1933.860 3088.670 ;
        RECT 1932.680 3071.090 1933.860 3072.270 ;
        RECT 1932.680 3069.490 1933.860 3070.670 ;
        RECT 1932.680 2945.090 1933.860 2946.270 ;
        RECT 1932.680 2943.490 1933.860 2944.670 ;
        RECT 1932.680 2927.090 1933.860 2928.270 ;
        RECT 1932.680 2925.490 1933.860 2926.670 ;
        RECT 1932.680 2909.090 1933.860 2910.270 ;
        RECT 1932.680 2907.490 1933.860 2908.670 ;
        RECT 1932.680 2891.090 1933.860 2892.270 ;
        RECT 1932.680 2889.490 1933.860 2890.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1552.620 2045.090 1553.800 2046.270 ;
        RECT 1552.620 2043.490 1553.800 2044.670 ;
        RECT 1552.620 2027.090 1553.800 2028.270 ;
        RECT 1552.620 2025.490 1553.800 2026.670 ;
        RECT 1552.620 2009.090 1553.800 2010.270 ;
        RECT 1552.620 2007.490 1553.800 2008.670 ;
        RECT 1552.620 1991.090 1553.800 1992.270 ;
        RECT 1552.620 1989.490 1553.800 1990.670 ;
        RECT 1552.620 1865.090 1553.800 1866.270 ;
        RECT 1552.620 1863.490 1553.800 1864.670 ;
        RECT 1552.620 1847.090 1553.800 1848.270 ;
        RECT 1552.620 1845.490 1553.800 1846.670 ;
        RECT 1552.620 1829.090 1553.800 1830.270 ;
        RECT 1552.620 1827.490 1553.800 1828.670 ;
        RECT 1552.620 1811.090 1553.800 1812.270 ;
        RECT 1552.620 1809.490 1553.800 1810.670 ;
        RECT 1552.620 1685.090 1553.800 1686.270 ;
        RECT 1552.620 1683.490 1553.800 1684.670 ;
        RECT 1552.620 1667.090 1553.800 1668.270 ;
        RECT 1552.620 1665.490 1553.800 1666.670 ;
        RECT 1552.620 1649.090 1553.800 1650.270 ;
        RECT 1552.620 1647.490 1553.800 1648.670 ;
        RECT 1552.620 1631.090 1553.800 1632.270 ;
        RECT 1552.620 1629.490 1553.800 1630.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2582.680 3125.090 2583.860 3126.270 ;
        RECT 2582.680 3123.490 2583.860 3124.670 ;
        RECT 2582.680 3107.090 2583.860 3108.270 ;
        RECT 2582.680 3105.490 2583.860 3106.670 ;
        RECT 2582.680 3089.090 2583.860 3090.270 ;
        RECT 2582.680 3087.490 2583.860 3088.670 ;
        RECT 2582.680 3071.090 2583.860 3072.270 ;
        RECT 2582.680 3069.490 2583.860 3070.670 ;
        RECT 2582.680 2945.090 2583.860 2946.270 ;
        RECT 2582.680 2943.490 2583.860 2944.670 ;
        RECT 2582.680 2927.090 2583.860 2928.270 ;
        RECT 2582.680 2925.490 2583.860 2926.670 ;
        RECT 2582.680 2909.090 2583.860 2910.270 ;
        RECT 2582.680 2907.490 2583.860 2908.670 ;
        RECT 2582.680 2891.090 2583.860 2892.270 ;
        RECT 2582.680 2889.490 2583.860 2890.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2582.680 2027.090 2583.860 2028.270 ;
        RECT 2582.680 2025.490 2583.860 2026.670 ;
        RECT 2582.680 2009.090 2583.860 2010.270 ;
        RECT 2582.680 2007.490 2583.860 2008.670 ;
        RECT 2582.680 1991.090 2583.860 1992.270 ;
        RECT 2582.680 1989.490 2583.860 1990.670 ;
        RECT 2582.680 1865.090 2583.860 1866.270 ;
        RECT 2582.680 1863.490 2583.860 1864.670 ;
        RECT 2582.680 1847.090 2583.860 1848.270 ;
        RECT 2582.680 1845.490 2583.860 1846.670 ;
        RECT 2582.680 1829.090 2583.860 1830.270 ;
        RECT 2582.680 1827.490 2583.860 1828.670 ;
        RECT 2582.680 1811.090 2583.860 1812.270 ;
        RECT 2582.680 1809.490 2583.860 1810.670 ;
        RECT 2582.680 1685.090 2583.860 1686.270 ;
        RECT 2582.680 1683.490 2583.860 1684.670 ;
        RECT 2582.680 1667.090 2583.860 1668.270 ;
        RECT 2582.680 1665.490 2583.860 1666.670 ;
        RECT 2582.680 1649.090 2583.860 1650.270 ;
        RECT 2582.680 1647.490 2583.860 1648.670 ;
        RECT 2582.680 1631.090 2583.860 1632.270 ;
        RECT 2582.680 1629.490 2583.860 1630.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1571.180 1469.090 1572.360 1470.270 ;
        RECT 1571.180 1467.490 1572.360 1468.670 ;
        RECT 1571.180 1451.090 1572.360 1452.270 ;
        RECT 1571.180 1449.490 1572.360 1450.670 ;
        RECT 1571.180 1325.090 1572.360 1326.270 ;
        RECT 1571.180 1323.490 1572.360 1324.670 ;
        RECT 1571.180 1307.090 1572.360 1308.270 ;
        RECT 1571.180 1305.490 1572.360 1306.670 ;
        RECT 1571.180 1289.090 1572.360 1290.270 ;
        RECT 1571.180 1287.490 1572.360 1288.670 ;
        RECT 1571.180 1271.090 1572.360 1272.270 ;
        RECT 1571.180 1269.490 1572.360 1270.670 ;
        RECT 1571.180 1145.090 1572.360 1146.270 ;
        RECT 1571.180 1143.490 1572.360 1144.670 ;
        RECT 1571.180 1127.090 1572.360 1128.270 ;
        RECT 1571.180 1125.490 1572.360 1126.670 ;
        RECT 1571.180 1109.090 1572.360 1110.270 ;
        RECT 1571.180 1107.490 1572.360 1108.670 ;
        RECT 1571.180 1091.090 1572.360 1092.270 ;
        RECT 1571.180 1089.490 1572.360 1090.670 ;
        RECT 1571.180 965.090 1572.360 966.270 ;
        RECT 1571.180 963.490 1572.360 964.670 ;
        RECT 1571.180 947.090 1572.360 948.270 ;
        RECT 1571.180 945.490 1572.360 946.670 ;
        RECT 1571.180 929.090 1572.360 930.270 ;
        RECT 1571.180 927.490 1572.360 928.670 ;
        RECT 1571.180 911.090 1572.360 912.270 ;
        RECT 1571.180 909.490 1572.360 910.670 ;
        RECT 1571.180 785.090 1572.360 786.270 ;
        RECT 1571.180 783.490 1572.360 784.670 ;
        RECT 1571.180 767.090 1572.360 768.270 ;
        RECT 1571.180 765.490 1572.360 766.670 ;
        RECT 1571.180 749.090 1572.360 750.270 ;
        RECT 1571.180 747.490 1572.360 748.670 ;
        RECT 1571.180 731.090 1572.360 732.270 ;
        RECT 1571.180 729.490 1572.360 730.670 ;
        RECT 1571.180 605.090 1572.360 606.270 ;
        RECT 1571.180 603.490 1572.360 604.670 ;
        RECT 1571.180 587.090 1572.360 588.270 ;
        RECT 1571.180 585.490 1572.360 586.670 ;
        RECT 1571.180 569.090 1572.360 570.270 ;
        RECT 1571.180 567.490 1572.360 568.670 ;
        RECT 1571.180 551.090 1572.360 552.270 ;
        RECT 1571.180 549.490 1572.360 550.670 ;
        RECT 1571.180 425.090 1572.360 426.270 ;
        RECT 1571.180 423.490 1572.360 424.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 682.470 3126.380 684.070 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 1332.470 3126.380 1334.070 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1932.470 3126.380 1934.070 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2582.470 3126.380 2584.070 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 682.470 3123.370 684.070 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 1332.470 3123.370 1334.070 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1932.470 3123.370 1934.070 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2582.470 3123.370 2584.070 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 682.470 3108.380 684.070 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 1332.470 3108.380 1334.070 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1932.470 3108.380 1934.070 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2582.470 3108.380 2584.070 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 682.470 3105.370 684.070 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 1332.470 3105.370 1334.070 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1932.470 3105.370 1934.070 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2582.470 3105.370 2584.070 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 682.470 3090.380 684.070 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1332.470 3090.380 1334.070 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1932.470 3090.380 1934.070 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2582.470 3090.380 2584.070 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 682.470 3087.370 684.070 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1332.470 3087.370 1334.070 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1932.470 3087.370 1934.070 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2582.470 3087.370 2584.070 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 682.470 3072.380 684.070 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1332.470 3072.380 1334.070 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1932.470 3072.380 1934.070 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2582.470 3072.380 2584.070 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 682.470 3069.370 684.070 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1332.470 3069.370 1334.070 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1932.470 3069.370 1934.070 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2582.470 3069.370 2584.070 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 682.470 2946.380 684.070 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 1332.470 2946.380 1334.070 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1932.470 2946.380 1934.070 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2582.470 2946.380 2584.070 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 682.470 2943.370 684.070 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 1332.470 2943.370 1334.070 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1932.470 2943.370 1934.070 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2582.470 2943.370 2584.070 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 682.470 2928.380 684.070 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 1332.470 2928.380 1334.070 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1932.470 2928.380 1934.070 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2582.470 2928.380 2584.070 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 682.470 2925.370 684.070 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 1332.470 2925.370 1334.070 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1932.470 2925.370 1934.070 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2582.470 2925.370 2584.070 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 682.470 2910.380 684.070 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1332.470 2910.380 1334.070 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1932.470 2910.380 1934.070 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2582.470 2910.380 2584.070 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 682.470 2907.370 684.070 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1332.470 2907.370 1334.070 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1932.470 2907.370 1934.070 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2582.470 2907.370 2584.070 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 682.470 2892.380 684.070 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1332.470 2892.380 1334.070 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1932.470 2892.380 1934.070 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2582.470 2892.380 2584.070 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 682.470 2889.370 684.070 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1332.470 2889.370 1334.070 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1932.470 2889.370 1934.070 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2582.470 2889.370 2584.070 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 320.970 2586.380 322.570 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 320.970 2583.370 322.570 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 320.970 2568.380 322.570 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 320.970 2565.370 322.570 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 320.970 2550.380 322.570 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 320.970 2547.370 322.570 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 320.970 2532.380 322.570 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 320.970 2529.370 322.570 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 320.970 2406.380 322.570 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 320.970 2403.370 322.570 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 320.970 2388.380 322.570 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 320.970 2385.370 322.570 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 320.970 2370.380 322.570 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 320.970 2367.370 322.570 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 320.970 2352.380 322.570 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 320.970 2349.370 322.570 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 320.970 2226.380 322.570 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 320.970 2223.370 322.570 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 320.970 2208.380 322.570 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 320.970 2205.370 322.570 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 320.970 2190.380 322.570 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 320.970 2187.370 322.570 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 320.970 2172.380 322.570 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 320.970 2169.370 322.570 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 320.970 2046.380 322.570 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1552.410 2046.380 1554.010 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 320.970 2043.370 322.570 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1552.410 2043.370 1554.010 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 320.970 2028.380 322.570 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1552.410 2028.380 1554.010 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2582.470 2028.380 2584.070 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 320.970 2025.370 322.570 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1552.410 2025.370 1554.010 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2582.470 2025.370 2584.070 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 320.970 2010.380 322.570 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1552.410 2010.380 1554.010 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2582.470 2010.380 2584.070 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 320.970 2007.370 322.570 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1552.410 2007.370 1554.010 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2582.470 2007.370 2584.070 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 320.970 1992.380 322.570 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1552.410 1992.380 1554.010 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2582.470 1992.380 2584.070 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 320.970 1989.370 322.570 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1552.410 1989.370 1554.010 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2582.470 1989.370 2584.070 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 320.970 1866.380 322.570 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1552.410 1866.380 1554.010 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2582.470 1866.380 2584.070 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 320.970 1863.370 322.570 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1552.410 1863.370 1554.010 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2582.470 1863.370 2584.070 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 320.970 1848.380 322.570 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1552.410 1848.380 1554.010 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2582.470 1848.380 2584.070 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 320.970 1845.370 322.570 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1552.410 1845.370 1554.010 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2582.470 1845.370 2584.070 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 320.970 1830.380 322.570 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1552.410 1830.380 1554.010 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2582.470 1830.380 2584.070 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 320.970 1827.370 322.570 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1552.410 1827.370 1554.010 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2582.470 1827.370 2584.070 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 320.970 1812.380 322.570 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1552.410 1812.380 1554.010 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2582.470 1812.380 2584.070 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 320.970 1809.370 322.570 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1552.410 1809.370 1554.010 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2582.470 1809.370 2584.070 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 320.970 1686.380 322.570 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1552.410 1686.380 1554.010 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2582.470 1686.380 2584.070 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 320.970 1683.370 322.570 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1552.410 1683.370 1554.010 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2582.470 1683.370 2584.070 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 320.970 1668.380 322.570 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1552.410 1668.380 1554.010 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2582.470 1668.380 2584.070 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 320.970 1665.370 322.570 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1552.410 1665.370 1554.010 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2582.470 1665.370 2584.070 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 320.970 1650.380 322.570 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1552.410 1650.380 1554.010 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2582.470 1650.380 2584.070 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 320.970 1647.370 322.570 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1552.410 1647.370 1554.010 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2582.470 1647.370 2584.070 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 320.970 1632.380 322.570 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1552.410 1632.380 1554.010 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2582.470 1632.380 2584.070 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 320.970 1629.370 322.570 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1552.410 1629.370 1554.010 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2582.470 1629.370 2584.070 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1570.970 1470.380 1572.570 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1570.970 1467.370 1572.570 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1570.970 1452.380 1572.570 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1570.970 1449.370 1572.570 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1570.970 1326.380 1572.570 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1570.970 1323.370 1572.570 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1570.970 1308.380 1572.570 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1570.970 1305.370 1572.570 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1570.970 1290.380 1572.570 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1570.970 1287.370 1572.570 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1570.970 1272.380 1572.570 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1570.970 1269.370 1572.570 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1570.970 1146.380 1572.570 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1570.970 1143.370 1572.570 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1570.970 1128.380 1572.570 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1570.970 1125.370 1572.570 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1570.970 1110.380 1572.570 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1570.970 1107.370 1572.570 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1570.970 1092.380 1572.570 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1570.970 1089.370 1572.570 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1570.970 966.380 1572.570 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1570.970 963.370 1572.570 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1570.970 948.380 1572.570 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1570.970 945.370 1572.570 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1570.970 930.380 1572.570 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1570.970 927.370 1572.570 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1570.970 912.380 1572.570 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1570.970 909.370 1572.570 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1570.970 786.380 1572.570 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1570.970 783.370 1572.570 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1570.970 768.380 1572.570 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1570.970 765.370 1572.570 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1570.970 750.380 1572.570 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1570.970 747.370 1572.570 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1570.970 732.380 1572.570 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1570.970 729.370 1572.570 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1570.970 606.380 1572.570 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1570.970 603.370 1572.570 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1570.970 588.380 1572.570 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1570.970 585.370 1572.570 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1570.970 570.380 1572.570 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1570.970 567.370 1572.570 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1570.970 552.380 1572.570 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1570.970 549.370 1572.570 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1570.970 426.380 1572.570 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1570.970 423.370 1572.570 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.040 3251.235 686.300 3252.140 ;
        RECT 1331.040 3251.235 1336.300 3252.140 ;
        RECT 1931.040 3251.235 1936.300 3252.140 ;
        RECT 2581.040 3251.235 2586.300 3252.140 ;
        RECT 681.480 3250.400 686.300 3251.235 ;
        RECT 1331.480 3250.400 1336.300 3251.235 ;
        RECT 1931.480 3250.400 1936.300 3251.235 ;
        RECT 2581.480 3250.400 2586.300 3251.235 ;
        RECT 2581.040 2051.235 2586.300 2052.140 ;
        RECT 2581.480 2050.400 2586.300 2051.235 ;
        RECT 1550.180 1605.000 1555.000 1605.835 ;
        RECT 1550.180 1604.095 1555.440 1605.000 ;
      LAYER via3 ;
        RECT 684.720 3250.440 686.240 3252.050 ;
        RECT 1334.720 3250.440 1336.240 3252.050 ;
        RECT 1934.720 3250.440 1936.240 3252.050 ;
        RECT 2584.720 3250.440 2586.240 3252.050 ;
        RECT 2584.720 2050.440 2586.240 2052.050 ;
        RECT 1550.240 1604.185 1551.760 1605.795 ;
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 292.020 3271.235 295.020 3538.400 ;
        RECT 310.020 3271.235 313.020 3547.800 ;
        RECT 328.020 3271.235 331.020 3557.200 ;
        RECT 454.020 3271.235 457.020 3529.000 ;
        RECT 472.020 3271.235 475.020 3538.400 ;
        RECT 490.020 3271.235 493.020 3547.800 ;
        RECT 508.020 3271.235 511.020 3557.200 ;
        RECT 634.020 3271.235 637.020 3529.000 ;
        RECT 652.020 3271.235 655.020 3538.400 ;
        RECT 670.020 3271.235 673.020 3547.800 ;
        RECT 688.020 3271.235 691.020 3557.200 ;
        RECT 684.690 2804.060 686.310 3252.140 ;
        RECT 814.020 2715.000 817.020 3529.000 ;
        RECT 832.020 2715.000 835.020 3538.400 ;
        RECT 850.020 2715.000 853.020 3547.800 ;
        RECT 868.020 2715.000 871.020 3557.200 ;
        RECT 994.020 3271.235 997.020 3529.000 ;
        RECT 1012.020 3271.235 1015.020 3538.400 ;
        RECT 1030.020 3271.235 1033.020 3547.800 ;
        RECT 1048.020 3271.235 1051.020 3557.200 ;
        RECT 1174.020 3271.235 1177.020 3529.000 ;
        RECT 1192.020 3271.235 1195.020 3538.400 ;
        RECT 1210.020 3271.235 1213.020 3547.800 ;
        RECT 1228.020 3271.235 1231.020 3557.200 ;
        RECT 1334.690 2804.060 1336.310 3252.140 ;
        RECT 1354.020 2715.000 1357.020 3529.000 ;
        RECT 1372.020 2715.000 1375.020 3538.400 ;
        RECT 1390.020 2715.000 1393.020 3547.800 ;
        RECT 1408.020 2715.000 1411.020 3557.200 ;
        RECT 1534.020 3271.235 1537.020 3529.000 ;
        RECT 1552.020 3271.235 1555.020 3538.400 ;
        RECT 1570.020 3271.235 1573.020 3547.800 ;
        RECT 1588.020 3271.235 1591.020 3557.200 ;
        RECT 1714.020 3271.235 1717.020 3529.000 ;
        RECT 1732.020 3271.235 1735.020 3538.400 ;
        RECT 1750.020 3271.235 1753.020 3547.800 ;
        RECT 1768.020 3271.235 1771.020 3557.200 ;
        RECT 1894.020 3271.235 1897.020 3529.000 ;
        RECT 1912.020 3271.235 1915.020 3538.400 ;
        RECT 1930.020 3271.235 1933.020 3547.800 ;
        RECT 1948.020 3271.235 1951.020 3557.200 ;
        RECT 1934.690 2804.060 1936.310 3252.140 ;
        RECT 397.770 1610.640 399.370 2688.240 ;
        RECT 1534.020 2071.235 1537.020 2785.000 ;
        RECT 1552.020 2071.235 1555.020 2785.000 ;
        RECT 1570.020 2071.235 1573.020 2785.000 ;
        RECT 1588.020 2071.235 1591.020 2785.000 ;
        RECT 1714.020 2071.235 1717.020 2785.000 ;
        RECT 1732.020 2071.235 1735.020 2785.000 ;
        RECT 1750.020 2071.235 1753.020 2785.000 ;
        RECT 1768.020 2071.235 1771.020 2785.000 ;
        RECT 1894.020 2071.235 1897.020 2785.000 ;
        RECT 1912.020 2071.235 1915.020 2785.000 ;
        RECT 1930.020 2071.235 1933.020 2785.000 ;
        RECT 1948.020 2071.235 1951.020 2785.000 ;
        RECT 1550.170 1604.095 1551.790 2052.175 ;
        RECT 292.020 -18.720 295.020 1585.000 ;
        RECT 310.020 -28.120 313.020 1585.000 ;
        RECT 328.020 -37.520 331.020 1585.000 ;
        RECT 454.020 -9.320 457.020 1585.000 ;
        RECT 472.020 -18.720 475.020 1585.000 ;
        RECT 490.020 -28.120 493.020 1585.000 ;
        RECT 508.020 -37.520 511.020 1585.000 ;
        RECT 634.020 -9.320 637.020 1585.000 ;
        RECT 652.020 -18.720 655.020 1585.000 ;
        RECT 670.020 -28.120 673.020 1585.000 ;
        RECT 688.020 -37.520 691.020 1585.000 ;
        RECT 814.020 -9.320 817.020 1585.000 ;
        RECT 832.020 -18.720 835.020 1585.000 ;
        RECT 850.020 -28.120 853.020 1585.000 ;
        RECT 868.020 -37.520 871.020 1585.000 ;
        RECT 994.020 -9.320 997.020 1585.000 ;
        RECT 1012.020 -18.720 1015.020 1585.000 ;
        RECT 1030.020 -28.120 1033.020 1585.000 ;
        RECT 1048.020 -37.520 1051.020 1585.000 ;
        RECT 1174.020 -9.320 1177.020 1585.000 ;
        RECT 1192.020 -18.720 1195.020 1585.000 ;
        RECT 1210.020 -28.120 1213.020 1585.000 ;
        RECT 1228.020 -37.520 1231.020 1585.000 ;
        RECT 1354.020 -9.320 1357.020 1585.000 ;
        RECT 1372.020 -18.720 1375.020 1585.000 ;
        RECT 1390.020 -28.120 1393.020 1585.000 ;
        RECT 1408.020 -37.520 1411.020 1585.000 ;
        RECT 1534.020 1515.000 1537.020 1585.000 ;
        RECT 1552.020 1515.000 1555.020 1585.000 ;
        RECT 1570.020 1515.000 1573.020 1585.000 ;
        RECT 1714.020 1515.000 1717.020 1585.000 ;
        RECT 1732.020 1515.000 1735.020 1585.000 ;
        RECT 1750.020 1515.000 1753.020 1585.000 ;
        RECT 1894.020 1515.000 1897.020 1585.000 ;
        RECT 1912.020 1515.000 1915.020 1585.000 ;
        RECT 1930.020 1515.000 1933.020 1585.000 ;
        RECT 2074.020 1515.000 2077.020 3529.000 ;
        RECT 2092.020 1515.000 2095.020 3538.400 ;
        RECT 2110.020 1515.000 2113.020 3547.800 ;
        RECT 2128.020 1515.000 2131.020 3557.200 ;
        RECT 2254.020 3271.235 2257.020 3529.000 ;
        RECT 2272.020 3271.235 2275.020 3538.400 ;
        RECT 2290.020 3271.235 2293.020 3547.800 ;
        RECT 2308.020 3271.235 2311.020 3557.200 ;
        RECT 2434.020 3271.235 2437.020 3529.000 ;
        RECT 2452.020 3271.235 2455.020 3538.400 ;
        RECT 2470.020 3271.235 2473.020 3547.800 ;
        RECT 2488.020 3271.235 2491.020 3557.200 ;
        RECT 2584.690 2804.060 2586.310 3252.140 ;
        RECT 2254.020 2071.235 2257.020 2785.000 ;
        RECT 2272.020 2071.235 2275.020 2785.000 ;
        RECT 2290.020 2071.235 2293.020 2785.000 ;
        RECT 2308.020 2071.235 2311.020 2785.000 ;
        RECT 2434.020 2071.235 2437.020 2785.000 ;
        RECT 2452.020 2071.235 2455.020 2785.000 ;
        RECT 2470.020 2071.235 2473.020 2785.000 ;
        RECT 2488.020 2071.235 2491.020 2785.000 ;
        RECT 2584.690 1604.060 2586.310 2052.140 ;
        RECT 2254.020 1515.000 2257.020 1585.000 ;
        RECT 2272.020 1515.000 2275.020 1585.000 ;
        RECT 2290.020 1515.000 2293.020 1585.000 ;
        RECT 2434.020 1515.000 2437.020 1585.000 ;
        RECT 2452.020 1515.000 2455.020 1585.000 ;
        RECT 2470.020 1515.000 2473.020 1585.000 ;
        RECT 2614.020 1515.000 2617.020 3529.000 ;
        RECT 2632.020 1515.000 2635.020 3538.400 ;
        RECT 2650.020 1515.000 2653.020 3547.800 ;
        RECT 1647.770 410.640 1649.370 1488.240 ;
        RECT 1534.020 -9.320 1537.020 385.000 ;
        RECT 1552.020 -18.720 1555.020 385.000 ;
        RECT 1570.020 -28.120 1573.020 385.000 ;
        RECT 1588.020 -37.520 1591.020 385.000 ;
        RECT 1714.020 -9.320 1717.020 385.000 ;
        RECT 1732.020 -18.720 1735.020 385.000 ;
        RECT 1750.020 -28.120 1753.020 385.000 ;
        RECT 1768.020 -37.520 1771.020 385.000 ;
        RECT 1894.020 -9.320 1897.020 385.000 ;
        RECT 1912.020 -18.720 1915.020 385.000 ;
        RECT 1930.020 -28.120 1933.020 385.000 ;
        RECT 1948.020 -37.520 1951.020 385.000 ;
        RECT 2074.020 -9.320 2077.020 385.000 ;
        RECT 2092.020 -18.720 2095.020 385.000 ;
        RECT 2110.020 -28.120 2113.020 385.000 ;
        RECT 2128.020 -37.520 2131.020 385.000 ;
        RECT 2254.020 -9.320 2257.020 385.000 ;
        RECT 2272.020 -18.720 2275.020 385.000 ;
        RECT 2290.020 -28.120 2293.020 385.000 ;
        RECT 2308.020 -37.520 2311.020 385.000 ;
        RECT 2434.020 -9.320 2437.020 385.000 ;
        RECT 2452.020 -18.720 2455.020 385.000 ;
        RECT 2470.020 -28.120 2473.020 385.000 ;
        RECT 2488.020 -37.520 2491.020 385.000 ;
        RECT 2614.020 -9.320 2617.020 385.000 ;
        RECT 2632.020 -18.720 2635.020 385.000 ;
        RECT 2650.020 -28.120 2653.020 385.000 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 684.910 3215.090 686.090 3216.270 ;
        RECT 684.910 3213.490 686.090 3214.670 ;
        RECT 684.910 3197.090 686.090 3198.270 ;
        RECT 684.910 3195.490 686.090 3196.670 ;
        RECT 684.910 3179.090 686.090 3180.270 ;
        RECT 684.910 3177.490 686.090 3178.670 ;
        RECT 684.910 3161.090 686.090 3162.270 ;
        RECT 684.910 3159.490 686.090 3160.670 ;
        RECT 684.910 3035.090 686.090 3036.270 ;
        RECT 684.910 3033.490 686.090 3034.670 ;
        RECT 684.910 3017.090 686.090 3018.270 ;
        RECT 684.910 3015.490 686.090 3016.670 ;
        RECT 684.910 2999.090 686.090 3000.270 ;
        RECT 684.910 2997.490 686.090 2998.670 ;
        RECT 684.910 2981.090 686.090 2982.270 ;
        RECT 684.910 2979.490 686.090 2980.670 ;
        RECT 684.910 2855.090 686.090 2856.270 ;
        RECT 684.910 2853.490 686.090 2854.670 ;
        RECT 684.910 2837.090 686.090 2838.270 ;
        RECT 684.910 2835.490 686.090 2836.670 ;
        RECT 684.910 2819.090 686.090 2820.270 ;
        RECT 684.910 2817.490 686.090 2818.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1334.910 3215.090 1336.090 3216.270 ;
        RECT 1334.910 3213.490 1336.090 3214.670 ;
        RECT 1334.910 3197.090 1336.090 3198.270 ;
        RECT 1334.910 3195.490 1336.090 3196.670 ;
        RECT 1334.910 3179.090 1336.090 3180.270 ;
        RECT 1334.910 3177.490 1336.090 3178.670 ;
        RECT 1334.910 3161.090 1336.090 3162.270 ;
        RECT 1334.910 3159.490 1336.090 3160.670 ;
        RECT 1334.910 3035.090 1336.090 3036.270 ;
        RECT 1334.910 3033.490 1336.090 3034.670 ;
        RECT 1334.910 3017.090 1336.090 3018.270 ;
        RECT 1334.910 3015.490 1336.090 3016.670 ;
        RECT 1334.910 2999.090 1336.090 3000.270 ;
        RECT 1334.910 2997.490 1336.090 2998.670 ;
        RECT 1334.910 2981.090 1336.090 2982.270 ;
        RECT 1334.910 2979.490 1336.090 2980.670 ;
        RECT 1334.910 2855.090 1336.090 2856.270 ;
        RECT 1334.910 2853.490 1336.090 2854.670 ;
        RECT 1334.910 2837.090 1336.090 2838.270 ;
        RECT 1334.910 2835.490 1336.090 2836.670 ;
        RECT 1334.910 2819.090 1336.090 2820.270 ;
        RECT 1334.910 2817.490 1336.090 2818.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1934.910 3215.090 1936.090 3216.270 ;
        RECT 1934.910 3213.490 1936.090 3214.670 ;
        RECT 1934.910 3197.090 1936.090 3198.270 ;
        RECT 1934.910 3195.490 1936.090 3196.670 ;
        RECT 1934.910 3179.090 1936.090 3180.270 ;
        RECT 1934.910 3177.490 1936.090 3178.670 ;
        RECT 1934.910 3161.090 1936.090 3162.270 ;
        RECT 1934.910 3159.490 1936.090 3160.670 ;
        RECT 1934.910 3035.090 1936.090 3036.270 ;
        RECT 1934.910 3033.490 1936.090 3034.670 ;
        RECT 1934.910 3017.090 1936.090 3018.270 ;
        RECT 1934.910 3015.490 1936.090 3016.670 ;
        RECT 1934.910 2999.090 1936.090 3000.270 ;
        RECT 1934.910 2997.490 1936.090 2998.670 ;
        RECT 1934.910 2981.090 1936.090 2982.270 ;
        RECT 1934.910 2979.490 1936.090 2980.670 ;
        RECT 1934.910 2855.090 1936.090 2856.270 ;
        RECT 1934.910 2853.490 1936.090 2854.670 ;
        RECT 1934.910 2837.090 1936.090 2838.270 ;
        RECT 1934.910 2835.490 1936.090 2836.670 ;
        RECT 1934.910 2819.090 1936.090 2820.270 ;
        RECT 1934.910 2817.490 1936.090 2818.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 397.980 2675.090 399.160 2676.270 ;
        RECT 397.980 2673.490 399.160 2674.670 ;
        RECT 397.980 2657.090 399.160 2658.270 ;
        RECT 397.980 2655.490 399.160 2656.670 ;
        RECT 397.980 2639.090 399.160 2640.270 ;
        RECT 397.980 2637.490 399.160 2638.670 ;
        RECT 397.980 2621.090 399.160 2622.270 ;
        RECT 397.980 2619.490 399.160 2620.670 ;
        RECT 397.980 2495.090 399.160 2496.270 ;
        RECT 397.980 2493.490 399.160 2494.670 ;
        RECT 397.980 2477.090 399.160 2478.270 ;
        RECT 397.980 2475.490 399.160 2476.670 ;
        RECT 397.980 2459.090 399.160 2460.270 ;
        RECT 397.980 2457.490 399.160 2458.670 ;
        RECT 397.980 2441.090 399.160 2442.270 ;
        RECT 397.980 2439.490 399.160 2440.670 ;
        RECT 397.980 2315.090 399.160 2316.270 ;
        RECT 397.980 2313.490 399.160 2314.670 ;
        RECT 397.980 2297.090 399.160 2298.270 ;
        RECT 397.980 2295.490 399.160 2296.670 ;
        RECT 397.980 2279.090 399.160 2280.270 ;
        RECT 397.980 2277.490 399.160 2278.670 ;
        RECT 397.980 2261.090 399.160 2262.270 ;
        RECT 397.980 2259.490 399.160 2260.670 ;
        RECT 397.980 2135.090 399.160 2136.270 ;
        RECT 397.980 2133.490 399.160 2134.670 ;
        RECT 397.980 2117.090 399.160 2118.270 ;
        RECT 397.980 2115.490 399.160 2116.670 ;
        RECT 397.980 2099.090 399.160 2100.270 ;
        RECT 397.980 2097.490 399.160 2098.670 ;
        RECT 397.980 2081.090 399.160 2082.270 ;
        RECT 397.980 2079.490 399.160 2080.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 397.980 1955.090 399.160 1956.270 ;
        RECT 397.980 1953.490 399.160 1954.670 ;
        RECT 397.980 1937.090 399.160 1938.270 ;
        RECT 397.980 1935.490 399.160 1936.670 ;
        RECT 397.980 1919.090 399.160 1920.270 ;
        RECT 397.980 1917.490 399.160 1918.670 ;
        RECT 397.980 1901.090 399.160 1902.270 ;
        RECT 397.980 1899.490 399.160 1900.670 ;
        RECT 397.980 1775.090 399.160 1776.270 ;
        RECT 397.980 1773.490 399.160 1774.670 ;
        RECT 397.980 1757.090 399.160 1758.270 ;
        RECT 397.980 1755.490 399.160 1756.670 ;
        RECT 397.980 1739.090 399.160 1740.270 ;
        RECT 397.980 1737.490 399.160 1738.670 ;
        RECT 397.980 1721.090 399.160 1722.270 ;
        RECT 397.980 1719.490 399.160 1720.670 ;
        RECT 1550.390 1955.090 1551.570 1956.270 ;
        RECT 1550.390 1953.490 1551.570 1954.670 ;
        RECT 1550.390 1937.090 1551.570 1938.270 ;
        RECT 1550.390 1935.490 1551.570 1936.670 ;
        RECT 1550.390 1919.090 1551.570 1920.270 ;
        RECT 1550.390 1917.490 1551.570 1918.670 ;
        RECT 1550.390 1901.090 1551.570 1902.270 ;
        RECT 1550.390 1899.490 1551.570 1900.670 ;
        RECT 1550.390 1775.090 1551.570 1776.270 ;
        RECT 1550.390 1773.490 1551.570 1774.670 ;
        RECT 1550.390 1757.090 1551.570 1758.270 ;
        RECT 1550.390 1755.490 1551.570 1756.670 ;
        RECT 1550.390 1739.090 1551.570 1740.270 ;
        RECT 1550.390 1737.490 1551.570 1738.670 ;
        RECT 1550.390 1721.090 1551.570 1722.270 ;
        RECT 1550.390 1719.490 1551.570 1720.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2584.910 3215.090 2586.090 3216.270 ;
        RECT 2584.910 3213.490 2586.090 3214.670 ;
        RECT 2584.910 3197.090 2586.090 3198.270 ;
        RECT 2584.910 3195.490 2586.090 3196.670 ;
        RECT 2584.910 3179.090 2586.090 3180.270 ;
        RECT 2584.910 3177.490 2586.090 3178.670 ;
        RECT 2584.910 3161.090 2586.090 3162.270 ;
        RECT 2584.910 3159.490 2586.090 3160.670 ;
        RECT 2584.910 3035.090 2586.090 3036.270 ;
        RECT 2584.910 3033.490 2586.090 3034.670 ;
        RECT 2584.910 3017.090 2586.090 3018.270 ;
        RECT 2584.910 3015.490 2586.090 3016.670 ;
        RECT 2584.910 2999.090 2586.090 3000.270 ;
        RECT 2584.910 2997.490 2586.090 2998.670 ;
        RECT 2584.910 2981.090 2586.090 2982.270 ;
        RECT 2584.910 2979.490 2586.090 2980.670 ;
        RECT 2584.910 2855.090 2586.090 2856.270 ;
        RECT 2584.910 2853.490 2586.090 2854.670 ;
        RECT 2584.910 2837.090 2586.090 2838.270 ;
        RECT 2584.910 2835.490 2586.090 2836.670 ;
        RECT 2584.910 2819.090 2586.090 2820.270 ;
        RECT 2584.910 2817.490 2586.090 2818.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2584.910 1955.090 2586.090 1956.270 ;
        RECT 2584.910 1953.490 2586.090 1954.670 ;
        RECT 2584.910 1937.090 2586.090 1938.270 ;
        RECT 2584.910 1935.490 2586.090 1936.670 ;
        RECT 2584.910 1919.090 2586.090 1920.270 ;
        RECT 2584.910 1917.490 2586.090 1918.670 ;
        RECT 2584.910 1901.090 2586.090 1902.270 ;
        RECT 2584.910 1899.490 2586.090 1900.670 ;
        RECT 2584.910 1775.090 2586.090 1776.270 ;
        RECT 2584.910 1773.490 2586.090 1774.670 ;
        RECT 2584.910 1757.090 2586.090 1758.270 ;
        RECT 2584.910 1755.490 2586.090 1756.670 ;
        RECT 2584.910 1739.090 2586.090 1740.270 ;
        RECT 2584.910 1737.490 2586.090 1738.670 ;
        RECT 2584.910 1721.090 2586.090 1722.270 ;
        RECT 2584.910 1719.490 2586.090 1720.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1647.980 1415.090 1649.160 1416.270 ;
        RECT 1647.980 1413.490 1649.160 1414.670 ;
        RECT 1647.980 1397.090 1649.160 1398.270 ;
        RECT 1647.980 1395.490 1649.160 1396.670 ;
        RECT 1647.980 1379.090 1649.160 1380.270 ;
        RECT 1647.980 1377.490 1649.160 1378.670 ;
        RECT 1647.980 1361.090 1649.160 1362.270 ;
        RECT 1647.980 1359.490 1649.160 1360.670 ;
        RECT 1647.980 1235.090 1649.160 1236.270 ;
        RECT 1647.980 1233.490 1649.160 1234.670 ;
        RECT 1647.980 1217.090 1649.160 1218.270 ;
        RECT 1647.980 1215.490 1649.160 1216.670 ;
        RECT 1647.980 1199.090 1649.160 1200.270 ;
        RECT 1647.980 1197.490 1649.160 1198.670 ;
        RECT 1647.980 1181.090 1649.160 1182.270 ;
        RECT 1647.980 1179.490 1649.160 1180.670 ;
        RECT 1647.980 1055.090 1649.160 1056.270 ;
        RECT 1647.980 1053.490 1649.160 1054.670 ;
        RECT 1647.980 1037.090 1649.160 1038.270 ;
        RECT 1647.980 1035.490 1649.160 1036.670 ;
        RECT 1647.980 1019.090 1649.160 1020.270 ;
        RECT 1647.980 1017.490 1649.160 1018.670 ;
        RECT 1647.980 1001.090 1649.160 1002.270 ;
        RECT 1647.980 999.490 1649.160 1000.670 ;
        RECT 1647.980 875.090 1649.160 876.270 ;
        RECT 1647.980 873.490 1649.160 874.670 ;
        RECT 1647.980 857.090 1649.160 858.270 ;
        RECT 1647.980 855.490 1649.160 856.670 ;
        RECT 1647.980 839.090 1649.160 840.270 ;
        RECT 1647.980 837.490 1649.160 838.670 ;
        RECT 1647.980 821.090 1649.160 822.270 ;
        RECT 1647.980 819.490 1649.160 820.670 ;
        RECT 1647.980 695.090 1649.160 696.270 ;
        RECT 1647.980 693.490 1649.160 694.670 ;
        RECT 1647.980 677.090 1649.160 678.270 ;
        RECT 1647.980 675.490 1649.160 676.670 ;
        RECT 1647.980 659.090 1649.160 660.270 ;
        RECT 1647.980 657.490 1649.160 658.670 ;
        RECT 1647.980 641.090 1649.160 642.270 ;
        RECT 1647.980 639.490 1649.160 640.670 ;
        RECT 1647.980 515.090 1649.160 516.270 ;
        RECT 1647.980 513.490 1649.160 514.670 ;
        RECT 1647.980 497.090 1649.160 498.270 ;
        RECT 1647.980 495.490 1649.160 496.670 ;
        RECT 1647.980 479.090 1649.160 480.270 ;
        RECT 1647.980 477.490 1649.160 478.670 ;
        RECT 1647.980 461.090 1649.160 462.270 ;
        RECT 1647.980 459.490 1649.160 460.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 684.690 3216.380 686.310 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1334.690 3216.380 1336.310 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1934.690 3216.380 1936.310 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2584.690 3216.380 2586.310 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 684.690 3213.370 686.310 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1334.690 3213.370 1336.310 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1934.690 3213.370 1936.310 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2584.690 3213.370 2586.310 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 684.690 3198.380 686.310 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1334.690 3198.380 1336.310 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1934.690 3198.380 1936.310 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2584.690 3198.380 2586.310 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 684.690 3195.370 686.310 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1334.690 3195.370 1336.310 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1934.690 3195.370 1936.310 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2584.690 3195.370 2586.310 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 684.690 3180.380 686.310 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1334.690 3180.380 1336.310 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1934.690 3180.380 1936.310 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2584.690 3180.380 2586.310 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 684.690 3177.370 686.310 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1334.690 3177.370 1336.310 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1934.690 3177.370 1936.310 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2584.690 3177.370 2586.310 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 684.690 3162.380 686.310 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 1334.690 3162.380 1336.310 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1934.690 3162.380 1936.310 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2584.690 3162.380 2586.310 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 684.690 3159.370 686.310 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 1334.690 3159.370 1336.310 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1934.690 3159.370 1936.310 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2584.690 3159.370 2586.310 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 684.690 3036.380 686.310 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1334.690 3036.380 1336.310 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1934.690 3036.380 1936.310 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2584.690 3036.380 2586.310 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 684.690 3033.370 686.310 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1334.690 3033.370 1336.310 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1934.690 3033.370 1936.310 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2584.690 3033.370 2586.310 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 684.690 3018.380 686.310 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1334.690 3018.380 1336.310 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1934.690 3018.380 1936.310 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2584.690 3018.380 2586.310 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 684.690 3015.370 686.310 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1334.690 3015.370 1336.310 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1934.690 3015.370 1936.310 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2584.690 3015.370 2586.310 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 684.690 3000.380 686.310 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1334.690 3000.380 1336.310 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1934.690 3000.380 1936.310 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2584.690 3000.380 2586.310 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 684.690 2997.370 686.310 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1334.690 2997.370 1336.310 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1934.690 2997.370 1936.310 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2584.690 2997.370 2586.310 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 684.690 2982.380 686.310 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 1334.690 2982.380 1336.310 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1934.690 2982.380 1936.310 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2584.690 2982.380 2586.310 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 684.690 2979.370 686.310 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 1334.690 2979.370 1336.310 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1934.690 2979.370 1936.310 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2584.690 2979.370 2586.310 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 684.690 2856.380 686.310 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1334.690 2856.380 1336.310 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1934.690 2856.380 1936.310 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2584.690 2856.380 2586.310 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 684.690 2853.370 686.310 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1334.690 2853.370 1336.310 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1934.690 2853.370 1936.310 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2584.690 2853.370 2586.310 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 684.690 2838.380 686.310 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1334.690 2838.380 1336.310 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1934.690 2838.380 1936.310 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2584.690 2838.380 2586.310 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 684.690 2835.370 686.310 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1334.690 2835.370 1336.310 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1934.690 2835.370 1936.310 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2584.690 2835.370 2586.310 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 684.690 2820.380 686.310 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1334.690 2820.380 1336.310 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1934.690 2820.380 1936.310 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2584.690 2820.380 2586.310 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 684.690 2817.370 686.310 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1334.690 2817.370 1336.310 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1934.690 2817.370 1936.310 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2584.690 2817.370 2586.310 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 397.770 2676.380 399.370 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 397.770 2673.370 399.370 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 397.770 2658.380 399.370 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 397.770 2655.370 399.370 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 397.770 2640.380 399.370 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 397.770 2637.370 399.370 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 397.770 2622.380 399.370 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 397.770 2619.370 399.370 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 397.770 2496.380 399.370 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 397.770 2493.370 399.370 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 397.770 2478.380 399.370 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 397.770 2475.370 399.370 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 397.770 2460.380 399.370 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 397.770 2457.370 399.370 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 397.770 2442.380 399.370 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 397.770 2439.370 399.370 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 397.770 2316.380 399.370 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 397.770 2313.370 399.370 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 397.770 2298.380 399.370 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 397.770 2295.370 399.370 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 397.770 2280.380 399.370 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 397.770 2277.370 399.370 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 397.770 2262.380 399.370 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 397.770 2259.370 399.370 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 397.770 2136.380 399.370 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 397.770 2133.370 399.370 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 397.770 2118.380 399.370 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 397.770 2115.370 399.370 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 397.770 2100.380 399.370 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 397.770 2097.370 399.370 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 397.770 2082.380 399.370 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 397.770 2079.370 399.370 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 397.770 1956.380 399.370 1956.390 ;
        RECT 1550.170 1956.380 1551.790 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2584.690 1956.380 2586.310 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 397.770 1953.370 399.370 1953.380 ;
        RECT 1550.170 1953.370 1551.790 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2584.690 1953.370 2586.310 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 397.770 1938.380 399.370 1938.390 ;
        RECT 1550.170 1938.380 1551.790 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2584.690 1938.380 2586.310 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 397.770 1935.370 399.370 1935.380 ;
        RECT 1550.170 1935.370 1551.790 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2584.690 1935.370 2586.310 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 397.770 1920.380 399.370 1920.390 ;
        RECT 1550.170 1920.380 1551.790 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2584.690 1920.380 2586.310 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 397.770 1917.370 399.370 1917.380 ;
        RECT 1550.170 1917.370 1551.790 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2584.690 1917.370 2586.310 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 397.770 1902.380 399.370 1902.390 ;
        RECT 1550.170 1902.380 1551.790 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2584.690 1902.380 2586.310 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 397.770 1899.370 399.370 1899.380 ;
        RECT 1550.170 1899.370 1551.790 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2584.690 1899.370 2586.310 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 397.770 1776.380 399.370 1776.390 ;
        RECT 1550.170 1776.380 1551.790 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2584.690 1776.380 2586.310 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 397.770 1773.370 399.370 1773.380 ;
        RECT 1550.170 1773.370 1551.790 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2584.690 1773.370 2586.310 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 397.770 1758.380 399.370 1758.390 ;
        RECT 1550.170 1758.380 1551.790 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2584.690 1758.380 2586.310 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 397.770 1755.370 399.370 1755.380 ;
        RECT 1550.170 1755.370 1551.790 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2584.690 1755.370 2586.310 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 397.770 1740.380 399.370 1740.390 ;
        RECT 1550.170 1740.380 1551.790 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2584.690 1740.380 2586.310 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 397.770 1737.370 399.370 1737.380 ;
        RECT 1550.170 1737.370 1551.790 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2584.690 1737.370 2586.310 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 397.770 1722.380 399.370 1722.390 ;
        RECT 1550.170 1722.380 1551.790 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2584.690 1722.380 2586.310 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 397.770 1719.370 399.370 1719.380 ;
        RECT 1550.170 1719.370 1551.790 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2584.690 1719.370 2586.310 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1647.770 1416.380 1649.370 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1647.770 1413.370 1649.370 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1647.770 1398.380 1649.370 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1647.770 1395.370 1649.370 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1647.770 1380.380 1649.370 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1647.770 1377.370 1649.370 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1647.770 1362.380 1649.370 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1647.770 1359.370 1649.370 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1647.770 1236.380 1649.370 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1647.770 1233.370 1649.370 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1647.770 1218.380 1649.370 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1647.770 1215.370 1649.370 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1647.770 1200.380 1649.370 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1647.770 1197.370 1649.370 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1647.770 1182.380 1649.370 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1647.770 1179.370 1649.370 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1647.770 1056.380 1649.370 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1647.770 1053.370 1649.370 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1647.770 1038.380 1649.370 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1647.770 1035.370 1649.370 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1647.770 1020.380 1649.370 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1647.770 1017.370 1649.370 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1647.770 1002.380 1649.370 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1647.770 999.370 1649.370 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1647.770 876.380 1649.370 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1647.770 873.370 1649.370 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1647.770 858.380 1649.370 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1647.770 855.370 1649.370 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1647.770 840.380 1649.370 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1647.770 837.370 1649.370 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1647.770 822.380 1649.370 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1647.770 819.370 1649.370 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1647.770 696.380 1649.370 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1647.770 693.370 1649.370 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1647.770 678.380 1649.370 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1647.770 675.370 1649.370 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1647.770 660.380 1649.370 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1647.770 657.370 1649.370 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1647.770 642.380 1649.370 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1647.770 639.370 1649.370 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1647.770 516.380 1649.370 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1647.770 513.370 1649.370 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1647.770 498.380 1649.370 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1647.770 495.370 1649.370 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1647.770 480.380 1649.370 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1647.770 477.370 1649.370 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1647.770 462.380 1649.370 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1647.770 459.370 1649.370 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 676.345 3263.065 676.515 3263.915 ;
        RECT 724.185 3263.065 724.355 3263.915 ;
        RECT 772.945 3263.065 773.115 3263.915 ;
        RECT 820.785 3263.065 820.955 3263.915 ;
        RECT 966.145 3263.065 966.315 3263.915 ;
        RECT 1013.985 3263.065 1014.155 3263.915 ;
        RECT 1062.745 3263.065 1062.915 3263.915 ;
        RECT 1110.585 3263.065 1110.755 3263.915 ;
        RECT 1159.345 3263.065 1159.515 3263.915 ;
        RECT 1207.185 3263.065 1207.355 3263.915 ;
        RECT 1317.585 3263.745 1317.755 3266.975 ;
        RECT 1014.445 3252.865 1014.615 3253.715 ;
      LAYER li1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER li1 ;
        RECT 724.645 3250.825 724.815 3252.015 ;
        RECT 748.565 3250.825 748.735 3252.015 ;
        RECT 772.945 3251.165 773.115 3252.355 ;
        RECT 883.345 3251.845 883.515 3252.695 ;
        RECT 917.845 3251.845 918.015 3252.695 ;
        RECT 959.245 3251.845 959.415 3252.695 ;
        RECT 1055.845 3252.185 1056.015 3253.715 ;
        RECT 1103.685 3252.185 1103.855 3253.035 ;
        RECT 1111.045 3252.865 1111.215 3253.715 ;
        RECT 1152.445 3252.185 1152.615 3253.715 ;
        RECT 1200.285 3252.185 1200.455 3253.035 ;
        RECT 1207.645 3252.185 1207.815 3253.375 ;
        RECT 1231.565 3252.185 1231.735 3253.375 ;
        RECT 1594.045 3253.205 1594.215 3254.055 ;
        RECT 1559.085 3252.865 1559.715 3253.035 ;
        RECT 1641.885 3252.865 1642.055 3254.055 ;
        RECT 1690.645 3253.205 1690.815 3254.055 ;
        RECT 1655.685 3252.865 1656.315 3253.035 ;
        RECT 1738.485 3252.865 1738.655 3254.055 ;
        RECT 1787.245 3253.205 1787.415 3254.055 ;
        RECT 1752.285 3252.865 1752.915 3253.035 ;
        RECT 1835.085 3252.865 1835.255 3254.055 ;
        RECT 2270.245 3253.205 2270.415 3254.055 ;
        RECT 1849.345 3252.865 1849.975 3253.035 ;
        RECT 2235.285 3252.865 2235.915 3253.035 ;
        RECT 2318.085 3252.865 2318.255 3254.055 ;
        RECT 2366.845 3253.205 2367.015 3254.055 ;
        RECT 2331.885 3252.865 2332.515 3253.035 ;
        RECT 2414.685 3252.865 2414.855 3254.055 ;
        RECT 2463.445 3253.205 2463.615 3254.055 ;
        RECT 2428.485 3252.865 2429.115 3253.035 ;
        RECT 2511.285 3252.865 2511.455 3254.055 ;
        RECT 2525.545 3252.865 2526.175 3253.035 ;
        RECT 1269.285 3252.185 1270.375 3252.355 ;
        RECT 1270.205 3251.505 1270.375 3252.185 ;
        RECT 1297.345 3251.845 1297.515 3252.695 ;
      LAYER li1 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER li1 ;
        RECT 1352.545 3251.165 1352.715 3252.015 ;
        RECT 1400.385 3250.825 1400.555 3252.015 ;
        RECT 1449.145 3251.505 1449.315 3252.355 ;
        RECT 1496.985 3251.505 1497.155 3252.695 ;
      LAYER li1 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER li1 ;
        RECT 1932.145 3251.165 1932.315 3252.355 ;
        RECT 1948.245 3251.165 1948.415 3252.695 ;
        RECT 1980.445 3251.505 1980.615 3252.695 ;
        RECT 2028.745 3250.825 2028.915 3251.675 ;
        RECT 2076.585 3250.825 2076.755 3252.015 ;
        RECT 2125.345 3251.505 2125.515 3252.355 ;
        RECT 2173.185 3251.505 2173.355 3252.695 ;
      LAYER li1 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER li1 ;
        RECT 391.145 2791.145 391.315 2793.015 ;
        RECT 477.625 2789.445 477.795 2792.335 ;
        RECT 504.765 2791.825 504.935 2793.695 ;
        RECT 1060.445 2791.825 1060.615 2794.375 ;
        RECT 1511.245 2793.525 1511.415 2794.375 ;
        RECT 1583.465 2793.525 1583.635 2794.375 ;
        RECT 1690.645 2793.525 1690.815 2795.055 ;
        RECT 1449.145 2792.165 1449.315 2793.015 ;
        RECT 1510.785 2792.845 1511.415 2793.015 ;
        RECT 1538.845 2792.165 1539.015 2793.015 ;
        RECT 1559.085 2792.505 1559.715 2792.675 ;
        RECT 1587.145 2792.505 1587.315 2793.355 ;
        RECT 1634.985 2792.505 1635.155 2793.355 ;
        RECT 1738.485 2793.185 1738.655 2795.055 ;
        RECT 1828.185 2793.185 1828.355 2794.375 ;
        RECT 1848.885 2793.185 1849.055 2794.375 ;
        RECT 2187.445 2793.185 2187.615 2794.375 ;
        RECT 2255.985 2793.185 2256.155 2794.375 ;
        RECT 2279.445 2794.205 2281.455 2794.375 ;
        RECT 2279.445 2793.525 2279.615 2794.205 ;
        RECT 1559.085 2792.165 1559.255 2792.505 ;
        RECT 1486.865 2788.085 1487.035 2789.275 ;
        RECT 1511.245 2788.425 1511.415 2791.655 ;
        RECT 1654.765 2789.785 1654.935 2791.655 ;
        RECT 1704.445 2790.125 1704.615 2792.675 ;
        RECT 1535.165 2788.085 1535.335 2788.935 ;
        RECT 1669.945 2788.085 1670.115 2789.955 ;
        RECT 1870.045 2788.425 1870.215 2791.315 ;
        RECT 1917.425 2788.255 1917.595 2791.315 ;
        RECT 2090.845 2788.765 2091.475 2788.935 ;
        RECT 2091.305 2788.425 2091.475 2788.765 ;
        RECT 1917.425 2788.085 1918.055 2788.255 ;
        RECT 1931.685 2788.085 1932.315 2788.255 ;
        RECT 1738.485 2787.745 1739.115 2787.915 ;
        RECT 1738.485 2787.405 1738.655 2787.745 ;
        RECT 1980.445 2787.065 1980.615 2787.915 ;
        RECT 2028.285 2787.065 2028.455 2788.255 ;
        RECT 2042.085 2788.085 2042.715 2788.255 ;
        RECT 2138.685 2788.085 2138.855 2791.655 ;
        RECT 2139.145 2788.085 2139.315 2791.655 ;
        RECT 2181.465 2787.745 2181.635 2791.655 ;
        RECT 2210.905 2788.765 2211.075 2792.675 ;
        RECT 2280.825 2792.165 2280.995 2793.695 ;
        RECT 2347.985 2792.335 2348.155 2794.035 ;
        RECT 2252.305 2788.425 2256.155 2788.595 ;
        RECT 2262.885 2788.425 2263.055 2791.655 ;
        RECT 2252.305 2787.745 2252.475 2788.425 ;
        RECT 2267.485 2788.085 2267.655 2788.935 ;
        RECT 2334.185 2788.255 2334.355 2792.335 ;
        RECT 2347.065 2792.165 2348.155 2792.335 ;
        RECT 2333.265 2788.085 2334.355 2788.255 ;
      LAYER li1 ;
        RECT 305.450 1610.795 1395.045 2688.085 ;
      LAYER li1 ;
        RECT 1409.125 2045.865 1409.295 2056.575 ;
      LAYER li1 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
        RECT 1555.450 410.795 2645.045 1488.085 ;
      LAYER mcon ;
        RECT 1317.585 3266.805 1317.755 3266.975 ;
        RECT 676.345 3263.745 676.515 3263.915 ;
        RECT 724.185 3263.745 724.355 3263.915 ;
        RECT 772.945 3263.745 773.115 3263.915 ;
        RECT 820.785 3263.745 820.955 3263.915 ;
        RECT 966.145 3263.745 966.315 3263.915 ;
        RECT 1013.985 3263.745 1014.155 3263.915 ;
        RECT 1062.745 3263.745 1062.915 3263.915 ;
        RECT 1110.585 3263.745 1110.755 3263.915 ;
        RECT 1159.345 3263.745 1159.515 3263.915 ;
        RECT 1207.185 3263.745 1207.355 3263.915 ;
        RECT 1594.045 3253.885 1594.215 3254.055 ;
        RECT 1014.445 3253.545 1014.615 3253.715 ;
        RECT 1055.845 3253.545 1056.015 3253.715 ;
        RECT 883.345 3252.525 883.515 3252.695 ;
        RECT 772.945 3252.185 773.115 3252.355 ;
        RECT 724.645 3251.845 724.815 3252.015 ;
        RECT 748.565 3251.845 748.735 3252.015 ;
        RECT 917.845 3252.525 918.015 3252.695 ;
        RECT 959.245 3252.525 959.415 3252.695 ;
        RECT 1111.045 3253.545 1111.215 3253.715 ;
        RECT 1103.685 3252.865 1103.855 3253.035 ;
        RECT 1152.445 3253.545 1152.615 3253.715 ;
        RECT 1207.645 3253.205 1207.815 3253.375 ;
        RECT 1200.285 3252.865 1200.455 3253.035 ;
        RECT 1231.565 3253.205 1231.735 3253.375 ;
        RECT 1641.885 3253.885 1642.055 3254.055 ;
        RECT 1690.645 3253.885 1690.815 3254.055 ;
        RECT 1738.485 3253.885 1738.655 3254.055 ;
        RECT 1787.245 3253.885 1787.415 3254.055 ;
        RECT 1835.085 3253.885 1835.255 3254.055 ;
        RECT 2270.245 3253.885 2270.415 3254.055 ;
        RECT 2318.085 3253.885 2318.255 3254.055 ;
        RECT 2366.845 3253.885 2367.015 3254.055 ;
        RECT 2414.685 3253.885 2414.855 3254.055 ;
        RECT 2463.445 3253.885 2463.615 3254.055 ;
        RECT 2511.285 3253.885 2511.455 3254.055 ;
        RECT 1559.545 3252.865 1559.715 3253.035 ;
        RECT 1656.145 3252.865 1656.315 3253.035 ;
        RECT 1752.745 3252.865 1752.915 3253.035 ;
        RECT 1849.805 3252.865 1849.975 3253.035 ;
        RECT 2235.745 3252.865 2235.915 3253.035 ;
        RECT 2332.345 3252.865 2332.515 3253.035 ;
        RECT 2428.945 3252.865 2429.115 3253.035 ;
        RECT 2526.005 3252.865 2526.175 3253.035 ;
        RECT 1297.345 3252.525 1297.515 3252.695 ;
        RECT 1496.985 3252.525 1497.155 3252.695 ;
        RECT 1449.145 3252.185 1449.315 3252.355 ;
        RECT 1352.545 3251.845 1352.715 3252.015 ;
        RECT 1400.385 3251.845 1400.555 3252.015 ;
        RECT 1948.245 3252.525 1948.415 3252.695 ;
        RECT 1932.145 3252.185 1932.315 3252.355 ;
        RECT 1980.445 3252.525 1980.615 3252.695 ;
        RECT 2173.185 3252.525 2173.355 3252.695 ;
        RECT 2125.345 3252.185 2125.515 3252.355 ;
        RECT 2076.585 3251.845 2076.755 3252.015 ;
        RECT 2028.745 3251.505 2028.915 3251.675 ;
        RECT 1690.645 2794.885 1690.815 2795.055 ;
        RECT 1060.445 2794.205 1060.615 2794.375 ;
        RECT 504.765 2793.525 504.935 2793.695 ;
        RECT 391.145 2792.845 391.315 2793.015 ;
        RECT 477.625 2792.165 477.795 2792.335 ;
        RECT 1511.245 2794.205 1511.415 2794.375 ;
        RECT 1583.465 2794.205 1583.635 2794.375 ;
        RECT 1738.485 2794.885 1738.655 2795.055 ;
        RECT 1587.145 2793.185 1587.315 2793.355 ;
        RECT 1449.145 2792.845 1449.315 2793.015 ;
        RECT 1511.245 2792.845 1511.415 2793.015 ;
        RECT 1538.845 2792.845 1539.015 2793.015 ;
        RECT 1559.545 2792.505 1559.715 2792.675 ;
        RECT 1634.985 2793.185 1635.155 2793.355 ;
        RECT 1828.185 2794.205 1828.355 2794.375 ;
        RECT 1848.885 2794.205 1849.055 2794.375 ;
        RECT 2187.445 2794.205 2187.615 2794.375 ;
        RECT 2255.985 2794.205 2256.155 2794.375 ;
        RECT 2281.285 2794.205 2281.455 2794.375 ;
        RECT 2347.985 2793.865 2348.155 2794.035 ;
        RECT 2280.825 2793.525 2280.995 2793.695 ;
        RECT 1704.445 2792.505 1704.615 2792.675 ;
        RECT 1511.245 2791.485 1511.415 2791.655 ;
        RECT 1486.865 2789.105 1487.035 2789.275 ;
        RECT 1654.765 2791.485 1654.935 2791.655 ;
        RECT 2210.905 2792.505 2211.075 2792.675 ;
        RECT 2138.685 2791.485 2138.855 2791.655 ;
        RECT 1870.045 2791.145 1870.215 2791.315 ;
        RECT 1669.945 2789.785 1670.115 2789.955 ;
        RECT 1535.165 2788.765 1535.335 2788.935 ;
        RECT 1917.425 2791.145 1917.595 2791.315 ;
        RECT 1917.885 2788.085 1918.055 2788.255 ;
        RECT 1932.145 2788.085 1932.315 2788.255 ;
        RECT 2028.285 2788.085 2028.455 2788.255 ;
        RECT 2042.545 2788.085 2042.715 2788.255 ;
        RECT 2139.145 2791.485 2139.315 2791.655 ;
        RECT 2181.465 2791.485 2181.635 2791.655 ;
        RECT 1738.945 2787.745 1739.115 2787.915 ;
        RECT 1980.445 2787.745 1980.615 2787.915 ;
        RECT 2334.185 2792.165 2334.355 2792.335 ;
        RECT 2262.885 2791.485 2263.055 2791.655 ;
        RECT 2255.985 2788.425 2256.155 2788.595 ;
        RECT 2267.485 2788.765 2267.655 2788.935 ;
        RECT 1409.125 2056.405 1409.295 2056.575 ;
      LAYER met1 ;
        RECT 1317.525 3266.960 1317.815 3267.005 ;
        RECT 1890.670 3266.960 1890.990 3267.020 ;
        RECT 1317.525 3266.820 1890.990 3266.960 ;
        RECT 1317.525 3266.775 1317.815 3266.820 ;
        RECT 1890.670 3266.760 1890.990 3266.820 ;
        RECT 1917.810 3266.960 1918.130 3267.020 ;
        RECT 2542.030 3266.960 2542.350 3267.020 ;
        RECT 1917.810 3266.820 2542.350 3266.960 ;
        RECT 1917.810 3266.760 1918.130 3266.820 ;
        RECT 2542.030 3266.760 2542.350 3266.820 ;
        RECT 1890.670 3264.580 1890.990 3264.640 ;
        RECT 1917.810 3264.580 1918.130 3264.640 ;
        RECT 1890.670 3264.440 1918.130 3264.580 ;
        RECT 1890.670 3264.380 1890.990 3264.440 ;
        RECT 1917.810 3264.380 1918.130 3264.440 ;
        RECT 2542.030 3264.240 2542.350 3264.300 ;
        RECT 2566.870 3264.240 2567.190 3264.300 ;
        RECT 2542.030 3264.100 2567.190 3264.240 ;
        RECT 2542.030 3264.040 2542.350 3264.100 ;
        RECT 2566.870 3264.040 2567.190 3264.100 ;
        RECT 646.370 3263.900 646.690 3263.960 ;
        RECT 667.990 3263.900 668.310 3263.960 ;
        RECT 676.285 3263.900 676.575 3263.945 ;
        RECT 646.370 3263.760 676.575 3263.900 ;
        RECT 646.370 3263.700 646.690 3263.760 ;
        RECT 667.990 3263.700 668.310 3263.760 ;
        RECT 676.285 3263.715 676.575 3263.760 ;
        RECT 724.125 3263.900 724.415 3263.945 ;
        RECT 772.885 3263.900 773.175 3263.945 ;
        RECT 724.125 3263.760 773.175 3263.900 ;
        RECT 724.125 3263.715 724.415 3263.760 ;
        RECT 772.885 3263.715 773.175 3263.760 ;
        RECT 820.725 3263.900 821.015 3263.945 ;
        RECT 966.085 3263.900 966.375 3263.945 ;
        RECT 820.725 3263.760 966.375 3263.900 ;
        RECT 820.725 3263.715 821.015 3263.760 ;
        RECT 966.085 3263.715 966.375 3263.760 ;
        RECT 1013.925 3263.900 1014.215 3263.945 ;
        RECT 1062.685 3263.900 1062.975 3263.945 ;
        RECT 1013.925 3263.760 1062.975 3263.900 ;
        RECT 1013.925 3263.715 1014.215 3263.760 ;
        RECT 1062.685 3263.715 1062.975 3263.760 ;
        RECT 1110.525 3263.900 1110.815 3263.945 ;
        RECT 1159.285 3263.900 1159.575 3263.945 ;
        RECT 1110.525 3263.760 1159.575 3263.900 ;
        RECT 1110.525 3263.715 1110.815 3263.760 ;
        RECT 1159.285 3263.715 1159.575 3263.760 ;
        RECT 1207.125 3263.900 1207.415 3263.945 ;
        RECT 1293.130 3263.900 1293.450 3263.960 ;
        RECT 1317.510 3263.900 1317.830 3263.960 ;
        RECT 1207.125 3263.760 1317.830 3263.900 ;
        RECT 2566.960 3263.900 2567.100 3264.040 ;
        RECT 2594.470 3263.900 2594.790 3263.960 ;
        RECT 2566.960 3263.760 2594.790 3263.900 ;
        RECT 1207.125 3263.715 1207.415 3263.760 ;
        RECT 1293.130 3263.700 1293.450 3263.760 ;
        RECT 1317.510 3263.700 1317.830 3263.760 ;
        RECT 2594.470 3263.700 2594.790 3263.760 ;
        RECT 676.285 3263.220 676.575 3263.265 ;
        RECT 696.970 3263.220 697.290 3263.280 ;
        RECT 724.125 3263.220 724.415 3263.265 ;
        RECT 676.285 3263.080 724.415 3263.220 ;
        RECT 676.285 3263.035 676.575 3263.080 ;
        RECT 696.970 3263.020 697.290 3263.080 ;
        RECT 724.125 3263.035 724.415 3263.080 ;
        RECT 772.885 3263.220 773.175 3263.265 ;
        RECT 820.725 3263.220 821.015 3263.265 ;
        RECT 772.885 3263.080 821.015 3263.220 ;
        RECT 772.885 3263.035 773.175 3263.080 ;
        RECT 820.725 3263.035 821.015 3263.080 ;
        RECT 966.085 3263.220 966.375 3263.265 ;
        RECT 1013.925 3263.220 1014.215 3263.265 ;
        RECT 966.085 3263.080 1014.215 3263.220 ;
        RECT 966.085 3263.035 966.375 3263.080 ;
        RECT 1013.925 3263.035 1014.215 3263.080 ;
        RECT 1062.685 3263.220 1062.975 3263.265 ;
        RECT 1110.525 3263.220 1110.815 3263.265 ;
        RECT 1062.685 3263.080 1110.815 3263.220 ;
        RECT 1062.685 3263.035 1062.975 3263.080 ;
        RECT 1110.525 3263.035 1110.815 3263.080 ;
        RECT 1159.285 3263.220 1159.575 3263.265 ;
        RECT 1207.125 3263.220 1207.415 3263.265 ;
        RECT 1159.285 3263.080 1207.415 3263.220 ;
        RECT 1159.285 3263.035 1159.575 3263.080 ;
        RECT 1207.125 3263.035 1207.415 3263.080 ;
        RECT 1593.985 3254.040 1594.275 3254.085 ;
        RECT 1641.825 3254.040 1642.115 3254.085 ;
        RECT 1593.985 3253.900 1642.115 3254.040 ;
        RECT 1593.985 3253.855 1594.275 3253.900 ;
        RECT 1641.825 3253.855 1642.115 3253.900 ;
        RECT 1690.585 3254.040 1690.875 3254.085 ;
        RECT 1738.425 3254.040 1738.715 3254.085 ;
        RECT 1690.585 3253.900 1738.715 3254.040 ;
        RECT 1690.585 3253.855 1690.875 3253.900 ;
        RECT 1738.425 3253.855 1738.715 3253.900 ;
        RECT 1787.185 3254.040 1787.475 3254.085 ;
        RECT 1835.025 3254.040 1835.315 3254.085 ;
        RECT 1787.185 3253.900 1835.315 3254.040 ;
        RECT 1787.185 3253.855 1787.475 3253.900 ;
        RECT 1835.025 3253.855 1835.315 3253.900 ;
        RECT 2270.185 3254.040 2270.475 3254.085 ;
        RECT 2318.025 3254.040 2318.315 3254.085 ;
        RECT 2270.185 3253.900 2318.315 3254.040 ;
        RECT 2270.185 3253.855 2270.475 3253.900 ;
        RECT 2318.025 3253.855 2318.315 3253.900 ;
        RECT 2366.785 3254.040 2367.075 3254.085 ;
        RECT 2414.625 3254.040 2414.915 3254.085 ;
        RECT 2366.785 3253.900 2414.915 3254.040 ;
        RECT 2366.785 3253.855 2367.075 3253.900 ;
        RECT 2414.625 3253.855 2414.915 3253.900 ;
        RECT 2463.385 3254.040 2463.675 3254.085 ;
        RECT 2511.225 3254.040 2511.515 3254.085 ;
        RECT 2463.385 3253.900 2511.515 3254.040 ;
        RECT 2463.385 3253.855 2463.675 3253.900 ;
        RECT 2511.225 3253.855 2511.515 3253.900 ;
        RECT 1014.385 3253.700 1014.675 3253.745 ;
        RECT 1055.785 3253.700 1056.075 3253.745 ;
        RECT 1014.385 3253.560 1056.075 3253.700 ;
        RECT 1014.385 3253.515 1014.675 3253.560 ;
        RECT 1055.785 3253.515 1056.075 3253.560 ;
        RECT 1110.985 3253.700 1111.275 3253.745 ;
        RECT 1152.385 3253.700 1152.675 3253.745 ;
        RECT 1110.985 3253.560 1152.675 3253.700 ;
        RECT 1110.985 3253.515 1111.275 3253.560 ;
        RECT 1152.385 3253.515 1152.675 3253.560 ;
        RECT 1207.585 3253.360 1207.875 3253.405 ;
        RECT 1231.505 3253.360 1231.795 3253.405 ;
        RECT 1593.985 3253.360 1594.275 3253.405 ;
        RECT 1690.585 3253.360 1690.875 3253.405 ;
        RECT 1787.185 3253.360 1787.475 3253.405 ;
        RECT 2270.185 3253.360 2270.475 3253.405 ;
        RECT 2366.785 3253.360 2367.075 3253.405 ;
        RECT 2463.385 3253.360 2463.675 3253.405 ;
        RECT 1207.585 3253.220 1231.795 3253.360 ;
        RECT 1207.585 3253.175 1207.875 3253.220 ;
        RECT 1231.505 3253.175 1231.795 3253.220 ;
        RECT 1565.540 3253.220 1594.275 3253.360 ;
        RECT 1007.100 3252.880 1014.140 3253.020 ;
        RECT 883.285 3252.680 883.575 3252.725 ;
        RECT 917.785 3252.680 918.075 3252.725 ;
        RECT 883.285 3252.540 918.075 3252.680 ;
        RECT 883.285 3252.495 883.575 3252.540 ;
        RECT 917.785 3252.495 918.075 3252.540 ;
        RECT 959.185 3252.680 959.475 3252.725 ;
        RECT 1007.100 3252.680 1007.240 3252.880 ;
        RECT 959.185 3252.540 1007.240 3252.680 ;
        RECT 1014.000 3252.680 1014.140 3252.880 ;
        RECT 1014.385 3252.835 1014.675 3253.065 ;
        RECT 1103.625 3253.020 1103.915 3253.065 ;
        RECT 1103.625 3252.880 1110.740 3253.020 ;
        RECT 1103.625 3252.835 1103.915 3252.880 ;
        RECT 1014.460 3252.680 1014.600 3252.835 ;
        RECT 1014.000 3252.540 1014.600 3252.680 ;
        RECT 1110.600 3252.680 1110.740 3252.880 ;
        RECT 1110.985 3252.835 1111.275 3253.065 ;
        RECT 1200.225 3253.020 1200.515 3253.065 ;
        RECT 1559.025 3253.020 1559.315 3253.065 ;
        RECT 1200.225 3252.880 1207.340 3253.020 ;
        RECT 1200.225 3252.835 1200.515 3252.880 ;
        RECT 1111.060 3252.680 1111.200 3252.835 ;
        RECT 1110.600 3252.540 1111.200 3252.680 ;
        RECT 1207.200 3252.680 1207.340 3252.880 ;
        RECT 1510.800 3252.880 1559.315 3253.020 ;
        RECT 1297.285 3252.680 1297.575 3252.725 ;
        RECT 1332.230 3252.680 1332.550 3252.740 ;
        RECT 1207.200 3252.540 1207.800 3252.680 ;
        RECT 959.185 3252.495 959.475 3252.540 ;
        RECT 1207.660 3252.385 1207.800 3252.540 ;
        RECT 1297.285 3252.540 1332.550 3252.680 ;
        RECT 1297.285 3252.495 1297.575 3252.540 ;
        RECT 1332.230 3252.480 1332.550 3252.540 ;
        RECT 1496.925 3252.680 1497.215 3252.725 ;
        RECT 1510.800 3252.680 1510.940 3252.880 ;
        RECT 1559.025 3252.835 1559.315 3252.880 ;
        RECT 1559.485 3253.020 1559.775 3253.065 ;
        RECT 1565.540 3253.020 1565.680 3253.220 ;
        RECT 1593.985 3253.175 1594.275 3253.220 ;
        RECT 1662.140 3253.220 1690.875 3253.360 ;
        RECT 1559.485 3252.880 1565.680 3253.020 ;
        RECT 1641.825 3253.020 1642.115 3253.065 ;
        RECT 1655.625 3253.020 1655.915 3253.065 ;
        RECT 1641.825 3252.880 1655.915 3253.020 ;
        RECT 1559.485 3252.835 1559.775 3252.880 ;
        RECT 1641.825 3252.835 1642.115 3252.880 ;
        RECT 1655.625 3252.835 1655.915 3252.880 ;
        RECT 1656.085 3253.020 1656.375 3253.065 ;
        RECT 1662.140 3253.020 1662.280 3253.220 ;
        RECT 1690.585 3253.175 1690.875 3253.220 ;
        RECT 1758.740 3253.220 1787.475 3253.360 ;
        RECT 1656.085 3252.880 1662.280 3253.020 ;
        RECT 1738.425 3253.020 1738.715 3253.065 ;
        RECT 1752.225 3253.020 1752.515 3253.065 ;
        RECT 1738.425 3252.880 1752.515 3253.020 ;
        RECT 1656.085 3252.835 1656.375 3252.880 ;
        RECT 1738.425 3252.835 1738.715 3252.880 ;
        RECT 1752.225 3252.835 1752.515 3252.880 ;
        RECT 1752.685 3253.020 1752.975 3253.065 ;
        RECT 1758.740 3253.020 1758.880 3253.220 ;
        RECT 1787.185 3253.175 1787.475 3253.220 ;
        RECT 2241.740 3253.220 2270.475 3253.360 ;
        RECT 1752.685 3252.880 1758.880 3253.020 ;
        RECT 1835.025 3253.020 1835.315 3253.065 ;
        RECT 1849.285 3253.020 1849.575 3253.065 ;
        RECT 1835.025 3252.880 1849.575 3253.020 ;
        RECT 1752.685 3252.835 1752.975 3252.880 ;
        RECT 1835.025 3252.835 1835.315 3252.880 ;
        RECT 1849.285 3252.835 1849.575 3252.880 ;
        RECT 1849.745 3253.020 1850.035 3253.065 ;
        RECT 2235.225 3253.020 2235.515 3253.065 ;
        RECT 1849.745 3252.880 1883.540 3253.020 ;
        RECT 1849.745 3252.835 1850.035 3252.880 ;
        RECT 1496.925 3252.540 1510.940 3252.680 ;
        RECT 1883.400 3252.680 1883.540 3252.880 ;
        RECT 2187.000 3252.880 2235.515 3253.020 ;
        RECT 1948.185 3252.680 1948.475 3252.725 ;
        RECT 1980.385 3252.680 1980.675 3252.725 ;
        RECT 1883.400 3252.540 1897.340 3252.680 ;
        RECT 1496.925 3252.495 1497.215 3252.540 ;
        RECT 724.200 3252.200 724.800 3252.340 ;
        RECT 688.230 3252.000 688.550 3252.060 ;
        RECT 724.200 3252.000 724.340 3252.200 ;
        RECT 724.660 3252.045 724.800 3252.200 ;
        RECT 772.885 3252.155 773.175 3252.385 ;
        RECT 1055.785 3252.340 1056.075 3252.385 ;
        RECT 1103.625 3252.340 1103.915 3252.385 ;
        RECT 1055.785 3252.200 1103.915 3252.340 ;
        RECT 1055.785 3252.155 1056.075 3252.200 ;
        RECT 1103.625 3252.155 1103.915 3252.200 ;
        RECT 1152.385 3252.340 1152.675 3252.385 ;
        RECT 1200.225 3252.340 1200.515 3252.385 ;
        RECT 1152.385 3252.200 1200.515 3252.340 ;
        RECT 1152.385 3252.155 1152.675 3252.200 ;
        RECT 1200.225 3252.155 1200.515 3252.200 ;
        RECT 1207.585 3252.155 1207.875 3252.385 ;
        RECT 1231.505 3252.340 1231.795 3252.385 ;
        RECT 1269.225 3252.340 1269.515 3252.385 ;
        RECT 1231.505 3252.200 1269.515 3252.340 ;
        RECT 1231.505 3252.155 1231.795 3252.200 ;
        RECT 1269.225 3252.155 1269.515 3252.200 ;
        RECT 1414.110 3252.340 1414.430 3252.400 ;
        RECT 1449.085 3252.340 1449.375 3252.385 ;
        RECT 1414.110 3252.200 1449.375 3252.340 ;
        RECT 1897.200 3252.340 1897.340 3252.540 ;
        RECT 1948.185 3252.540 1980.675 3252.680 ;
        RECT 1948.185 3252.495 1948.475 3252.540 ;
        RECT 1980.385 3252.495 1980.675 3252.540 ;
        RECT 2173.125 3252.680 2173.415 3252.725 ;
        RECT 2187.000 3252.680 2187.140 3252.880 ;
        RECT 2235.225 3252.835 2235.515 3252.880 ;
        RECT 2235.685 3253.020 2235.975 3253.065 ;
        RECT 2241.740 3253.020 2241.880 3253.220 ;
        RECT 2270.185 3253.175 2270.475 3253.220 ;
        RECT 2338.340 3253.220 2367.075 3253.360 ;
        RECT 2235.685 3252.880 2241.880 3253.020 ;
        RECT 2318.025 3253.020 2318.315 3253.065 ;
        RECT 2331.825 3253.020 2332.115 3253.065 ;
        RECT 2318.025 3252.880 2332.115 3253.020 ;
        RECT 2235.685 3252.835 2235.975 3252.880 ;
        RECT 2318.025 3252.835 2318.315 3252.880 ;
        RECT 2331.825 3252.835 2332.115 3252.880 ;
        RECT 2332.285 3253.020 2332.575 3253.065 ;
        RECT 2338.340 3253.020 2338.480 3253.220 ;
        RECT 2366.785 3253.175 2367.075 3253.220 ;
        RECT 2434.940 3253.220 2463.675 3253.360 ;
        RECT 2332.285 3252.880 2338.480 3253.020 ;
        RECT 2414.625 3253.020 2414.915 3253.065 ;
        RECT 2428.425 3253.020 2428.715 3253.065 ;
        RECT 2414.625 3252.880 2428.715 3253.020 ;
        RECT 2332.285 3252.835 2332.575 3252.880 ;
        RECT 2414.625 3252.835 2414.915 3252.880 ;
        RECT 2428.425 3252.835 2428.715 3252.880 ;
        RECT 2428.885 3253.020 2429.175 3253.065 ;
        RECT 2434.940 3253.020 2435.080 3253.220 ;
        RECT 2463.385 3253.175 2463.675 3253.220 ;
        RECT 2428.885 3252.880 2435.080 3253.020 ;
        RECT 2511.225 3253.020 2511.515 3253.065 ;
        RECT 2525.485 3253.020 2525.775 3253.065 ;
        RECT 2511.225 3252.880 2525.775 3253.020 ;
        RECT 2428.885 3252.835 2429.175 3252.880 ;
        RECT 2511.225 3252.835 2511.515 3252.880 ;
        RECT 2525.485 3252.835 2525.775 3252.880 ;
        RECT 2525.945 3253.020 2526.235 3253.065 ;
        RECT 2525.945 3252.880 2559.740 3253.020 ;
        RECT 2525.945 3252.835 2526.235 3252.880 ;
        RECT 2173.125 3252.540 2187.140 3252.680 ;
        RECT 2559.600 3252.680 2559.740 3252.880 ;
        RECT 2559.600 3252.540 2573.540 3252.680 ;
        RECT 2173.125 3252.495 2173.415 3252.540 ;
        RECT 1932.085 3252.340 1932.375 3252.385 ;
        RECT 2125.285 3252.340 2125.575 3252.385 ;
        RECT 1897.200 3252.200 1932.375 3252.340 ;
        RECT 688.230 3251.860 724.340 3252.000 ;
        RECT 688.230 3251.800 688.550 3251.860 ;
        RECT 724.585 3251.815 724.875 3252.045 ;
        RECT 748.505 3252.000 748.795 3252.045 ;
        RECT 772.960 3252.000 773.100 3252.155 ;
        RECT 1414.110 3252.140 1414.430 3252.200 ;
        RECT 1449.085 3252.155 1449.375 3252.200 ;
        RECT 1932.085 3252.155 1932.375 3252.200 ;
        RECT 2090.400 3252.200 2125.575 3252.340 ;
        RECT 2573.400 3252.340 2573.540 3252.540 ;
        RECT 2582.050 3252.340 2582.370 3252.400 ;
        RECT 2573.400 3252.200 2582.370 3252.340 ;
        RECT 748.505 3251.860 773.100 3252.000 ;
        RECT 869.010 3252.000 869.330 3252.060 ;
        RECT 883.285 3252.000 883.575 3252.045 ;
        RECT 869.010 3251.860 883.575 3252.000 ;
        RECT 748.505 3251.815 748.795 3251.860 ;
        RECT 869.010 3251.800 869.330 3251.860 ;
        RECT 883.285 3251.815 883.575 3251.860 ;
        RECT 917.785 3252.000 918.075 3252.045 ;
        RECT 959.185 3252.000 959.475 3252.045 ;
        RECT 917.785 3251.860 959.475 3252.000 ;
        RECT 917.785 3251.815 918.075 3251.860 ;
        RECT 959.185 3251.815 959.475 3251.860 ;
        RECT 1297.285 3251.815 1297.575 3252.045 ;
        RECT 1352.485 3252.000 1352.775 3252.045 ;
        RECT 1400.325 3252.000 1400.615 3252.045 ;
        RECT 1352.485 3251.860 1400.615 3252.000 ;
        RECT 1352.485 3251.815 1352.775 3251.860 ;
        RECT 1400.325 3251.815 1400.615 3251.860 ;
        RECT 2076.525 3252.000 2076.815 3252.045 ;
        RECT 2090.400 3252.000 2090.540 3252.200 ;
        RECT 2125.285 3252.155 2125.575 3252.200 ;
        RECT 2582.050 3252.140 2582.370 3252.200 ;
        RECT 2076.525 3251.860 2090.540 3252.000 ;
        RECT 2076.525 3251.815 2076.815 3251.860 ;
        RECT 1270.145 3251.660 1270.435 3251.705 ;
        RECT 1297.360 3251.660 1297.500 3251.815 ;
        RECT 820.800 3251.520 821.400 3251.660 ;
        RECT 772.885 3251.320 773.175 3251.365 ;
        RECT 820.800 3251.320 820.940 3251.520 ;
        RECT 821.260 3251.380 821.400 3251.520 ;
        RECT 1270.145 3251.520 1297.500 3251.660 ;
        RECT 1449.085 3251.660 1449.375 3251.705 ;
        RECT 1496.925 3251.660 1497.215 3251.705 ;
        RECT 1449.085 3251.520 1497.215 3251.660 ;
        RECT 1270.145 3251.475 1270.435 3251.520 ;
        RECT 1449.085 3251.475 1449.375 3251.520 ;
        RECT 1496.925 3251.475 1497.215 3251.520 ;
        RECT 1980.385 3251.660 1980.675 3251.705 ;
        RECT 2028.685 3251.660 2028.975 3251.705 ;
        RECT 1980.385 3251.520 2028.975 3251.660 ;
        RECT 1980.385 3251.475 1980.675 3251.520 ;
        RECT 2028.685 3251.475 2028.975 3251.520 ;
        RECT 2125.285 3251.660 2125.575 3251.705 ;
        RECT 2173.125 3251.660 2173.415 3251.705 ;
        RECT 2125.285 3251.520 2173.415 3251.660 ;
        RECT 2125.285 3251.475 2125.575 3251.520 ;
        RECT 2173.125 3251.475 2173.415 3251.520 ;
      LAYER met1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met1 ;
        RECT 772.885 3251.180 820.940 3251.320 ;
        RECT 772.885 3251.135 773.175 3251.180 ;
        RECT 821.170 3251.120 821.490 3251.380 ;
        RECT 1332.230 3251.320 1332.550 3251.380 ;
        RECT 1352.485 3251.320 1352.775 3251.365 ;
        RECT 724.585 3250.980 724.875 3251.025 ;
        RECT 748.505 3250.980 748.795 3251.025 ;
        RECT 724.585 3250.840 748.795 3250.980 ;
        RECT 724.585 3250.795 724.875 3250.840 ;
        RECT 748.505 3250.795 748.795 3250.840 ;
        RECT 927.890 2898.400 928.210 2898.460 ;
        RECT 939.390 2898.400 939.710 2898.460 ;
        RECT 927.890 2898.260 939.710 2898.400 ;
        RECT 927.890 2898.200 928.210 2898.260 ;
        RECT 939.390 2898.200 939.710 2898.260 ;
      LAYER met1 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met1 ;
        RECT 1332.230 3251.180 1352.775 3251.320 ;
        RECT 1932.085 3251.320 1932.375 3251.365 ;
        RECT 1935.750 3251.320 1936.070 3251.380 ;
        RECT 1948.185 3251.320 1948.475 3251.365 ;
        RECT 1332.230 3251.120 1332.550 3251.180 ;
        RECT 1352.485 3251.135 1352.775 3251.180 ;
        RECT 1400.325 3250.980 1400.615 3251.025 ;
        RECT 1407.670 3250.980 1407.990 3251.040 ;
        RECT 1414.110 3250.980 1414.430 3251.040 ;
        RECT 1400.325 3250.840 1414.430 3250.980 ;
        RECT 1400.325 3250.795 1400.615 3250.840 ;
        RECT 1407.670 3250.780 1407.990 3250.840 ;
        RECT 1414.110 3250.780 1414.430 3250.840 ;
        RECT 1472.990 3229.560 1473.310 3229.620 ;
        RECT 1536.930 3229.560 1537.250 3229.620 ;
        RECT 1472.990 3229.420 1537.250 3229.560 ;
        RECT 1472.990 3229.360 1473.310 3229.420 ;
        RECT 1536.930 3229.360 1537.250 3229.420 ;
        RECT 1459.190 3222.420 1459.510 3222.480 ;
        RECT 1535.550 3222.420 1535.870 3222.480 ;
        RECT 1459.190 3222.280 1535.870 3222.420 ;
        RECT 1459.190 3222.220 1459.510 3222.280 ;
        RECT 1535.550 3222.220 1535.870 3222.280 ;
        RECT 1452.290 3215.620 1452.610 3215.680 ;
        RECT 1535.550 3215.620 1535.870 3215.680 ;
        RECT 1452.290 3215.480 1535.870 3215.620 ;
        RECT 1452.290 3215.420 1452.610 3215.480 ;
        RECT 1535.550 3215.420 1535.870 3215.480 ;
        RECT 1438.490 3208.820 1438.810 3208.880 ;
        RECT 1538.310 3208.820 1538.630 3208.880 ;
        RECT 1438.490 3208.680 1538.630 3208.820 ;
        RECT 1438.490 3208.620 1438.810 3208.680 ;
        RECT 1538.310 3208.620 1538.630 3208.680 ;
        RECT 1431.590 3201.680 1431.910 3201.740 ;
        RECT 1538.310 3201.680 1538.630 3201.740 ;
        RECT 1431.590 3201.540 1538.630 3201.680 ;
        RECT 1431.590 3201.480 1431.910 3201.540 ;
        RECT 1538.310 3201.480 1538.630 3201.540 ;
        RECT 1424.690 3194.880 1425.010 3194.940 ;
        RECT 1533.250 3194.880 1533.570 3194.940 ;
        RECT 1424.690 3194.740 1533.570 3194.880 ;
        RECT 1424.690 3194.680 1425.010 3194.740 ;
        RECT 1533.250 3194.680 1533.570 3194.740 ;
        RECT 1473.450 3188.080 1473.770 3188.140 ;
        RECT 1534.170 3188.080 1534.490 3188.140 ;
        RECT 1473.450 3187.940 1534.490 3188.080 ;
        RECT 1473.450 3187.880 1473.770 3187.940 ;
        RECT 1534.170 3187.880 1534.490 3187.940 ;
        RECT 1352.010 2901.460 1352.330 2901.520 ;
        RECT 1397.550 2901.460 1397.870 2901.520 ;
        RECT 1352.010 2901.320 1397.870 2901.460 ;
        RECT 1352.010 2901.260 1352.330 2901.320 ;
        RECT 1397.550 2901.260 1397.870 2901.320 ;
        RECT 1459.650 2898.400 1459.970 2898.460 ;
        RECT 1538.310 2898.400 1538.630 2898.460 ;
        RECT 1459.650 2898.260 1538.630 2898.400 ;
        RECT 1459.650 2898.200 1459.970 2898.260 ;
        RECT 1538.310 2898.200 1538.630 2898.260 ;
      LAYER met1 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met1 ;
        RECT 1932.085 3251.180 1948.475 3251.320 ;
        RECT 1932.085 3251.135 1932.375 3251.180 ;
        RECT 1935.750 3251.120 1936.070 3251.180 ;
        RECT 1948.185 3251.135 1948.475 3251.180 ;
        RECT 2028.685 3250.980 2028.975 3251.025 ;
        RECT 2076.525 3250.980 2076.815 3251.025 ;
        RECT 2028.685 3250.840 2076.815 3250.980 ;
        RECT 2028.685 3250.795 2028.975 3250.840 ;
        RECT 2076.525 3250.795 2076.815 3250.840 ;
      LAYER met1 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met1 ;
        RECT 1690.585 2795.040 1690.875 2795.085 ;
        RECT 1732.890 2795.040 1733.210 2795.100 ;
        RECT 1738.425 2795.040 1738.715 2795.085 ;
        RECT 1690.585 2794.900 1738.715 2795.040 ;
        RECT 1690.585 2794.855 1690.875 2794.900 ;
        RECT 1732.890 2794.840 1733.210 2794.900 ;
        RECT 1738.425 2794.855 1738.715 2794.900 ;
        RECT 2279.920 2794.560 2280.980 2794.700 ;
        RECT 386.930 2794.360 387.250 2794.420 ;
        RECT 432.010 2794.360 432.330 2794.420 ;
        RECT 433.390 2794.360 433.710 2794.420 ;
        RECT 386.930 2794.220 433.710 2794.360 ;
        RECT 386.930 2794.160 387.250 2794.220 ;
        RECT 432.010 2794.160 432.330 2794.220 ;
        RECT 433.390 2794.160 433.710 2794.220 ;
        RECT 482.610 2794.360 482.930 2794.420 ;
        RECT 500.550 2794.360 500.870 2794.420 ;
        RECT 482.610 2794.220 500.870 2794.360 ;
        RECT 482.610 2794.160 482.930 2794.220 ;
        RECT 500.550 2794.160 500.870 2794.220 ;
        RECT 648.210 2794.360 648.530 2794.420 ;
        RECT 1053.010 2794.360 1053.330 2794.420 ;
        RECT 1060.385 2794.360 1060.675 2794.405 ;
        RECT 648.210 2794.220 1060.675 2794.360 ;
        RECT 648.210 2794.160 648.530 2794.220 ;
        RECT 1053.010 2794.160 1053.330 2794.220 ;
        RECT 1060.385 2794.175 1060.675 2794.220 ;
        RECT 1418.710 2794.360 1419.030 2794.420 ;
        RECT 1511.185 2794.360 1511.475 2794.405 ;
        RECT 1418.710 2794.220 1511.475 2794.360 ;
        RECT 1418.710 2794.160 1419.030 2794.220 ;
        RECT 1511.185 2794.175 1511.475 2794.220 ;
        RECT 1583.405 2794.360 1583.695 2794.405 ;
        RECT 1828.125 2794.360 1828.415 2794.405 ;
        RECT 1583.405 2794.220 1828.415 2794.360 ;
        RECT 1583.405 2794.175 1583.695 2794.220 ;
        RECT 1828.125 2794.175 1828.415 2794.220 ;
        RECT 1848.825 2794.360 1849.115 2794.405 ;
        RECT 2187.385 2794.360 2187.675 2794.405 ;
        RECT 1848.825 2794.220 2187.675 2794.360 ;
        RECT 1848.825 2794.175 1849.115 2794.220 ;
        RECT 2187.385 2794.175 2187.675 2794.220 ;
        RECT 2255.925 2794.360 2256.215 2794.405 ;
        RECT 2279.920 2794.360 2280.060 2794.560 ;
        RECT 2255.925 2794.220 2280.060 2794.360 ;
        RECT 2255.925 2794.175 2256.215 2794.220 ;
        RECT 462.370 2794.020 462.690 2794.080 ;
        RECT 503.770 2794.020 504.090 2794.080 ;
        RECT 513.890 2794.020 514.210 2794.080 ;
        RECT 676.270 2794.020 676.590 2794.080 ;
        RECT 462.370 2793.880 504.090 2794.020 ;
        RECT 462.370 2793.820 462.690 2793.880 ;
        RECT 503.770 2793.820 504.090 2793.880 ;
        RECT 504.320 2793.880 676.590 2794.020 ;
        RECT 374.970 2793.680 375.290 2793.740 ;
        RECT 420.970 2793.680 421.290 2793.740 ;
        RECT 466.510 2793.680 466.830 2793.740 ;
        RECT 504.320 2793.680 504.460 2793.880 ;
        RECT 513.890 2793.820 514.210 2793.880 ;
        RECT 676.270 2793.820 676.590 2793.880 ;
        RECT 1419.170 2794.020 1419.490 2794.080 ;
        RECT 2280.840 2794.020 2280.980 2794.560 ;
        RECT 2281.225 2794.360 2281.515 2794.405 ;
        RECT 2415.070 2794.360 2415.390 2794.420 ;
        RECT 2281.225 2794.220 2415.390 2794.360 ;
        RECT 2281.225 2794.175 2281.515 2794.220 ;
        RECT 2415.070 2794.160 2415.390 2794.220 ;
        RECT 2284.430 2794.020 2284.750 2794.080 ;
        RECT 1419.170 2793.880 2280.060 2794.020 ;
        RECT 2280.840 2793.880 2284.750 2794.020 ;
        RECT 1419.170 2793.820 1419.490 2793.880 ;
        RECT 374.970 2793.540 504.460 2793.680 ;
        RECT 504.705 2793.680 504.995 2793.725 ;
        RECT 526.770 2793.680 527.090 2793.740 ;
        RECT 696.970 2793.680 697.290 2793.740 ;
        RECT 504.705 2793.540 697.290 2793.680 ;
        RECT 374.970 2793.480 375.290 2793.540 ;
        RECT 420.970 2793.480 421.290 2793.540 ;
        RECT 466.510 2793.480 466.830 2793.540 ;
        RECT 504.705 2793.495 504.995 2793.540 ;
        RECT 526.770 2793.480 527.090 2793.540 ;
        RECT 696.970 2793.480 697.290 2793.540 ;
        RECT 700.190 2793.680 700.510 2793.740 ;
        RECT 1001.030 2793.680 1001.350 2793.740 ;
        RECT 700.190 2793.540 1001.350 2793.680 ;
        RECT 700.190 2793.480 700.510 2793.540 ;
        RECT 1001.030 2793.480 1001.350 2793.540 ;
        RECT 1090.270 2793.680 1090.590 2793.740 ;
        RECT 1094.410 2793.680 1094.730 2793.740 ;
        RECT 1139.950 2793.680 1140.270 2793.740 ;
        RECT 1186.870 2793.680 1187.190 2793.740 ;
        RECT 1090.270 2793.540 1187.190 2793.680 ;
        RECT 1090.270 2793.480 1090.590 2793.540 ;
        RECT 1094.410 2793.480 1094.730 2793.540 ;
        RECT 1139.950 2793.480 1140.270 2793.540 ;
        RECT 1186.870 2793.480 1187.190 2793.540 ;
        RECT 1511.185 2793.680 1511.475 2793.725 ;
        RECT 1583.405 2793.680 1583.695 2793.725 ;
        RECT 1511.185 2793.540 1583.695 2793.680 ;
        RECT 1511.185 2793.495 1511.475 2793.540 ;
        RECT 1583.405 2793.495 1583.695 2793.540 ;
        RECT 1642.730 2793.680 1643.050 2793.740 ;
        RECT 1687.810 2793.680 1688.130 2793.740 ;
        RECT 1642.730 2793.540 1688.130 2793.680 ;
        RECT 1642.730 2793.480 1643.050 2793.540 ;
        RECT 1687.810 2793.480 1688.130 2793.540 ;
        RECT 1689.190 2793.680 1689.510 2793.740 ;
        RECT 1690.585 2793.680 1690.875 2793.725 ;
        RECT 1689.190 2793.540 1690.875 2793.680 ;
        RECT 1689.190 2793.480 1689.510 2793.540 ;
        RECT 1690.585 2793.495 1690.875 2793.540 ;
        RECT 1723.690 2793.680 1724.010 2793.740 ;
        RECT 1766.470 2793.680 1766.790 2793.740 ;
        RECT 1723.690 2793.540 1766.790 2793.680 ;
        RECT 1723.690 2793.480 1724.010 2793.540 ;
        RECT 1766.470 2793.480 1766.790 2793.540 ;
        RECT 2245.790 2793.680 2246.110 2793.740 ;
        RECT 2279.385 2793.680 2279.675 2793.725 ;
        RECT 2245.790 2793.540 2279.675 2793.680 ;
        RECT 2245.790 2793.480 2246.110 2793.540 ;
        RECT 2279.385 2793.495 2279.675 2793.540 ;
        RECT 380.030 2793.340 380.350 2793.400 ;
        RECT 426.950 2793.340 427.270 2793.400 ;
        RECT 475.250 2793.340 475.570 2793.400 ;
        RECT 380.030 2793.200 475.570 2793.340 ;
        RECT 380.030 2793.140 380.350 2793.200 ;
        RECT 426.950 2793.140 427.270 2793.200 ;
        RECT 475.250 2793.140 475.570 2793.200 ;
        RECT 503.770 2793.340 504.090 2793.400 ;
        RECT 508.830 2793.340 509.150 2793.400 ;
        RECT 662.470 2793.340 662.790 2793.400 ;
        RECT 503.770 2793.200 662.790 2793.340 ;
        RECT 503.770 2793.140 504.090 2793.200 ;
        RECT 508.830 2793.140 509.150 2793.200 ;
        RECT 662.470 2793.140 662.790 2793.200 ;
        RECT 686.390 2793.340 686.710 2793.400 ;
        RECT 986.770 2793.340 987.090 2793.400 ;
        RECT 686.390 2793.200 987.090 2793.340 ;
        RECT 686.390 2793.140 686.710 2793.200 ;
        RECT 986.770 2793.140 987.090 2793.200 ;
        RECT 1083.370 2793.340 1083.690 2793.400 ;
        RECT 1129.370 2793.340 1129.690 2793.400 ;
        RECT 1173.070 2793.340 1173.390 2793.400 ;
        RECT 1083.370 2793.200 1173.390 2793.340 ;
        RECT 1083.370 2793.140 1083.690 2793.200 ;
        RECT 1129.370 2793.140 1129.690 2793.200 ;
        RECT 1173.070 2793.140 1173.390 2793.200 ;
        RECT 1587.085 2793.340 1587.375 2793.385 ;
        RECT 1634.925 2793.340 1635.215 2793.385 ;
        RECT 1587.085 2793.200 1635.215 2793.340 ;
        RECT 1587.085 2793.155 1587.375 2793.200 ;
        RECT 1634.925 2793.155 1635.215 2793.200 ;
        RECT 1738.425 2793.340 1738.715 2793.385 ;
        RECT 1780.270 2793.340 1780.590 2793.400 ;
        RECT 1738.425 2793.200 1780.590 2793.340 ;
        RECT 1738.425 2793.155 1738.715 2793.200 ;
        RECT 1780.270 2793.140 1780.590 2793.200 ;
        RECT 1828.125 2793.340 1828.415 2793.385 ;
        RECT 1848.825 2793.340 1849.115 2793.385 ;
        RECT 1828.125 2793.200 1849.115 2793.340 ;
        RECT 1828.125 2793.155 1828.415 2793.200 ;
        RECT 1848.825 2793.155 1849.115 2793.200 ;
        RECT 2187.385 2793.340 2187.675 2793.385 ;
        RECT 2255.925 2793.340 2256.215 2793.385 ;
        RECT 2187.385 2793.200 2256.215 2793.340 ;
        RECT 2279.920 2793.340 2280.060 2793.880 ;
        RECT 2284.430 2793.820 2284.750 2793.880 ;
        RECT 2300.990 2794.020 2301.310 2794.080 ;
        RECT 2304.210 2794.020 2304.530 2794.080 ;
        RECT 2347.450 2794.020 2347.770 2794.080 ;
        RECT 2300.990 2793.880 2347.770 2794.020 ;
        RECT 2300.990 2793.820 2301.310 2793.880 ;
        RECT 2304.210 2793.820 2304.530 2793.880 ;
        RECT 2347.450 2793.820 2347.770 2793.880 ;
        RECT 2347.925 2794.020 2348.215 2794.065 ;
        RECT 2385.630 2794.020 2385.950 2794.080 ;
        RECT 2428.870 2794.020 2429.190 2794.080 ;
        RECT 2347.925 2793.880 2429.190 2794.020 ;
        RECT 2347.925 2793.835 2348.215 2793.880 ;
        RECT 2385.630 2793.820 2385.950 2793.880 ;
        RECT 2428.870 2793.820 2429.190 2793.880 ;
        RECT 2280.765 2793.680 2281.055 2793.725 ;
        RECT 2308.810 2793.680 2309.130 2793.740 ;
        RECT 2356.650 2793.680 2356.970 2793.740 ;
        RECT 2402.650 2793.680 2402.970 2793.740 ;
        RECT 2280.765 2793.540 2402.970 2793.680 ;
        RECT 2280.765 2793.495 2281.055 2793.540 ;
        RECT 2308.810 2793.480 2309.130 2793.540 ;
        RECT 2356.650 2793.480 2356.970 2793.540 ;
        RECT 2402.650 2793.480 2402.970 2793.540 ;
        RECT 2298.230 2793.340 2298.550 2793.400 ;
        RECT 2343.770 2793.340 2344.090 2793.400 ;
        RECT 2391.610 2793.340 2391.930 2793.400 ;
        RECT 2435.770 2793.340 2436.090 2793.400 ;
        RECT 2279.920 2793.200 2436.090 2793.340 ;
        RECT 2187.385 2793.155 2187.675 2793.200 ;
        RECT 2255.925 2793.155 2256.215 2793.200 ;
        RECT 2298.230 2793.140 2298.550 2793.200 ;
        RECT 2343.770 2793.140 2344.090 2793.200 ;
        RECT 2391.610 2793.140 2391.930 2793.200 ;
        RECT 2435.770 2793.140 2436.090 2793.200 ;
        RECT 391.085 2793.000 391.375 2793.045 ;
        RECT 409.930 2793.000 410.250 2793.060 ;
        RECT 455.470 2793.000 455.790 2793.060 ;
        RECT 391.085 2792.860 455.790 2793.000 ;
        RECT 391.085 2792.815 391.375 2792.860 ;
        RECT 409.930 2792.800 410.250 2792.860 ;
        RECT 455.470 2792.800 455.790 2792.860 ;
        RECT 537.350 2793.000 537.670 2793.060 ;
        RECT 865.790 2793.000 866.110 2793.060 ;
        RECT 537.350 2792.860 866.110 2793.000 ;
        RECT 537.350 2792.800 537.670 2792.860 ;
        RECT 865.790 2792.800 866.110 2792.860 ;
        RECT 1122.010 2793.000 1122.330 2793.060 ;
        RECT 1166.170 2793.000 1166.490 2793.060 ;
        RECT 1122.010 2792.860 1166.490 2793.000 ;
        RECT 1122.010 2792.800 1122.330 2792.860 ;
        RECT 1166.170 2792.800 1166.490 2792.860 ;
        RECT 1449.085 2793.000 1449.375 2793.045 ;
        RECT 1510.725 2793.000 1511.015 2793.045 ;
        RECT 1449.085 2792.860 1511.015 2793.000 ;
        RECT 1449.085 2792.815 1449.375 2792.860 ;
        RECT 1510.725 2792.815 1511.015 2792.860 ;
        RECT 1511.185 2793.000 1511.475 2793.045 ;
        RECT 1538.785 2793.000 1539.075 2793.045 ;
        RECT 1511.185 2792.860 1539.075 2793.000 ;
        RECT 1511.185 2792.815 1511.475 2792.860 ;
        RECT 1538.785 2792.815 1539.075 2792.860 ;
        RECT 1677.230 2793.000 1677.550 2793.060 ;
        RECT 1723.690 2793.000 1724.010 2793.060 ;
        RECT 1677.230 2792.860 1724.010 2793.000 ;
        RECT 1677.230 2792.800 1677.550 2792.860 ;
        RECT 1723.690 2792.800 1724.010 2792.860 ;
        RECT 1741.170 2793.000 1741.490 2793.060 ;
        RECT 1787.170 2793.000 1787.490 2793.060 ;
        RECT 1741.170 2792.860 1787.490 2793.000 ;
        RECT 1741.170 2792.800 1741.490 2792.860 ;
        RECT 1787.170 2792.800 1787.490 2792.860 ;
        RECT 2273.390 2793.000 2273.710 2793.060 ;
        RECT 2321.690 2793.000 2322.010 2793.060 ;
        RECT 2367.230 2793.000 2367.550 2793.060 ;
        RECT 2415.070 2793.000 2415.390 2793.060 ;
        RECT 2273.390 2792.860 2415.390 2793.000 ;
        RECT 2273.390 2792.800 2273.710 2792.860 ;
        RECT 2321.690 2792.800 2322.010 2792.860 ;
        RECT 2367.230 2792.800 2367.550 2792.860 ;
        RECT 2415.070 2792.800 2415.390 2792.860 ;
        RECT 397.050 2792.660 397.370 2792.720 ;
        RECT 444.430 2792.660 444.750 2792.720 ;
        RECT 492.730 2792.660 493.050 2792.720 ;
        RECT 539.190 2792.660 539.510 2792.720 ;
        RECT 397.050 2792.520 539.510 2792.660 ;
        RECT 397.050 2792.460 397.370 2792.520 ;
        RECT 444.430 2792.460 444.750 2792.520 ;
        RECT 492.730 2792.460 493.050 2792.520 ;
        RECT 539.190 2792.460 539.510 2792.520 ;
        RECT 544.250 2792.660 544.570 2792.720 ;
        RECT 872.690 2792.660 873.010 2792.720 ;
        RECT 544.250 2792.520 873.010 2792.660 ;
        RECT 544.250 2792.460 544.570 2792.520 ;
        RECT 872.690 2792.460 873.010 2792.520 ;
        RECT 1042.430 2792.660 1042.750 2792.720 ;
        RECT 1087.510 2792.660 1087.830 2792.720 ;
        RECT 1135.810 2792.660 1136.130 2792.720 ;
        RECT 1179.970 2792.660 1180.290 2792.720 ;
        RECT 1042.430 2792.520 1180.290 2792.660 ;
        RECT 1042.430 2792.460 1042.750 2792.520 ;
        RECT 1087.510 2792.460 1087.830 2792.520 ;
        RECT 1135.810 2792.460 1136.130 2792.520 ;
        RECT 1179.970 2792.460 1180.290 2792.520 ;
        RECT 1559.485 2792.660 1559.775 2792.705 ;
        RECT 1559.485 2792.520 1586.840 2792.660 ;
        RECT 1559.485 2792.475 1559.775 2792.520 ;
        RECT 392.450 2792.320 392.770 2792.380 ;
        RECT 439.370 2792.320 439.690 2792.380 ;
        RECT 477.565 2792.320 477.855 2792.365 ;
        RECT 392.450 2792.180 477.855 2792.320 ;
        RECT 392.450 2792.120 392.770 2792.180 ;
        RECT 439.370 2792.120 439.690 2792.180 ;
        RECT 477.565 2792.135 477.855 2792.180 ;
        RECT 524.010 2792.320 524.330 2792.380 ;
        RECT 858.890 2792.320 859.210 2792.380 ;
        RECT 524.010 2792.180 859.210 2792.320 ;
        RECT 524.010 2792.120 524.330 2792.180 ;
        RECT 858.890 2792.120 859.210 2792.180 ;
        RECT 1055.770 2792.320 1056.090 2792.380 ;
        RECT 1058.990 2792.320 1059.310 2792.380 ;
        RECT 1105.450 2792.320 1105.770 2792.380 ;
        RECT 1152.370 2792.320 1152.690 2792.380 ;
        RECT 1055.770 2792.180 1152.690 2792.320 ;
        RECT 1055.770 2792.120 1056.090 2792.180 ;
        RECT 1058.990 2792.120 1059.310 2792.180 ;
        RECT 1105.450 2792.120 1105.770 2792.180 ;
        RECT 1152.370 2792.120 1152.690 2792.180 ;
        RECT 1420.550 2792.320 1420.870 2792.380 ;
        RECT 1449.085 2792.320 1449.375 2792.365 ;
        RECT 1420.550 2792.180 1449.375 2792.320 ;
        RECT 1420.550 2792.120 1420.870 2792.180 ;
        RECT 1449.085 2792.135 1449.375 2792.180 ;
        RECT 1538.785 2792.320 1539.075 2792.365 ;
        RECT 1559.025 2792.320 1559.315 2792.365 ;
        RECT 1538.785 2792.180 1559.315 2792.320 ;
        RECT 1586.700 2792.320 1586.840 2792.520 ;
        RECT 1587.085 2792.475 1587.375 2792.705 ;
        RECT 1634.925 2792.660 1635.215 2792.705 ;
        RECT 1652.850 2792.660 1653.170 2792.720 ;
        RECT 1690.570 2792.660 1690.890 2792.720 ;
        RECT 1695.170 2792.660 1695.490 2792.720 ;
        RECT 1704.385 2792.660 1704.675 2792.705 ;
        RECT 1634.925 2792.520 1655.840 2792.660 ;
        RECT 1634.925 2792.475 1635.215 2792.520 ;
        RECT 1587.160 2792.320 1587.300 2792.475 ;
        RECT 1652.850 2792.460 1653.170 2792.520 ;
        RECT 1586.700 2792.180 1587.300 2792.320 ;
        RECT 1538.785 2792.135 1539.075 2792.180 ;
        RECT 1559.025 2792.135 1559.315 2792.180 ;
        RECT 368.530 2791.980 368.850 2792.040 ;
        RECT 433.390 2791.980 433.710 2792.040 ;
        RECT 478.470 2791.980 478.790 2792.040 ;
        RECT 504.705 2791.980 504.995 2792.025 ;
        RECT 368.530 2791.840 403.720 2791.980 ;
        RECT 368.530 2791.780 368.850 2791.840 ;
        RECT 362.090 2791.300 362.410 2791.360 ;
        RECT 391.085 2791.300 391.375 2791.345 ;
        RECT 362.090 2791.160 391.375 2791.300 ;
        RECT 403.580 2791.300 403.720 2791.840 ;
        RECT 433.390 2791.840 504.995 2791.980 ;
        RECT 433.390 2791.780 433.710 2791.840 ;
        RECT 478.470 2791.780 478.790 2791.840 ;
        RECT 504.705 2791.795 504.995 2791.840 ;
        RECT 510.210 2791.980 510.530 2792.040 ;
        RECT 851.990 2791.980 852.310 2792.040 ;
        RECT 510.210 2791.840 852.310 2791.980 ;
        RECT 510.210 2791.780 510.530 2791.840 ;
        RECT 851.990 2791.780 852.310 2791.840 ;
        RECT 1060.385 2791.980 1060.675 2792.025 ;
        RECT 1100.850 2791.980 1101.170 2792.040 ;
        RECT 1146.390 2791.980 1146.710 2792.040 ;
        RECT 1060.385 2791.840 1146.710 2791.980 ;
        RECT 1060.385 2791.795 1060.675 2791.840 ;
        RECT 1100.850 2791.780 1101.170 2791.840 ;
        RECT 1146.390 2791.780 1146.710 2791.840 ;
        RECT 1549.350 2791.980 1549.670 2792.040 ;
        RECT 1596.270 2791.980 1596.590 2792.040 ;
        RECT 1549.350 2791.840 1596.590 2791.980 ;
        RECT 1655.700 2791.980 1655.840 2792.520 ;
        RECT 1690.570 2792.520 1704.675 2792.660 ;
        RECT 1690.570 2792.460 1690.890 2792.520 ;
        RECT 1695.170 2792.460 1695.490 2792.520 ;
        RECT 1704.385 2792.475 1704.675 2792.520 ;
        RECT 2210.845 2792.660 2211.135 2792.705 ;
        RECT 2268.330 2792.660 2268.650 2792.720 ;
        RECT 2315.250 2792.660 2315.570 2792.720 ;
        RECT 2361.250 2792.660 2361.570 2792.720 ;
        RECT 2408.170 2792.660 2408.490 2792.720 ;
        RECT 2210.845 2792.520 2408.490 2792.660 ;
        RECT 2210.845 2792.475 2211.135 2792.520 ;
        RECT 2268.330 2792.460 2268.650 2792.520 ;
        RECT 2315.250 2792.460 2315.570 2792.520 ;
        RECT 2361.250 2792.460 2361.570 2792.520 ;
        RECT 2408.170 2792.460 2408.490 2792.520 ;
        RECT 1662.510 2792.320 1662.830 2792.380 ;
        RECT 1706.210 2792.320 1706.530 2792.380 ;
        RECT 1752.670 2792.320 1752.990 2792.380 ;
        RECT 1662.510 2792.180 1752.990 2792.320 ;
        RECT 1662.510 2792.120 1662.830 2792.180 ;
        RECT 1706.210 2792.120 1706.530 2792.180 ;
        RECT 1752.670 2792.120 1752.990 2792.180 ;
        RECT 2266.490 2792.320 2266.810 2792.380 ;
        RECT 2280.765 2792.320 2281.055 2792.365 ;
        RECT 2266.490 2792.180 2281.055 2792.320 ;
        RECT 2266.490 2792.120 2266.810 2792.180 ;
        RECT 2280.765 2792.135 2281.055 2792.180 ;
        RECT 2284.430 2792.320 2284.750 2792.380 ;
        RECT 2333.650 2792.320 2333.970 2792.380 ;
        RECT 2284.430 2792.180 2333.970 2792.320 ;
        RECT 2284.430 2792.120 2284.750 2792.180 ;
        RECT 2333.650 2792.120 2333.970 2792.180 ;
        RECT 2334.125 2792.320 2334.415 2792.365 ;
        RECT 2340.090 2792.320 2340.410 2792.380 ;
        RECT 2347.005 2792.320 2347.295 2792.365 ;
        RECT 2334.125 2792.180 2347.295 2792.320 ;
        RECT 2334.125 2792.135 2334.415 2792.180 ;
        RECT 2340.090 2792.120 2340.410 2792.180 ;
        RECT 2347.005 2792.135 2347.295 2792.180 ;
        RECT 2347.450 2792.320 2347.770 2792.380 ;
        RECT 2394.830 2792.320 2395.150 2792.380 ;
        RECT 2347.450 2792.180 2395.150 2792.320 ;
        RECT 2347.450 2792.120 2347.770 2792.180 ;
        RECT 2394.830 2792.120 2395.150 2792.180 ;
        RECT 1699.310 2791.980 1699.630 2792.040 ;
        RECT 2326.750 2791.980 2327.070 2792.040 ;
        RECT 2374.130 2791.980 2374.450 2792.040 ;
        RECT 2415.070 2791.980 2415.390 2792.040 ;
        RECT 1655.700 2791.840 1738.640 2791.980 ;
        RECT 1549.350 2791.780 1549.670 2791.840 ;
        RECT 1596.270 2791.780 1596.590 2791.840 ;
        RECT 1699.310 2791.780 1699.630 2791.840 ;
        RECT 403.950 2791.640 404.270 2791.700 ;
        RECT 450.410 2791.640 450.730 2791.700 ;
        RECT 501.010 2791.640 501.330 2791.700 ;
        RECT 403.950 2791.500 501.330 2791.640 ;
        RECT 403.950 2791.440 404.270 2791.500 ;
        RECT 450.410 2791.440 450.730 2791.500 ;
        RECT 501.010 2791.440 501.330 2791.500 ;
        RECT 501.930 2791.640 502.250 2791.700 ;
        RECT 845.090 2791.640 845.410 2791.700 ;
        RECT 1065.430 2791.640 1065.750 2791.700 ;
        RECT 1111.430 2791.640 1111.750 2791.700 ;
        RECT 1159.270 2791.640 1159.590 2791.700 ;
        RECT 501.930 2791.500 845.410 2791.640 ;
        RECT 501.930 2791.440 502.250 2791.500 ;
        RECT 845.090 2791.440 845.410 2791.500 ;
        RECT 1034.240 2791.500 1159.590 2791.640 ;
        RECT 414.530 2791.300 414.850 2791.360 ;
        RECT 462.370 2791.300 462.690 2791.360 ;
        RECT 403.580 2791.160 462.690 2791.300 ;
        RECT 362.090 2791.100 362.410 2791.160 ;
        RECT 391.085 2791.115 391.375 2791.160 ;
        RECT 414.530 2791.100 414.850 2791.160 ;
        RECT 462.370 2791.100 462.690 2791.160 ;
        RECT 489.050 2791.300 489.370 2791.360 ;
        RECT 838.190 2791.300 838.510 2791.360 ;
        RECT 489.050 2791.160 838.510 2791.300 ;
        RECT 489.050 2791.100 489.370 2791.160 ;
        RECT 838.190 2791.100 838.510 2791.160 ;
        RECT 371.290 2790.960 371.610 2791.020 ;
        RECT 745.270 2790.960 745.590 2791.020 ;
        RECT 371.290 2790.820 745.590 2790.960 ;
        RECT 371.290 2790.760 371.610 2790.820 ;
        RECT 745.270 2790.760 745.590 2790.820 ;
        RECT 1018.970 2790.960 1019.290 2791.020 ;
        RECT 1034.240 2790.960 1034.380 2791.500 ;
        RECT 1065.430 2791.440 1065.750 2791.500 ;
        RECT 1111.430 2791.440 1111.750 2791.500 ;
        RECT 1159.270 2791.440 1159.590 2791.500 ;
        RECT 1511.185 2791.640 1511.475 2791.685 ;
        RECT 1654.705 2791.640 1654.995 2791.685 ;
        RECT 1511.185 2791.500 1654.995 2791.640 ;
        RECT 1511.185 2791.455 1511.475 2791.500 ;
        RECT 1654.705 2791.455 1654.995 2791.500 ;
        RECT 1682.290 2791.640 1682.610 2791.700 ;
        RECT 1728.750 2791.640 1729.070 2791.700 ;
        RECT 1682.290 2791.500 1729.070 2791.640 ;
        RECT 1738.500 2791.640 1738.640 2791.840 ;
        RECT 2279.920 2791.840 2415.390 2791.980 ;
        RECT 2279.920 2791.700 2280.060 2791.840 ;
        RECT 2326.750 2791.780 2327.070 2791.840 ;
        RECT 2374.130 2791.780 2374.450 2791.840 ;
        RECT 2415.070 2791.780 2415.390 2791.840 ;
        RECT 1747.610 2791.640 1747.930 2791.700 ;
        RECT 1794.070 2791.640 1794.390 2791.700 ;
        RECT 1738.500 2791.500 1794.390 2791.640 ;
        RECT 1682.290 2791.440 1682.610 2791.500 ;
        RECT 1728.750 2791.440 1729.070 2791.500 ;
        RECT 1747.610 2791.440 1747.930 2791.500 ;
        RECT 1794.070 2791.440 1794.390 2791.500 ;
        RECT 2090.770 2791.640 2091.090 2791.700 ;
        RECT 2138.625 2791.640 2138.915 2791.685 ;
        RECT 2090.770 2791.500 2138.915 2791.640 ;
        RECT 2090.770 2791.440 2091.090 2791.500 ;
        RECT 2138.625 2791.455 2138.915 2791.500 ;
        RECT 2139.085 2791.640 2139.375 2791.685 ;
        RECT 2181.405 2791.640 2181.695 2791.685 ;
        RECT 2139.085 2791.500 2181.695 2791.640 ;
        RECT 2139.085 2791.455 2139.375 2791.500 ;
        RECT 2181.405 2791.455 2181.695 2791.500 ;
        RECT 2262.825 2791.640 2263.115 2791.685 ;
        RECT 2279.830 2791.640 2280.150 2791.700 ;
        RECT 2262.825 2791.500 2280.150 2791.640 ;
        RECT 2262.825 2791.455 2263.115 2791.500 ;
        RECT 2279.830 2791.440 2280.150 2791.500 ;
        RECT 2301.450 2791.640 2301.770 2791.700 ;
        RECT 2435.770 2791.640 2436.090 2791.700 ;
        RECT 2301.450 2791.500 2436.090 2791.640 ;
        RECT 2301.450 2791.440 2301.770 2791.500 ;
        RECT 2435.770 2791.440 2436.090 2791.500 ;
        RECT 1034.610 2791.300 1034.930 2791.360 ;
        RECT 1076.470 2791.300 1076.790 2791.360 ;
        RECT 1122.010 2791.300 1122.330 2791.360 ;
        RECT 1034.610 2791.160 1122.330 2791.300 ;
        RECT 1034.610 2791.100 1034.930 2791.160 ;
        RECT 1076.470 2791.100 1076.790 2791.160 ;
        RECT 1122.010 2791.100 1122.330 2791.160 ;
        RECT 1146.390 2791.300 1146.710 2791.360 ;
        RECT 1193.770 2791.300 1194.090 2791.360 ;
        RECT 1146.390 2791.160 1194.090 2791.300 ;
        RECT 1146.390 2791.100 1146.710 2791.160 ;
        RECT 1193.770 2791.100 1194.090 2791.160 ;
        RECT 1411.350 2791.300 1411.670 2791.360 ;
        RECT 1587.070 2791.300 1587.390 2791.360 ;
        RECT 1670.330 2791.300 1670.650 2791.360 ;
        RECT 1718.170 2791.300 1718.490 2791.360 ;
        RECT 1724.610 2791.300 1724.930 2791.360 ;
        RECT 1411.350 2791.160 1587.390 2791.300 ;
        RECT 1411.350 2791.100 1411.670 2791.160 ;
        RECT 1587.070 2791.100 1587.390 2791.160 ;
        RECT 1669.040 2791.160 1724.930 2791.300 ;
        RECT 1728.840 2791.300 1728.980 2791.440 ;
        RECT 1773.370 2791.300 1773.690 2791.360 ;
        RECT 1728.840 2791.160 1773.690 2791.300 ;
        RECT 1018.970 2790.820 1034.380 2790.960 ;
        RECT 1069.570 2790.960 1069.890 2791.020 ;
        RECT 1118.330 2790.960 1118.650 2791.020 ;
        RECT 1159.270 2790.960 1159.590 2791.020 ;
        RECT 1069.570 2790.820 1159.590 2790.960 ;
        RECT 1018.970 2790.760 1019.290 2790.820 ;
        RECT 1069.570 2790.760 1069.890 2790.820 ;
        RECT 1118.330 2790.760 1118.650 2790.820 ;
        RECT 1159.270 2790.760 1159.590 2790.820 ;
        RECT 1425.150 2790.960 1425.470 2791.020 ;
        RECT 1600.870 2790.960 1601.190 2791.020 ;
        RECT 1659.290 2790.960 1659.610 2791.020 ;
        RECT 1662.510 2790.960 1662.830 2791.020 ;
        RECT 1425.150 2790.820 1601.190 2790.960 ;
        RECT 1425.150 2790.760 1425.470 2790.820 ;
        RECT 1600.870 2790.760 1601.190 2790.820 ;
        RECT 1624.420 2790.820 1662.830 2790.960 ;
        RECT 384.630 2790.620 384.950 2790.680 ;
        RECT 765.970 2790.620 766.290 2790.680 ;
        RECT 384.630 2790.480 766.290 2790.620 ;
        RECT 384.630 2790.420 384.950 2790.480 ;
        RECT 765.970 2790.420 766.290 2790.480 ;
        RECT 1411.810 2790.620 1412.130 2790.680 ;
        RECT 1613.290 2790.620 1613.610 2790.680 ;
        RECT 1624.420 2790.620 1624.560 2790.820 ;
        RECT 1659.290 2790.760 1659.610 2790.820 ;
        RECT 1662.510 2790.760 1662.830 2790.820 ;
        RECT 1411.810 2790.480 1624.560 2790.620 ;
        RECT 1624.790 2790.620 1625.110 2790.680 ;
        RECT 1669.040 2790.620 1669.180 2791.160 ;
        RECT 1670.330 2791.100 1670.650 2791.160 ;
        RECT 1718.170 2791.100 1718.490 2791.160 ;
        RECT 1724.610 2791.100 1724.930 2791.160 ;
        RECT 1773.370 2791.100 1773.690 2791.160 ;
        RECT 1869.985 2791.300 1870.275 2791.345 ;
        RECT 1917.365 2791.300 1917.655 2791.345 ;
        RECT 1869.985 2791.160 1917.655 2791.300 ;
        RECT 1869.985 2791.115 1870.275 2791.160 ;
        RECT 1917.365 2791.115 1917.655 2791.160 ;
        RECT 2266.950 2791.300 2267.270 2791.360 ;
        RECT 2428.870 2791.300 2429.190 2791.360 ;
        RECT 2266.950 2791.160 2429.190 2791.300 ;
        RECT 2266.950 2791.100 2267.270 2791.160 ;
        RECT 2428.870 2791.100 2429.190 2791.160 ;
        RECT 1669.410 2790.960 1669.730 2791.020 ;
        RECT 1712.650 2790.960 1712.970 2791.020 ;
        RECT 1759.570 2790.960 1759.890 2791.020 ;
        RECT 1669.410 2790.820 1759.890 2790.960 ;
        RECT 1669.410 2790.760 1669.730 2790.820 ;
        RECT 1712.650 2790.760 1712.970 2790.820 ;
        RECT 1759.570 2790.760 1759.890 2790.820 ;
        RECT 1797.290 2790.960 1797.610 2791.020 ;
        RECT 2387.470 2790.960 2387.790 2791.020 ;
        RECT 1797.290 2790.820 2387.790 2790.960 ;
        RECT 1797.290 2790.760 1797.610 2790.820 ;
        RECT 2387.470 2790.760 2387.790 2790.820 ;
        RECT 2394.830 2790.960 2395.150 2791.020 ;
        RECT 2442.670 2790.960 2442.990 2791.020 ;
        RECT 2394.830 2790.820 2442.990 2790.960 ;
        RECT 2394.830 2790.760 2395.150 2790.820 ;
        RECT 2442.670 2790.760 2442.990 2790.820 ;
        RECT 1624.790 2790.480 1669.180 2790.620 ;
        RECT 1724.610 2790.620 1724.930 2790.680 ;
        RECT 1760.030 2790.620 1760.350 2790.680 ;
        RECT 1724.610 2790.480 1760.350 2790.620 ;
        RECT 1411.810 2790.420 1412.130 2790.480 ;
        RECT 1613.290 2790.420 1613.610 2790.480 ;
        RECT 1624.790 2790.420 1625.110 2790.480 ;
        RECT 1724.610 2790.420 1724.930 2790.480 ;
        RECT 1760.030 2790.420 1760.350 2790.480 ;
        RECT 1783.490 2790.620 1783.810 2790.680 ;
        RECT 2373.670 2790.620 2373.990 2790.680 ;
        RECT 1783.490 2790.480 2373.990 2790.620 ;
        RECT 1783.490 2790.420 1783.810 2790.480 ;
        RECT 2373.670 2790.420 2373.990 2790.480 ;
        RECT 2377.350 2790.620 2377.670 2790.680 ;
        RECT 2421.970 2790.620 2422.290 2790.680 ;
        RECT 2377.350 2790.480 2422.290 2790.620 ;
        RECT 2377.350 2790.420 2377.670 2790.480 ;
        RECT 2421.970 2790.420 2422.290 2790.480 ;
        RECT 396.590 2790.280 396.910 2790.340 ;
        RECT 786.670 2790.280 786.990 2790.340 ;
        RECT 396.590 2790.140 786.990 2790.280 ;
        RECT 396.590 2790.080 396.910 2790.140 ;
        RECT 786.670 2790.080 786.990 2790.140 ;
        RECT 1420.090 2790.280 1420.410 2790.340 ;
        RECT 1636.750 2790.280 1637.070 2790.340 ;
        RECT 1420.090 2790.140 1637.070 2790.280 ;
        RECT 1420.090 2790.080 1420.410 2790.140 ;
        RECT 1636.750 2790.080 1637.070 2790.140 ;
        RECT 1704.385 2790.280 1704.675 2790.325 ;
        RECT 1741.170 2790.280 1741.490 2790.340 ;
        RECT 1704.385 2790.140 1741.490 2790.280 ;
        RECT 1704.385 2790.095 1704.675 2790.140 ;
        RECT 1741.170 2790.080 1741.490 2790.140 ;
        RECT 1790.390 2790.280 1790.710 2790.340 ;
        RECT 2380.570 2790.280 2380.890 2790.340 ;
        RECT 1790.390 2790.140 2380.890 2790.280 ;
        RECT 1790.390 2790.080 1790.710 2790.140 ;
        RECT 2380.570 2790.080 2380.890 2790.140 ;
        RECT 406.250 2789.940 406.570 2790.000 ;
        RECT 807.370 2789.940 807.690 2790.000 ;
        RECT 406.250 2789.800 807.690 2789.940 ;
        RECT 406.250 2789.740 406.570 2789.800 ;
        RECT 807.370 2789.740 807.690 2789.800 ;
        RECT 1419.630 2789.940 1419.950 2790.000 ;
        RECT 1642.730 2789.940 1643.050 2790.000 ;
        RECT 1419.630 2789.800 1643.050 2789.940 ;
        RECT 1419.630 2789.740 1419.950 2789.800 ;
        RECT 1642.730 2789.740 1643.050 2789.800 ;
        RECT 1654.705 2789.940 1654.995 2789.985 ;
        RECT 1669.885 2789.940 1670.175 2789.985 ;
        RECT 1654.705 2789.800 1670.175 2789.940 ;
        RECT 1654.705 2789.755 1654.995 2789.800 ;
        RECT 1669.885 2789.755 1670.175 2789.800 ;
        RECT 1797.750 2789.940 1798.070 2790.000 ;
        RECT 2394.370 2789.940 2394.690 2790.000 ;
        RECT 1797.750 2789.800 2394.690 2789.940 ;
        RECT 1797.750 2789.740 1798.070 2789.800 ;
        RECT 2394.370 2789.740 2394.690 2789.800 ;
        RECT 477.565 2789.600 477.855 2789.645 ;
        RECT 484.910 2789.600 485.230 2789.660 ;
        RECT 534.590 2789.600 534.910 2789.660 ;
        RECT 477.565 2789.460 534.910 2789.600 ;
        RECT 477.565 2789.415 477.855 2789.460 ;
        RECT 484.910 2789.400 485.230 2789.460 ;
        RECT 534.590 2789.400 534.910 2789.460 ;
        RECT 539.190 2789.600 539.510 2789.660 ;
        RECT 717.670 2789.600 717.990 2789.660 ;
        RECT 539.190 2789.460 717.990 2789.600 ;
        RECT 539.190 2789.400 539.510 2789.460 ;
        RECT 717.670 2789.400 717.990 2789.460 ;
        RECT 1549.810 2789.600 1550.130 2789.660 ;
        RECT 1642.270 2789.600 1642.590 2789.660 ;
        RECT 1549.810 2789.460 1642.590 2789.600 ;
        RECT 1549.810 2789.400 1550.130 2789.460 ;
        RECT 1642.270 2789.400 1642.590 2789.460 ;
        RECT 1645.490 2789.600 1645.810 2789.660 ;
        RECT 1648.250 2789.600 1648.570 2789.660 ;
        RECT 1690.570 2789.600 1690.890 2789.660 ;
        RECT 1645.490 2789.460 1690.890 2789.600 ;
        RECT 1645.490 2789.400 1645.810 2789.460 ;
        RECT 1648.250 2789.400 1648.570 2789.460 ;
        RECT 1690.570 2789.400 1690.890 2789.460 ;
        RECT 1762.790 2789.600 1763.110 2789.660 ;
        RECT 2380.570 2789.600 2380.890 2789.660 ;
        RECT 1762.790 2789.460 2380.890 2789.600 ;
        RECT 1762.790 2789.400 1763.110 2789.460 ;
        RECT 2380.570 2789.400 2380.890 2789.460 ;
        RECT 418.670 2789.260 418.990 2789.320 ;
        RECT 828.070 2789.260 828.390 2789.320 ;
        RECT 418.670 2789.120 828.390 2789.260 ;
        RECT 418.670 2789.060 418.990 2789.120 ;
        RECT 828.070 2789.060 828.390 2789.120 ;
        RECT 1010.690 2789.260 1011.010 2789.320 ;
        RECT 1055.770 2789.260 1056.090 2789.320 ;
        RECT 1010.690 2789.120 1056.090 2789.260 ;
        RECT 1010.690 2789.060 1011.010 2789.120 ;
        RECT 1055.770 2789.060 1056.090 2789.120 ;
        RECT 1410.890 2789.260 1411.210 2789.320 ;
        RECT 1486.805 2789.260 1487.095 2789.305 ;
        RECT 2218.190 2789.260 2218.510 2789.320 ;
        RECT 2402.650 2789.260 2402.970 2789.320 ;
        RECT 1410.890 2789.120 1487.095 2789.260 ;
        RECT 1410.890 2789.060 1411.210 2789.120 ;
        RECT 1486.805 2789.075 1487.095 2789.120 ;
        RECT 1583.020 2789.120 2211.520 2789.260 ;
        RECT 413.610 2788.920 413.930 2788.980 ;
        RECT 465.590 2788.920 465.910 2788.980 ;
        RECT 413.610 2788.780 465.910 2788.920 ;
        RECT 413.610 2788.720 413.930 2788.780 ;
        RECT 465.590 2788.720 465.910 2788.780 ;
        RECT 475.250 2788.920 475.570 2788.980 ;
        RECT 520.790 2788.920 521.110 2788.980 ;
        RECT 475.250 2788.780 521.110 2788.920 ;
        RECT 475.250 2788.720 475.570 2788.780 ;
        RECT 520.790 2788.720 521.110 2788.780 ;
        RECT 627.510 2788.920 627.830 2788.980 ;
        RECT 1042.430 2788.920 1042.750 2788.980 ;
        RECT 627.510 2788.780 1042.750 2788.920 ;
        RECT 627.510 2788.720 627.830 2788.780 ;
        RECT 1042.430 2788.720 1042.750 2788.780 ;
        RECT 1417.790 2788.920 1418.110 2788.980 ;
        RECT 1535.105 2788.920 1535.395 2788.965 ;
        RECT 1583.020 2788.920 1583.160 2789.120 ;
        RECT 2090.785 2788.920 2091.075 2788.965 ;
        RECT 2210.845 2788.920 2211.135 2788.965 ;
        RECT 1417.790 2788.780 1512.320 2788.920 ;
        RECT 1417.790 2788.720 1418.110 2788.780 ;
        RECT 399.810 2788.580 400.130 2788.640 ;
        RECT 444.890 2788.580 445.210 2788.640 ;
        RECT 399.810 2788.440 445.210 2788.580 ;
        RECT 399.810 2788.380 400.130 2788.440 ;
        RECT 444.890 2788.380 445.210 2788.440 ;
        RECT 606.810 2788.580 607.130 2788.640 ;
        RECT 1034.610 2788.580 1034.930 2788.640 ;
        RECT 606.810 2788.440 1034.930 2788.580 ;
        RECT 606.810 2788.380 607.130 2788.440 ;
        RECT 1034.610 2788.380 1034.930 2788.440 ;
        RECT 1045.190 2788.580 1045.510 2788.640 ;
        RECT 1090.270 2788.580 1090.590 2788.640 ;
        RECT 1045.190 2788.440 1090.590 2788.580 ;
        RECT 1045.190 2788.380 1045.510 2788.440 ;
        RECT 1090.270 2788.380 1090.590 2788.440 ;
        RECT 1418.250 2788.580 1418.570 2788.640 ;
        RECT 1511.185 2788.580 1511.475 2788.625 ;
        RECT 1418.250 2788.440 1511.475 2788.580 ;
        RECT 1512.180 2788.580 1512.320 2788.780 ;
        RECT 1535.105 2788.780 1583.160 2788.920 ;
        RECT 1583.480 2788.780 2091.075 2788.920 ;
        RECT 1535.105 2788.735 1535.395 2788.780 ;
        RECT 1583.480 2788.580 1583.620 2788.780 ;
        RECT 2090.785 2788.735 2091.075 2788.780 ;
        RECT 2186.540 2788.780 2211.135 2788.920 ;
        RECT 2211.380 2788.920 2211.520 2789.120 ;
        RECT 2218.190 2789.120 2402.970 2789.260 ;
        RECT 2218.190 2789.060 2218.510 2789.120 ;
        RECT 2402.650 2789.060 2402.970 2789.120 ;
        RECT 2235.670 2788.920 2235.990 2788.980 ;
        RECT 2211.380 2788.780 2235.990 2788.920 ;
        RECT 1512.180 2788.440 1583.620 2788.580 ;
        RECT 1418.250 2788.380 1418.570 2788.440 ;
        RECT 1511.185 2788.395 1511.475 2788.440 ;
        RECT 1869.985 2788.395 1870.275 2788.625 ;
        RECT 2091.245 2788.580 2091.535 2788.625 ;
        RECT 2186.540 2788.580 2186.680 2788.780 ;
        RECT 2210.845 2788.735 2211.135 2788.780 ;
        RECT 2235.670 2788.720 2235.990 2788.780 ;
        RECT 2238.890 2788.920 2239.210 2788.980 ;
        RECT 2267.425 2788.920 2267.715 2788.965 ;
        RECT 2408.170 2788.920 2408.490 2788.980 ;
        RECT 2238.890 2788.780 2263.500 2788.920 ;
        RECT 2238.890 2788.720 2239.210 2788.780 ;
        RECT 2076.600 2788.440 2091.000 2788.580 ;
        RECT 378.650 2788.240 378.970 2788.300 ;
        RECT 424.190 2788.240 424.510 2788.300 ;
        RECT 378.650 2788.100 424.510 2788.240 ;
        RECT 378.650 2788.040 378.970 2788.100 ;
        RECT 424.190 2788.040 424.510 2788.100 ;
        RECT 455.470 2788.240 455.790 2788.300 ;
        RECT 500.090 2788.240 500.410 2788.300 ;
        RECT 455.470 2788.100 500.410 2788.240 ;
        RECT 455.470 2788.040 455.790 2788.100 ;
        RECT 500.090 2788.040 500.410 2788.100 ;
        RECT 501.010 2788.240 501.330 2788.300 ;
        RECT 541.490 2788.240 541.810 2788.300 ;
        RECT 501.010 2788.100 541.810 2788.240 ;
        RECT 501.010 2788.040 501.330 2788.100 ;
        RECT 541.490 2788.040 541.810 2788.100 ;
        RECT 586.110 2788.240 586.430 2788.300 ;
        RECT 1018.970 2788.240 1019.290 2788.300 ;
        RECT 586.110 2788.100 1019.290 2788.240 ;
        RECT 586.110 2788.040 586.430 2788.100 ;
        RECT 1018.970 2788.040 1019.290 2788.100 ;
        RECT 1024.490 2788.240 1024.810 2788.300 ;
        RECT 1069.570 2788.240 1069.890 2788.300 ;
        RECT 1024.490 2788.100 1069.890 2788.240 ;
        RECT 1024.490 2788.040 1024.810 2788.100 ;
        RECT 1069.570 2788.040 1069.890 2788.100 ;
        RECT 1486.805 2788.240 1487.095 2788.285 ;
        RECT 1535.105 2788.240 1535.395 2788.285 ;
        RECT 1486.805 2788.100 1535.395 2788.240 ;
        RECT 1486.805 2788.055 1487.095 2788.100 ;
        RECT 1535.105 2788.055 1535.395 2788.100 ;
        RECT 1617.890 2788.240 1618.210 2788.300 ;
        RECT 1669.410 2788.240 1669.730 2788.300 ;
        RECT 1617.890 2788.100 1669.730 2788.240 ;
        RECT 1617.890 2788.040 1618.210 2788.100 ;
        RECT 1669.410 2788.040 1669.730 2788.100 ;
        RECT 1669.885 2788.240 1670.175 2788.285 ;
        RECT 1669.885 2788.100 1702.300 2788.240 ;
        RECT 1669.885 2788.055 1670.175 2788.100 ;
        RECT 390.610 2787.900 390.930 2787.960 ;
        RECT 431.090 2787.900 431.410 2787.960 ;
        RECT 390.610 2787.760 431.410 2787.900 ;
        RECT 390.610 2787.700 390.930 2787.760 ;
        RECT 431.090 2787.700 431.410 2787.760 ;
        RECT 479.390 2787.900 479.710 2787.960 ;
        RECT 1007.470 2787.900 1007.790 2787.960 ;
        RECT 479.390 2787.760 1007.790 2787.900 ;
        RECT 479.390 2787.700 479.710 2787.760 ;
        RECT 1007.470 2787.700 1007.790 2787.760 ;
        RECT 1038.290 2787.900 1038.610 2787.960 ;
        RECT 1083.370 2787.900 1083.690 2787.960 ;
        RECT 1038.290 2787.760 1083.690 2787.900 ;
        RECT 1038.290 2787.700 1038.610 2787.760 ;
        RECT 1083.370 2787.700 1083.690 2787.760 ;
        RECT 1548.890 2787.900 1549.210 2787.960 ;
        RECT 1628.470 2787.900 1628.790 2787.960 ;
        RECT 1548.890 2787.760 1628.790 2787.900 ;
        RECT 1548.890 2787.700 1549.210 2787.760 ;
        RECT 1628.470 2787.700 1628.790 2787.760 ;
        RECT 1631.690 2787.900 1632.010 2787.960 ;
        RECT 1677.230 2787.900 1677.550 2787.960 ;
        RECT 1631.690 2787.760 1677.550 2787.900 ;
        RECT 1631.690 2787.700 1632.010 2787.760 ;
        RECT 1677.230 2787.700 1677.550 2787.760 ;
        RECT 1702.160 2787.560 1702.300 2788.100 ;
        RECT 1745.400 2788.100 1780.500 2788.240 ;
        RECT 1738.885 2787.900 1739.175 2787.945 ;
        RECT 1745.400 2787.900 1745.540 2788.100 ;
        RECT 1738.885 2787.760 1745.540 2787.900 ;
        RECT 1738.885 2787.715 1739.175 2787.760 ;
        RECT 1738.425 2787.560 1738.715 2787.605 ;
        RECT 1702.160 2787.420 1738.715 2787.560 ;
        RECT 1780.360 2787.560 1780.500 2788.100 ;
        RECT 1828.110 2788.040 1828.430 2788.300 ;
        RECT 1869.510 2788.240 1869.830 2788.300 ;
        RECT 1870.060 2788.240 1870.200 2788.395 ;
        RECT 1869.510 2788.100 1870.200 2788.240 ;
        RECT 1917.825 2788.240 1918.115 2788.285 ;
        RECT 1931.625 2788.240 1931.915 2788.285 ;
        RECT 1917.825 2788.100 1931.915 2788.240 ;
        RECT 1869.510 2788.040 1869.830 2788.100 ;
        RECT 1917.825 2788.055 1918.115 2788.100 ;
        RECT 1931.625 2788.055 1931.915 2788.100 ;
        RECT 1932.085 2788.240 1932.375 2788.285 ;
        RECT 2028.225 2788.240 2028.515 2788.285 ;
        RECT 2042.025 2788.240 2042.315 2788.285 ;
        RECT 1932.085 2788.100 1966.340 2788.240 ;
        RECT 1932.085 2788.055 1932.375 2788.100 ;
        RECT 1828.200 2787.560 1828.340 2788.040 ;
        RECT 1966.200 2787.900 1966.340 2788.100 ;
        RECT 2028.225 2788.100 2042.315 2788.240 ;
        RECT 2028.225 2788.055 2028.515 2788.100 ;
        RECT 2042.025 2788.055 2042.315 2788.100 ;
        RECT 2042.485 2788.240 2042.775 2788.285 ;
        RECT 2076.600 2788.240 2076.740 2788.440 ;
        RECT 2090.860 2788.300 2091.000 2788.440 ;
        RECT 2091.245 2788.440 2186.680 2788.580 ;
        RECT 2255.925 2788.580 2256.215 2788.625 ;
        RECT 2262.825 2788.580 2263.115 2788.625 ;
        RECT 2255.925 2788.440 2263.115 2788.580 ;
        RECT 2263.360 2788.580 2263.500 2788.780 ;
        RECT 2267.425 2788.780 2408.490 2788.920 ;
        RECT 2267.425 2788.735 2267.715 2788.780 ;
        RECT 2408.170 2788.720 2408.490 2788.780 ;
        RECT 2415.070 2788.580 2415.390 2788.640 ;
        RECT 2263.360 2788.440 2415.390 2788.580 ;
        RECT 2091.245 2788.395 2091.535 2788.440 ;
        RECT 2255.925 2788.395 2256.215 2788.440 ;
        RECT 2262.825 2788.395 2263.115 2788.440 ;
        RECT 2415.070 2788.380 2415.390 2788.440 ;
        RECT 2042.485 2788.100 2076.740 2788.240 ;
        RECT 2042.485 2788.055 2042.775 2788.100 ;
        RECT 2090.770 2788.040 2091.090 2788.300 ;
        RECT 2138.625 2788.240 2138.915 2788.285 ;
        RECT 2139.085 2788.240 2139.375 2788.285 ;
        RECT 2138.625 2788.100 2139.375 2788.240 ;
        RECT 2138.625 2788.055 2138.915 2788.100 ;
        RECT 2139.085 2788.055 2139.375 2788.100 ;
        RECT 2231.990 2788.240 2232.310 2788.300 ;
        RECT 2267.425 2788.240 2267.715 2788.285 ;
        RECT 2231.990 2788.100 2267.715 2788.240 ;
        RECT 2231.990 2788.040 2232.310 2788.100 ;
        RECT 2267.425 2788.055 2267.715 2788.100 ;
        RECT 2294.090 2788.240 2294.410 2788.300 ;
        RECT 2333.205 2788.240 2333.495 2788.285 ;
        RECT 2294.090 2788.100 2333.495 2788.240 ;
        RECT 2294.090 2788.040 2294.410 2788.100 ;
        RECT 2333.205 2788.055 2333.495 2788.100 ;
        RECT 2333.650 2788.240 2333.970 2788.300 ;
        RECT 2377.350 2788.240 2377.670 2788.300 ;
        RECT 2333.650 2788.100 2377.670 2788.240 ;
        RECT 2333.650 2788.040 2333.970 2788.100 ;
        RECT 2377.350 2788.040 2377.670 2788.100 ;
        RECT 1980.385 2787.900 1980.675 2787.945 ;
        RECT 1966.200 2787.760 1980.675 2787.900 ;
        RECT 1980.385 2787.715 1980.675 2787.760 ;
        RECT 2181.405 2787.900 2181.695 2787.945 ;
        RECT 2252.245 2787.900 2252.535 2787.945 ;
        RECT 2181.405 2787.760 2252.535 2787.900 ;
        RECT 2181.405 2787.715 2181.695 2787.760 ;
        RECT 2252.245 2787.715 2252.535 2787.760 ;
        RECT 2252.690 2787.900 2253.010 2787.960 ;
        RECT 2421.970 2787.900 2422.290 2787.960 ;
        RECT 2252.690 2787.760 2422.290 2787.900 ;
        RECT 2252.690 2787.700 2253.010 2787.760 ;
        RECT 2421.970 2787.700 2422.290 2787.760 ;
        RECT 1780.360 2787.420 1828.340 2787.560 ;
        RECT 1738.425 2787.375 1738.715 2787.420 ;
        RECT 1980.385 2787.220 1980.675 2787.265 ;
        RECT 2028.225 2787.220 2028.515 2787.265 ;
        RECT 1980.385 2787.080 2028.515 2787.220 ;
        RECT 1980.385 2787.035 1980.675 2787.080 ;
        RECT 2028.225 2787.035 2028.515 2787.080 ;
        RECT 365.310 2731.800 365.630 2731.860 ;
        RECT 740.670 2731.800 740.990 2731.860 ;
        RECT 365.310 2731.660 740.990 2731.800 ;
        RECT 365.310 2731.600 365.630 2731.660 ;
        RECT 740.670 2731.600 740.990 2731.660 ;
        RECT 427.410 2731.460 427.730 2731.520 ;
        RECT 844.170 2731.460 844.490 2731.520 ;
        RECT 427.410 2731.320 844.490 2731.460 ;
        RECT 427.410 2731.260 427.730 2731.320 ;
        RECT 844.170 2731.260 844.490 2731.320 ;
        RECT 433.850 2731.120 434.170 2731.180 ;
        RECT 854.750 2731.120 855.070 2731.180 ;
        RECT 433.850 2730.980 855.070 2731.120 ;
        RECT 433.850 2730.920 434.170 2730.980 ;
        RECT 854.750 2730.920 855.070 2730.980 ;
        RECT 434.310 2730.780 434.630 2730.840 ;
        RECT 865.330 2730.780 865.650 2730.840 ;
        RECT 434.310 2730.640 865.650 2730.780 ;
        RECT 434.310 2730.580 434.630 2730.640 ;
        RECT 865.330 2730.580 865.650 2730.640 ;
        RECT 441.210 2730.440 441.530 2730.500 ;
        RECT 875.450 2730.440 875.770 2730.500 ;
        RECT 441.210 2730.300 875.770 2730.440 ;
        RECT 441.210 2730.240 441.530 2730.300 ;
        RECT 875.450 2730.240 875.770 2730.300 ;
        RECT 455.010 2730.100 455.330 2730.160 ;
        RECT 896.150 2730.100 896.470 2730.160 ;
        RECT 455.010 2729.960 896.470 2730.100 ;
        RECT 455.010 2729.900 455.330 2729.960 ;
        RECT 896.150 2729.900 896.470 2729.960 ;
        RECT 448.110 2729.760 448.430 2729.820 ;
        RECT 886.030 2729.760 886.350 2729.820 ;
        RECT 448.110 2729.620 886.350 2729.760 ;
        RECT 448.110 2729.560 448.430 2729.620 ;
        RECT 886.030 2729.560 886.350 2729.620 ;
        RECT 461.910 2729.420 462.230 2729.480 ;
        RECT 906.730 2729.420 907.050 2729.480 ;
        RECT 461.910 2729.280 907.050 2729.420 ;
        RECT 461.910 2729.220 462.230 2729.280 ;
        RECT 906.730 2729.220 907.050 2729.280 ;
        RECT 468.810 2729.080 469.130 2729.140 ;
        RECT 916.850 2729.080 917.170 2729.140 ;
        RECT 468.810 2728.940 917.170 2729.080 ;
        RECT 468.810 2728.880 469.130 2728.940 ;
        RECT 916.850 2728.880 917.170 2728.940 ;
        RECT 468.350 2728.740 468.670 2728.800 ;
        RECT 927.430 2728.740 927.750 2728.800 ;
        RECT 468.350 2728.600 927.750 2728.740 ;
        RECT 468.350 2728.540 468.670 2728.600 ;
        RECT 927.430 2728.540 927.750 2728.600 ;
        RECT 288.950 2725.340 289.270 2725.400 ;
        RECT 553.910 2725.340 554.230 2725.400 ;
        RECT 288.950 2725.200 554.230 2725.340 ;
        RECT 288.950 2725.140 289.270 2725.200 ;
        RECT 553.910 2725.140 554.230 2725.200 ;
        RECT 289.410 2725.000 289.730 2725.060 ;
        RECT 564.030 2725.000 564.350 2725.060 ;
        RECT 289.410 2724.860 564.350 2725.000 ;
        RECT 289.410 2724.800 289.730 2724.860 ;
        RECT 564.030 2724.800 564.350 2724.860 ;
        RECT 475.710 2724.660 476.030 2724.720 ;
        RECT 937.550 2724.660 937.870 2724.720 ;
        RECT 475.710 2724.520 937.870 2724.660 ;
        RECT 475.710 2724.460 476.030 2724.520 ;
        RECT 937.550 2724.460 937.870 2724.520 ;
        RECT 481.230 2724.320 481.550 2724.380 ;
        RECT 941.690 2724.320 942.010 2724.380 ;
        RECT 481.230 2724.180 942.010 2724.320 ;
        RECT 481.230 2724.120 481.550 2724.180 ;
        RECT 941.690 2724.120 942.010 2724.180 ;
        RECT 470.650 2723.980 470.970 2724.040 ;
        RECT 942.150 2723.980 942.470 2724.040 ;
        RECT 470.650 2723.840 942.470 2723.980 ;
        RECT 470.650 2723.780 470.970 2723.840 ;
        RECT 942.150 2723.780 942.470 2723.840 ;
        RECT 460.530 2723.640 460.850 2723.700 ;
        RECT 942.610 2723.640 942.930 2723.700 ;
        RECT 460.530 2723.500 942.930 2723.640 ;
        RECT 460.530 2723.440 460.850 2723.500 ;
        RECT 942.610 2723.440 942.930 2723.500 ;
        RECT 449.950 2723.300 450.270 2723.360 ;
        RECT 943.070 2723.300 943.390 2723.360 ;
        RECT 449.950 2723.160 943.390 2723.300 ;
        RECT 449.950 2723.100 450.270 2723.160 ;
        RECT 943.070 2723.100 943.390 2723.160 ;
        RECT 439.830 2722.960 440.150 2723.020 ;
        RECT 943.530 2722.960 943.850 2723.020 ;
        RECT 439.830 2722.820 943.850 2722.960 ;
        RECT 439.830 2722.760 440.150 2722.820 ;
        RECT 943.530 2722.760 943.850 2722.820 ;
        RECT 429.250 2722.620 429.570 2722.680 ;
        RECT 943.990 2722.620 944.310 2722.680 ;
        RECT 429.250 2722.480 944.310 2722.620 ;
        RECT 429.250 2722.420 429.570 2722.480 ;
        RECT 943.990 2722.420 944.310 2722.480 ;
        RECT 419.130 2722.280 419.450 2722.340 ;
        RECT 944.450 2722.280 944.770 2722.340 ;
        RECT 419.130 2722.140 944.770 2722.280 ;
        RECT 419.130 2722.080 419.450 2722.140 ;
        RECT 944.450 2722.080 944.770 2722.140 ;
        RECT 408.550 2721.940 408.870 2722.000 ;
        RECT 979.870 2721.940 980.190 2722.000 ;
        RECT 408.550 2721.800 980.190 2721.940 ;
        RECT 408.550 2721.740 408.870 2721.800 ;
        RECT 979.870 2721.740 980.190 2721.800 ;
        RECT 288.490 2721.600 288.810 2721.660 ;
        RECT 543.330 2721.600 543.650 2721.660 ;
        RECT 288.490 2721.460 543.650 2721.600 ;
        RECT 288.490 2721.400 288.810 2721.460 ;
        RECT 543.330 2721.400 543.650 2721.460 ;
        RECT 288.030 2721.260 288.350 2721.320 ;
        RECT 533.210 2721.260 533.530 2721.320 ;
        RECT 288.030 2721.120 533.530 2721.260 ;
        RECT 288.030 2721.060 288.350 2721.120 ;
        RECT 533.210 2721.060 533.530 2721.120 ;
        RECT 287.570 2720.920 287.890 2720.980 ;
        RECT 522.630 2720.920 522.950 2720.980 ;
        RECT 287.570 2720.780 522.950 2720.920 ;
        RECT 287.570 2720.720 287.890 2720.780 ;
        RECT 522.630 2720.720 522.950 2720.780 ;
        RECT 287.110 2720.580 287.430 2720.640 ;
        RECT 512.510 2720.580 512.830 2720.640 ;
        RECT 287.110 2720.440 512.830 2720.580 ;
        RECT 287.110 2720.380 287.430 2720.440 ;
        RECT 512.510 2720.380 512.830 2720.440 ;
        RECT 358.410 2718.540 358.730 2718.600 ;
        RECT 377.270 2718.540 377.590 2718.600 ;
        RECT 358.410 2718.400 377.590 2718.540 ;
        RECT 358.410 2718.340 358.730 2718.400 ;
        RECT 377.270 2718.340 377.590 2718.400 ;
        RECT 636.710 2718.540 637.030 2718.600 ;
        RECT 1045.190 2718.540 1045.510 2718.600 ;
        RECT 636.710 2718.400 1045.510 2718.540 ;
        RECT 636.710 2718.340 637.030 2718.400 ;
        RECT 1045.190 2718.340 1045.510 2718.400 ;
        RECT 1145.010 2718.540 1145.330 2718.600 ;
        RECT 1300.950 2718.540 1301.270 2718.600 ;
        RECT 1145.010 2718.400 1301.270 2718.540 ;
        RECT 1145.010 2718.340 1145.330 2718.400 ;
        RECT 1300.950 2718.340 1301.270 2718.400 ;
        RECT 616.010 2718.200 616.330 2718.260 ;
        RECT 1038.290 2718.200 1038.610 2718.260 ;
        RECT 616.010 2718.060 1038.610 2718.200 ;
        RECT 616.010 2718.000 616.330 2718.060 ;
        RECT 1038.290 2718.000 1038.610 2718.060 ;
        RECT 1138.110 2718.200 1138.430 2718.260 ;
        RECT 1290.370 2718.200 1290.690 2718.260 ;
        RECT 1138.110 2718.060 1290.690 2718.200 ;
        RECT 1138.110 2718.000 1138.430 2718.060 ;
        RECT 1290.370 2718.000 1290.690 2718.060 ;
        RECT 351.050 2717.860 351.370 2717.920 ;
        RECT 356.570 2717.860 356.890 2717.920 ;
        RECT 351.050 2717.720 356.890 2717.860 ;
        RECT 351.050 2717.660 351.370 2717.720 ;
        RECT 356.570 2717.660 356.890 2717.720 ;
        RECT 595.310 2717.860 595.630 2717.920 ;
        RECT 1024.490 2717.860 1024.810 2717.920 ;
        RECT 595.310 2717.720 1024.810 2717.860 ;
        RECT 595.310 2717.660 595.630 2717.720 ;
        RECT 1024.490 2717.660 1024.810 2717.720 ;
        RECT 1041.510 2717.860 1041.830 2717.920 ;
        RECT 1114.190 2717.860 1114.510 2717.920 ;
        RECT 1041.510 2717.720 1114.510 2717.860 ;
        RECT 1041.510 2717.660 1041.830 2717.720 ;
        RECT 1114.190 2717.660 1114.510 2717.720 ;
        RECT 1158.810 2717.860 1159.130 2717.920 ;
        RECT 1321.650 2717.860 1321.970 2717.920 ;
        RECT 1158.810 2717.720 1321.970 2717.860 ;
        RECT 1158.810 2717.660 1159.130 2717.720 ;
        RECT 1321.650 2717.660 1321.970 2717.720 ;
        RECT 574.610 2717.520 574.930 2717.580 ;
        RECT 1010.690 2717.520 1011.010 2717.580 ;
        RECT 574.610 2717.380 1011.010 2717.520 ;
        RECT 574.610 2717.320 574.930 2717.380 ;
        RECT 1010.690 2717.320 1011.010 2717.380 ;
        RECT 1048.410 2717.520 1048.730 2717.580 ;
        RECT 1124.310 2717.520 1124.630 2717.580 ;
        RECT 1048.410 2717.380 1124.630 2717.520 ;
        RECT 1048.410 2717.320 1048.730 2717.380 ;
        RECT 1124.310 2717.320 1124.630 2717.380 ;
        RECT 1151.910 2717.520 1152.230 2717.580 ;
        RECT 1311.070 2717.520 1311.390 2717.580 ;
        RECT 1151.910 2717.380 1311.390 2717.520 ;
        RECT 1151.910 2717.320 1152.230 2717.380 ;
        RECT 1311.070 2717.320 1311.390 2717.380 ;
        RECT 500.550 2717.180 500.870 2717.240 ;
        RECT 948.130 2717.180 948.450 2717.240 ;
        RECT 500.550 2717.040 948.450 2717.180 ;
        RECT 500.550 2716.980 500.870 2717.040 ;
        RECT 948.130 2716.980 948.450 2717.040 ;
        RECT 1055.310 2717.180 1055.630 2717.240 ;
        RECT 1134.890 2717.180 1135.210 2717.240 ;
        RECT 1055.310 2717.040 1135.210 2717.180 ;
        RECT 1055.310 2716.980 1055.630 2717.040 ;
        RECT 1134.890 2716.980 1135.210 2717.040 ;
        RECT 1165.710 2717.180 1166.030 2717.240 ;
        RECT 1332.230 2717.180 1332.550 2717.240 ;
        RECT 1165.710 2717.040 1332.550 2717.180 ;
        RECT 1165.710 2716.980 1166.030 2717.040 ;
        RECT 1332.230 2716.980 1332.550 2717.040 ;
        RECT 315.170 2716.840 315.490 2716.900 ;
        RECT 410.390 2716.840 410.710 2716.900 ;
        RECT 315.170 2716.700 410.710 2716.840 ;
        RECT 315.170 2716.640 315.490 2716.700 ;
        RECT 410.390 2716.640 410.710 2716.700 ;
        RECT 496.410 2716.840 496.730 2716.900 ;
        RECT 968.830 2716.840 969.150 2716.900 ;
        RECT 496.410 2716.700 969.150 2716.840 ;
        RECT 496.410 2716.640 496.730 2716.700 ;
        RECT 968.830 2716.640 969.150 2716.700 ;
        RECT 1062.210 2716.840 1062.530 2716.900 ;
        RECT 1155.590 2716.840 1155.910 2716.900 ;
        RECT 1062.210 2716.700 1155.910 2716.840 ;
        RECT 1062.210 2716.640 1062.530 2716.700 ;
        RECT 1155.590 2716.640 1155.910 2716.700 ;
        RECT 1165.250 2716.840 1165.570 2716.900 ;
        RECT 1342.350 2716.840 1342.670 2716.900 ;
        RECT 1165.250 2716.700 1342.670 2716.840 ;
        RECT 1165.250 2716.640 1165.570 2716.700 ;
        RECT 1342.350 2716.640 1342.670 2716.700 ;
        RECT 286.190 2716.500 286.510 2716.560 ;
        RECT 398.430 2716.500 398.750 2716.560 ;
        RECT 286.190 2716.360 398.750 2716.500 ;
        RECT 286.190 2716.300 286.510 2716.360 ;
        RECT 398.430 2716.300 398.750 2716.360 ;
        RECT 509.750 2716.500 510.070 2716.560 ;
        RECT 989.530 2716.500 989.850 2716.560 ;
        RECT 509.750 2716.360 989.850 2716.500 ;
        RECT 509.750 2716.300 510.070 2716.360 ;
        RECT 989.530 2716.300 989.850 2716.360 ;
        RECT 1076.010 2716.500 1076.330 2716.560 ;
        RECT 1176.290 2716.500 1176.610 2716.560 ;
        RECT 1076.010 2716.360 1176.610 2716.500 ;
        RECT 1076.010 2716.300 1076.330 2716.360 ;
        RECT 1176.290 2716.300 1176.610 2716.360 ;
        RECT 1179.510 2716.500 1179.830 2716.560 ;
        RECT 1363.050 2716.500 1363.370 2716.560 ;
        RECT 1179.510 2716.360 1363.370 2716.500 ;
        RECT 1179.510 2716.300 1179.830 2716.360 ;
        RECT 1363.050 2716.300 1363.370 2716.360 ;
        RECT 335.870 2716.160 336.190 2716.220 ;
        RECT 479.390 2716.160 479.710 2716.220 ;
        RECT 335.870 2716.020 479.710 2716.160 ;
        RECT 335.870 2715.960 336.190 2716.020 ;
        RECT 479.390 2715.960 479.710 2716.020 ;
        RECT 517.110 2716.160 517.430 2716.220 ;
        RECT 1010.230 2716.160 1010.550 2716.220 ;
        RECT 517.110 2716.020 1010.550 2716.160 ;
        RECT 517.110 2715.960 517.430 2716.020 ;
        RECT 1010.230 2715.960 1010.550 2716.020 ;
        RECT 1054.850 2716.160 1055.170 2716.220 ;
        RECT 1145.470 2716.160 1145.790 2716.220 ;
        RECT 1054.850 2716.020 1145.790 2716.160 ;
        RECT 1054.850 2715.960 1055.170 2716.020 ;
        RECT 1145.470 2715.960 1145.790 2716.020 ;
        RECT 1172.610 2716.160 1172.930 2716.220 ;
        RECT 1352.930 2716.160 1353.250 2716.220 ;
        RECT 1172.610 2716.020 1353.250 2716.160 ;
        RECT 1172.610 2715.960 1172.930 2716.020 ;
        RECT 1352.930 2715.960 1353.250 2716.020 ;
        RECT 337.710 2715.820 338.030 2715.880 ;
        RECT 491.810 2715.820 492.130 2715.880 ;
        RECT 337.710 2715.680 492.130 2715.820 ;
        RECT 337.710 2715.620 338.030 2715.680 ;
        RECT 491.810 2715.620 492.130 2715.680 ;
        RECT 530.910 2715.820 531.230 2715.880 ;
        RECT 1030.930 2715.820 1031.250 2715.880 ;
        RECT 530.910 2715.680 1031.250 2715.820 ;
        RECT 530.910 2715.620 531.230 2715.680 ;
        RECT 1030.930 2715.620 1031.250 2715.680 ;
        RECT 1069.110 2715.820 1069.430 2715.880 ;
        RECT 1166.170 2715.820 1166.490 2715.880 ;
        RECT 1069.110 2715.680 1166.490 2715.820 ;
        RECT 1069.110 2715.620 1069.430 2715.680 ;
        RECT 1166.170 2715.620 1166.490 2715.680 ;
        RECT 1186.410 2715.820 1186.730 2715.880 ;
        RECT 1373.630 2715.820 1373.950 2715.880 ;
        RECT 1186.410 2715.680 1373.950 2715.820 ;
        RECT 1186.410 2715.620 1186.730 2715.680 ;
        RECT 1373.630 2715.620 1373.950 2715.680 ;
        RECT 286.650 2715.480 286.970 2715.540 ;
        RECT 501.930 2715.480 502.250 2715.540 ;
        RECT 286.650 2715.340 502.250 2715.480 ;
        RECT 286.650 2715.280 286.970 2715.340 ;
        RECT 501.930 2715.280 502.250 2715.340 ;
        RECT 551.610 2715.480 551.930 2715.540 ;
        RECT 1062.210 2715.480 1062.530 2715.540 ;
        RECT 551.610 2715.340 1062.530 2715.480 ;
        RECT 551.610 2715.280 551.930 2715.340 ;
        RECT 1062.210 2715.280 1062.530 2715.340 ;
        RECT 1082.910 2715.480 1083.230 2715.540 ;
        RECT 1186.870 2715.480 1187.190 2715.540 ;
        RECT 1082.910 2715.340 1187.190 2715.480 ;
        RECT 1082.910 2715.280 1083.230 2715.340 ;
        RECT 1186.870 2715.280 1187.190 2715.340 ;
        RECT 1193.310 2715.480 1193.630 2715.540 ;
        RECT 1383.750 2715.480 1384.070 2715.540 ;
        RECT 1193.310 2715.340 1384.070 2715.480 ;
        RECT 1193.310 2715.280 1193.630 2715.340 ;
        RECT 1383.750 2715.280 1384.070 2715.340 ;
        RECT 387.850 2715.140 388.170 2715.200 ;
        RECT 927.890 2715.140 928.210 2715.200 ;
        RECT 387.850 2715.000 928.210 2715.140 ;
        RECT 387.850 2714.940 388.170 2715.000 ;
        RECT 927.890 2714.940 928.210 2715.000 ;
        RECT 1013.910 2715.140 1014.230 2715.200 ;
        RECT 1072.790 2715.140 1073.110 2715.200 ;
        RECT 1013.910 2715.000 1073.110 2715.140 ;
        RECT 1013.910 2714.940 1014.230 2715.000 ;
        RECT 1072.790 2714.940 1073.110 2715.000 ;
        RECT 1089.350 2715.140 1089.670 2715.200 ;
        RECT 1196.990 2715.140 1197.310 2715.200 ;
        RECT 1089.350 2715.000 1197.310 2715.140 ;
        RECT 1089.350 2714.940 1089.670 2715.000 ;
        RECT 1196.990 2714.940 1197.310 2715.000 ;
        RECT 1200.210 2715.140 1200.530 2715.200 ;
        RECT 1394.330 2715.140 1394.650 2715.200 ;
        RECT 1200.210 2715.000 1394.650 2715.140 ;
        RECT 1200.210 2714.940 1200.530 2715.000 ;
        RECT 1394.330 2714.940 1394.650 2715.000 ;
        RECT 325.750 2714.800 326.070 2714.860 ;
        RECT 700.190 2714.800 700.510 2714.860 ;
        RECT 325.750 2714.660 700.510 2714.800 ;
        RECT 325.750 2714.600 326.070 2714.660 ;
        RECT 700.190 2714.600 700.510 2714.660 ;
        RECT 872.690 2714.800 873.010 2714.860 ;
        RECT 1052.090 2714.800 1052.410 2714.860 ;
        RECT 872.690 2714.660 1052.410 2714.800 ;
        RECT 872.690 2714.600 873.010 2714.660 ;
        RECT 1052.090 2714.600 1052.410 2714.660 ;
        RECT 1103.610 2714.800 1103.930 2714.860 ;
        RECT 1131.210 2714.800 1131.530 2714.860 ;
        RECT 1280.250 2714.800 1280.570 2714.860 ;
        RECT 1103.610 2714.660 1104.300 2714.800 ;
        RECT 1103.610 2714.600 1103.930 2714.660 ;
        RECT 444.890 2714.460 445.210 2714.520 ;
        RECT 802.770 2714.460 803.090 2714.520 ;
        RECT 444.890 2714.320 803.090 2714.460 ;
        RECT 444.890 2714.260 445.210 2714.320 ;
        RECT 802.770 2714.260 803.090 2714.320 ;
        RECT 865.790 2714.460 866.110 2714.520 ;
        RECT 1041.510 2714.460 1041.830 2714.520 ;
        RECT 865.790 2714.320 1041.830 2714.460 ;
        RECT 865.790 2714.260 866.110 2714.320 ;
        RECT 1041.510 2714.260 1041.830 2714.320 ;
        RECT 351.510 2714.120 351.830 2714.180 ;
        RECT 367.150 2714.120 367.470 2714.180 ;
        RECT 351.510 2713.980 367.470 2714.120 ;
        RECT 351.510 2713.920 351.830 2713.980 ;
        RECT 367.150 2713.920 367.470 2713.980 ;
        RECT 465.590 2714.120 465.910 2714.180 ;
        RECT 823.470 2714.120 823.790 2714.180 ;
        RECT 465.590 2713.980 823.790 2714.120 ;
        RECT 465.590 2713.920 465.910 2713.980 ;
        RECT 823.470 2713.920 823.790 2713.980 ;
        RECT 858.890 2714.120 859.210 2714.180 ;
        RECT 1020.810 2714.120 1021.130 2714.180 ;
        RECT 858.890 2713.980 1021.130 2714.120 ;
        RECT 858.890 2713.920 859.210 2713.980 ;
        RECT 1020.810 2713.920 1021.130 2713.980 ;
        RECT 1034.610 2714.120 1034.930 2714.180 ;
        RECT 1103.610 2714.120 1103.930 2714.180 ;
        RECT 1034.610 2713.980 1103.930 2714.120 ;
        RECT 1034.610 2713.920 1034.930 2713.980 ;
        RECT 1103.610 2713.920 1103.930 2713.980 ;
        RECT 431.090 2713.780 431.410 2713.840 ;
        RECT 782.070 2713.780 782.390 2713.840 ;
        RECT 431.090 2713.640 782.390 2713.780 ;
        RECT 431.090 2713.580 431.410 2713.640 ;
        RECT 782.070 2713.580 782.390 2713.640 ;
        RECT 851.990 2713.780 852.310 2713.840 ;
        RECT 1000.110 2713.780 1000.430 2713.840 ;
        RECT 851.990 2713.640 1000.430 2713.780 ;
        RECT 851.990 2713.580 852.310 2713.640 ;
        RECT 1000.110 2713.580 1000.430 2713.640 ;
        RECT 1027.710 2713.780 1028.030 2713.840 ;
        RECT 1093.490 2713.780 1093.810 2713.840 ;
        RECT 1027.710 2713.640 1093.810 2713.780 ;
        RECT 1027.710 2713.580 1028.030 2713.640 ;
        RECT 1093.490 2713.580 1093.810 2713.640 ;
        RECT 424.190 2713.440 424.510 2713.500 ;
        RECT 761.370 2713.440 761.690 2713.500 ;
        RECT 424.190 2713.300 761.690 2713.440 ;
        RECT 424.190 2713.240 424.510 2713.300 ;
        RECT 761.370 2713.240 761.690 2713.300 ;
        RECT 845.090 2713.440 845.410 2713.500 ;
        RECT 979.410 2713.440 979.730 2713.500 ;
        RECT 845.090 2713.300 979.730 2713.440 ;
        RECT 845.090 2713.240 845.410 2713.300 ;
        RECT 979.410 2713.240 979.730 2713.300 ;
        RECT 1021.270 2713.440 1021.590 2713.500 ;
        RECT 1082.910 2713.440 1083.230 2713.500 ;
        RECT 1021.270 2713.300 1083.230 2713.440 ;
        RECT 1104.160 2713.440 1104.300 2714.660 ;
        RECT 1131.210 2714.660 1280.570 2714.800 ;
        RECT 1131.210 2714.600 1131.530 2714.660 ;
        RECT 1280.250 2714.600 1280.570 2714.660 ;
        RECT 1130.750 2714.460 1131.070 2714.520 ;
        RECT 1269.670 2714.460 1269.990 2714.520 ;
        RECT 1130.750 2714.320 1269.990 2714.460 ;
        RECT 1130.750 2714.260 1131.070 2714.320 ;
        RECT 1269.670 2714.260 1269.990 2714.320 ;
        RECT 1117.410 2714.120 1117.730 2714.180 ;
        RECT 1248.970 2714.120 1249.290 2714.180 ;
        RECT 1117.410 2713.980 1249.290 2714.120 ;
        RECT 1117.410 2713.920 1117.730 2713.980 ;
        RECT 1248.970 2713.920 1249.290 2713.980 ;
        RECT 1123.390 2713.780 1123.710 2713.840 ;
        RECT 1259.550 2713.780 1259.870 2713.840 ;
        RECT 1123.390 2713.640 1259.870 2713.780 ;
        RECT 1123.390 2713.580 1123.710 2713.640 ;
        RECT 1259.550 2713.580 1259.870 2713.640 ;
        RECT 1228.270 2713.440 1228.590 2713.500 ;
        RECT 1104.160 2713.300 1228.590 2713.440 ;
        RECT 1021.270 2713.240 1021.590 2713.300 ;
        RECT 1082.910 2713.240 1083.230 2713.300 ;
        RECT 1228.270 2713.240 1228.590 2713.300 ;
        RECT 541.490 2713.100 541.810 2713.160 ;
        RECT 730.090 2713.100 730.410 2713.160 ;
        RECT 541.490 2712.960 730.410 2713.100 ;
        RECT 541.490 2712.900 541.810 2712.960 ;
        RECT 730.090 2712.900 730.410 2712.960 ;
        RECT 838.190 2713.100 838.510 2713.160 ;
        RECT 958.710 2713.100 959.030 2713.160 ;
        RECT 838.190 2712.960 959.030 2713.100 ;
        RECT 838.190 2712.900 838.510 2712.960 ;
        RECT 958.710 2712.900 959.030 2712.960 ;
        RECT 1110.510 2713.100 1110.830 2713.160 ;
        RECT 1238.850 2713.100 1239.170 2713.160 ;
        RECT 1110.510 2712.960 1239.170 2713.100 ;
        RECT 1110.510 2712.900 1110.830 2712.960 ;
        RECT 1238.850 2712.900 1239.170 2712.960 ;
        RECT 534.590 2712.760 534.910 2712.820 ;
        RECT 709.390 2712.760 709.710 2712.820 ;
        RECT 534.590 2712.620 709.710 2712.760 ;
        RECT 534.590 2712.560 534.910 2712.620 ;
        RECT 709.390 2712.560 709.710 2712.620 ;
        RECT 1089.810 2712.760 1090.130 2712.820 ;
        RECT 1207.570 2712.760 1207.890 2712.820 ;
        RECT 1089.810 2712.620 1207.890 2712.760 ;
        RECT 1089.810 2712.560 1090.130 2712.620 ;
        RECT 1207.570 2712.560 1207.890 2712.620 ;
        RECT 520.790 2712.420 521.110 2712.480 ;
        RECT 688.690 2712.420 689.010 2712.480 ;
        RECT 520.790 2712.280 689.010 2712.420 ;
        RECT 520.790 2712.220 521.110 2712.280 ;
        RECT 688.690 2712.220 689.010 2712.280 ;
        RECT 1096.710 2712.420 1097.030 2712.480 ;
        RECT 1217.690 2712.420 1218.010 2712.480 ;
        RECT 1096.710 2712.280 1218.010 2712.420 ;
        RECT 1096.710 2712.220 1097.030 2712.280 ;
        RECT 1217.690 2712.220 1218.010 2712.280 ;
        RECT 500.090 2712.080 500.410 2712.140 ;
        RECT 657.410 2712.080 657.730 2712.140 ;
        RECT 500.090 2711.940 657.730 2712.080 ;
        RECT 500.090 2711.880 500.410 2711.940 ;
        RECT 657.410 2711.880 657.730 2711.940 ;
      LAYER met1 ;
        RECT 300.000 1607.860 1397.420 2689.320 ;
      LAYER met1 ;
        RECT 1410.430 2152.780 1410.750 2152.840 ;
        RECT 2307.890 2152.780 2308.210 2152.840 ;
        RECT 1410.430 2152.640 2308.210 2152.780 ;
        RECT 1410.430 2152.580 1410.750 2152.640 ;
        RECT 2307.890 2152.580 2308.210 2152.640 ;
        RECT 1414.110 2145.640 1414.430 2145.700 ;
        RECT 2301.450 2145.640 2301.770 2145.700 ;
        RECT 1414.110 2145.500 2301.770 2145.640 ;
        RECT 1414.110 2145.440 1414.430 2145.500 ;
        RECT 2301.450 2145.440 2301.770 2145.500 ;
        RECT 1414.110 2138.840 1414.430 2138.900 ;
        RECT 2266.950 2138.840 2267.270 2138.900 ;
        RECT 1414.110 2138.700 2267.270 2138.840 ;
        RECT 1414.110 2138.640 1414.430 2138.700 ;
        RECT 2266.950 2138.640 2267.270 2138.700 ;
        RECT 1413.650 2138.500 1413.970 2138.560 ;
        RECT 2252.690 2138.500 2253.010 2138.560 ;
        RECT 1413.650 2138.360 2253.010 2138.500 ;
        RECT 1413.650 2138.300 1413.970 2138.360 ;
        RECT 2252.690 2138.300 2253.010 2138.360 ;
        RECT 1410.430 2132.040 1410.750 2132.100 ;
        RECT 2245.790 2132.040 2246.110 2132.100 ;
        RECT 1410.430 2131.900 2246.110 2132.040 ;
        RECT 1410.430 2131.840 1410.750 2131.900 ;
        RECT 2245.790 2131.840 2246.110 2131.900 ;
        RECT 1414.110 2125.240 1414.430 2125.300 ;
        RECT 2238.890 2125.240 2239.210 2125.300 ;
        RECT 1414.110 2125.100 2239.210 2125.240 ;
        RECT 1414.110 2125.040 1414.430 2125.100 ;
        RECT 2238.890 2125.040 2239.210 2125.100 ;
        RECT 1414.110 2118.100 1414.430 2118.160 ;
        RECT 2231.990 2118.100 2232.310 2118.160 ;
        RECT 1414.110 2117.960 2232.310 2118.100 ;
        RECT 1414.110 2117.900 1414.430 2117.960 ;
        RECT 2231.990 2117.900 2232.310 2117.960 ;
        RECT 1410.430 2117.760 1410.750 2117.820 ;
        RECT 2218.190 2117.760 2218.510 2117.820 ;
        RECT 1410.430 2117.620 2218.510 2117.760 ;
        RECT 1410.430 2117.560 1410.750 2117.620 ;
        RECT 2218.190 2117.560 2218.510 2117.620 ;
        RECT 1414.110 2111.300 1414.430 2111.360 ;
        RECT 1797.750 2111.300 1798.070 2111.360 ;
        RECT 1414.110 2111.160 1798.070 2111.300 ;
        RECT 1414.110 2111.100 1414.430 2111.160 ;
        RECT 1797.750 2111.100 1798.070 2111.160 ;
        RECT 1414.110 2104.500 1414.430 2104.560 ;
        RECT 1797.290 2104.500 1797.610 2104.560 ;
        RECT 1414.110 2104.360 1797.610 2104.500 ;
        RECT 1414.110 2104.300 1414.430 2104.360 ;
        RECT 1797.290 2104.300 1797.610 2104.360 ;
        RECT 1414.110 2097.360 1414.430 2097.420 ;
        RECT 1790.390 2097.360 1790.710 2097.420 ;
        RECT 1414.110 2097.220 1790.710 2097.360 ;
        RECT 1414.110 2097.160 1414.430 2097.220 ;
        RECT 1790.390 2097.160 1790.710 2097.220 ;
        RECT 1410.430 2097.020 1410.750 2097.080 ;
        RECT 1762.790 2097.020 1763.110 2097.080 ;
        RECT 1410.430 2096.880 1763.110 2097.020 ;
        RECT 1410.430 2096.820 1410.750 2096.880 ;
        RECT 1762.790 2096.820 1763.110 2096.880 ;
        RECT 1409.510 2090.560 1409.830 2090.620 ;
        RECT 1783.490 2090.560 1783.810 2090.620 ;
        RECT 1409.510 2090.420 1783.810 2090.560 ;
        RECT 1409.510 2090.360 1409.830 2090.420 ;
        RECT 1783.490 2090.360 1783.810 2090.420 ;
        RECT 1425.610 2087.840 1425.930 2087.900 ;
        RECT 1593.970 2087.840 1594.290 2087.900 ;
        RECT 1425.610 2087.700 1594.290 2087.840 ;
        RECT 1425.610 2087.640 1425.930 2087.700 ;
        RECT 1593.970 2087.640 1594.290 2087.700 ;
        RECT 1422.390 2087.500 1422.710 2087.560 ;
        RECT 1617.890 2087.500 1618.210 2087.560 ;
        RECT 1422.390 2087.360 1618.210 2087.500 ;
        RECT 1422.390 2087.300 1422.710 2087.360 ;
        RECT 1617.890 2087.300 1618.210 2087.360 ;
        RECT 1416.870 2087.160 1417.190 2087.220 ;
        RECT 1645.490 2087.160 1645.810 2087.220 ;
        RECT 1416.870 2087.020 1645.810 2087.160 ;
        RECT 1416.870 2086.960 1417.190 2087.020 ;
        RECT 1645.490 2086.960 1645.810 2087.020 ;
        RECT 1414.110 2083.760 1414.430 2083.820 ;
        RECT 2366.770 2083.760 2367.090 2083.820 ;
        RECT 1414.110 2083.620 2367.090 2083.760 ;
        RECT 1414.110 2083.560 1414.430 2083.620 ;
        RECT 2366.770 2083.560 2367.090 2083.620 ;
        RECT 1436.650 2083.420 1436.970 2083.480 ;
        RECT 2263.270 2083.420 2263.590 2083.480 ;
        RECT 1436.650 2083.280 2263.590 2083.420 ;
        RECT 1436.650 2083.220 1436.970 2083.280 ;
        RECT 2263.270 2083.220 2263.590 2083.280 ;
        RECT 1436.190 2083.080 1436.510 2083.140 ;
        RECT 2263.730 2083.080 2264.050 2083.140 ;
        RECT 1436.190 2082.940 2264.050 2083.080 ;
        RECT 1436.190 2082.880 1436.510 2082.940 ;
        RECT 2263.730 2082.880 2264.050 2082.940 ;
        RECT 1412.730 2082.740 1413.050 2082.800 ;
        RECT 2266.490 2082.740 2266.810 2082.800 ;
        RECT 1412.730 2082.600 2266.810 2082.740 ;
        RECT 1412.730 2082.540 1413.050 2082.600 ;
        RECT 2266.490 2082.540 2266.810 2082.600 ;
        RECT 1412.270 2082.400 1412.590 2082.460 ;
        RECT 2270.170 2082.400 2270.490 2082.460 ;
        RECT 1412.270 2082.260 2270.490 2082.400 ;
        RECT 1412.270 2082.200 1412.590 2082.260 ;
        RECT 2270.170 2082.200 2270.490 2082.260 ;
        RECT 1435.730 2082.060 1436.050 2082.120 ;
        RECT 2305.130 2082.060 2305.450 2082.120 ;
        RECT 1435.730 2081.920 2305.450 2082.060 ;
        RECT 1435.730 2081.860 1436.050 2081.920 ;
        RECT 2305.130 2081.860 2305.450 2081.920 ;
        RECT 1421.930 2081.720 1422.250 2081.780 ;
        RECT 2297.770 2081.720 2298.090 2081.780 ;
        RECT 1421.930 2081.580 2298.090 2081.720 ;
        RECT 1421.930 2081.520 1422.250 2081.580 ;
        RECT 2297.770 2081.520 2298.090 2081.580 ;
        RECT 1414.570 2081.380 1414.890 2081.440 ;
        RECT 2318.470 2081.380 2318.790 2081.440 ;
        RECT 1414.570 2081.240 2318.790 2081.380 ;
        RECT 1414.570 2081.180 1414.890 2081.240 ;
        RECT 2318.470 2081.180 2318.790 2081.240 ;
        RECT 1409.510 2081.040 1409.830 2081.100 ;
        RECT 2325.370 2081.040 2325.690 2081.100 ;
        RECT 1409.510 2080.900 2325.690 2081.040 ;
        RECT 1409.510 2080.840 1409.830 2080.900 ;
        RECT 2325.370 2080.840 2325.690 2080.900 ;
        RECT 1408.590 2080.700 1408.910 2080.760 ;
        RECT 2332.270 2080.700 2332.590 2080.760 ;
        RECT 1408.590 2080.560 2332.590 2080.700 ;
        RECT 1408.590 2080.500 1408.910 2080.560 ;
        RECT 2332.270 2080.500 2332.590 2080.560 ;
        RECT 1409.050 2080.360 1409.370 2080.420 ;
        RECT 2339.630 2080.360 2339.950 2080.420 ;
        RECT 1409.050 2080.220 2339.950 2080.360 ;
        RECT 1409.050 2080.160 1409.370 2080.220 ;
        RECT 2339.630 2080.160 2339.950 2080.220 ;
        RECT 1440.330 2080.020 1440.650 2080.080 ;
        RECT 1662.970 2080.020 1663.290 2080.080 ;
        RECT 1440.330 2079.880 1663.290 2080.020 ;
        RECT 1440.330 2079.820 1440.650 2079.880 ;
        RECT 1662.970 2079.820 1663.290 2079.880 ;
        RECT 1439.410 2079.680 1439.730 2079.740 ;
        RECT 1656.070 2079.680 1656.390 2079.740 ;
        RECT 1439.410 2079.540 1656.390 2079.680 ;
        RECT 1439.410 2079.480 1439.730 2079.540 ;
        RECT 1656.070 2079.480 1656.390 2079.540 ;
        RECT 1417.330 2079.340 1417.650 2079.400 ;
        RECT 1624.790 2079.340 1625.110 2079.400 ;
        RECT 1417.330 2079.200 1625.110 2079.340 ;
        RECT 1417.330 2079.140 1417.650 2079.200 ;
        RECT 1624.790 2079.140 1625.110 2079.200 ;
        RECT 1494.150 2079.000 1494.470 2079.060 ;
        RECT 1631.690 2079.000 1632.010 2079.060 ;
        RECT 1494.150 2078.860 1632.010 2079.000 ;
        RECT 1494.150 2078.800 1494.470 2078.860 ;
        RECT 1631.690 2078.800 1632.010 2078.860 ;
        RECT 1414.110 2076.960 1414.430 2077.020 ;
        RECT 2359.870 2076.960 2360.190 2077.020 ;
        RECT 1414.110 2076.820 2360.190 2076.960 ;
        RECT 1414.110 2076.760 1414.430 2076.820 ;
        RECT 2359.870 2076.760 2360.190 2076.820 ;
        RECT 1413.650 2076.620 1413.970 2076.680 ;
        RECT 2352.970 2076.620 2353.290 2076.680 ;
        RECT 1413.650 2076.480 2353.290 2076.620 ;
        RECT 1413.650 2076.420 1413.970 2076.480 ;
        RECT 2352.970 2076.420 2353.290 2076.480 ;
        RECT 1429.750 2076.280 1430.070 2076.340 ;
        RECT 1745.770 2076.280 1746.090 2076.340 ;
        RECT 1429.750 2076.140 1746.090 2076.280 ;
        RECT 1429.750 2076.080 1430.070 2076.140 ;
        RECT 1745.770 2076.080 1746.090 2076.140 ;
        RECT 1440.790 2075.940 1441.110 2076.000 ;
        RECT 1760.490 2075.940 1760.810 2076.000 ;
        RECT 1440.790 2075.800 1760.810 2075.940 ;
        RECT 1440.790 2075.740 1441.110 2075.800 ;
        RECT 1760.490 2075.740 1760.810 2075.800 ;
        RECT 1428.830 2075.600 1429.150 2075.660 ;
        RECT 1752.670 2075.600 1752.990 2075.660 ;
        RECT 1428.830 2075.460 1752.990 2075.600 ;
        RECT 1428.830 2075.400 1429.150 2075.460 ;
        RECT 1752.670 2075.400 1752.990 2075.460 ;
        RECT 1441.250 2075.260 1441.570 2075.320 ;
        RECT 1766.470 2075.260 1766.790 2075.320 ;
        RECT 1441.250 2075.120 1766.790 2075.260 ;
        RECT 1441.250 2075.060 1441.570 2075.120 ;
        RECT 1766.470 2075.060 1766.790 2075.120 ;
        RECT 1441.710 2074.920 1442.030 2074.980 ;
        RECT 1773.830 2074.920 1774.150 2074.980 ;
        RECT 1441.710 2074.780 1774.150 2074.920 ;
        RECT 1441.710 2074.720 1442.030 2074.780 ;
        RECT 1773.830 2074.720 1774.150 2074.780 ;
        RECT 1428.370 2074.580 1428.690 2074.640 ;
        RECT 1760.030 2074.580 1760.350 2074.640 ;
        RECT 1428.370 2074.440 1760.350 2074.580 ;
        RECT 1428.370 2074.380 1428.690 2074.440 ;
        RECT 1760.030 2074.380 1760.350 2074.440 ;
        RECT 1438.030 2074.240 1438.350 2074.300 ;
        RECT 1780.270 2074.240 1780.590 2074.300 ;
        RECT 1438.030 2074.100 1780.590 2074.240 ;
        RECT 1438.030 2074.040 1438.350 2074.100 ;
        RECT 1780.270 2074.040 1780.590 2074.100 ;
        RECT 1437.570 2073.900 1437.890 2073.960 ;
        RECT 1787.170 2073.900 1787.490 2073.960 ;
        RECT 1437.570 2073.760 1787.490 2073.900 ;
        RECT 1437.570 2073.700 1437.890 2073.760 ;
        RECT 1787.170 2073.700 1787.490 2073.760 ;
        RECT 1437.110 2073.560 1437.430 2073.620 ;
        RECT 1794.530 2073.560 1794.850 2073.620 ;
        RECT 1437.110 2073.420 1794.850 2073.560 ;
        RECT 1437.110 2073.360 1437.430 2073.420 ;
        RECT 1794.530 2073.360 1794.850 2073.420 ;
        RECT 1430.210 2073.220 1430.530 2073.280 ;
        RECT 1738.870 2073.220 1739.190 2073.280 ;
        RECT 1430.210 2073.080 1739.190 2073.220 ;
        RECT 1430.210 2073.020 1430.530 2073.080 ;
        RECT 1738.870 2073.020 1739.190 2073.080 ;
        RECT 1439.870 2072.880 1440.190 2072.940 ;
        RECT 1649.170 2072.880 1649.490 2072.940 ;
        RECT 1439.870 2072.740 1649.490 2072.880 ;
        RECT 1439.870 2072.680 1440.190 2072.740 ;
        RECT 1649.170 2072.680 1649.490 2072.740 ;
        RECT 1432.510 2072.540 1432.830 2072.600 ;
        RECT 1621.570 2072.540 1621.890 2072.600 ;
        RECT 1432.510 2072.400 1621.890 2072.540 ;
        RECT 1432.510 2072.340 1432.830 2072.400 ;
        RECT 1621.570 2072.340 1621.890 2072.400 ;
        RECT 1494.610 2072.200 1494.930 2072.260 ;
        RECT 1649.630 2072.200 1649.950 2072.260 ;
        RECT 1494.610 2072.060 1649.950 2072.200 ;
        RECT 1494.610 2072.000 1494.930 2072.060 ;
        RECT 1649.630 2072.000 1649.950 2072.060 ;
        RECT 1414.110 2069.820 1414.430 2069.880 ;
        RECT 2346.070 2069.820 2346.390 2069.880 ;
        RECT 1414.110 2069.680 2346.390 2069.820 ;
        RECT 1414.110 2069.620 1414.430 2069.680 ;
        RECT 2346.070 2069.620 2346.390 2069.680 ;
        RECT 1433.430 2069.480 1433.750 2069.540 ;
        RECT 1684.130 2069.480 1684.450 2069.540 ;
        RECT 1433.430 2069.340 1684.450 2069.480 ;
        RECT 1433.430 2069.280 1433.750 2069.340 ;
        RECT 1684.130 2069.280 1684.450 2069.340 ;
        RECT 1434.350 2069.140 1434.670 2069.200 ;
        RECT 1697.470 2069.140 1697.790 2069.200 ;
        RECT 1434.350 2069.000 1697.790 2069.140 ;
        RECT 1434.350 2068.940 1434.670 2069.000 ;
        RECT 1697.470 2068.940 1697.790 2069.000 ;
        RECT 1416.410 2068.800 1416.730 2068.860 ;
        RECT 1683.670 2068.800 1683.990 2068.860 ;
        RECT 1416.410 2068.660 1683.990 2068.800 ;
        RECT 1416.410 2068.600 1416.730 2068.660 ;
        RECT 1683.670 2068.600 1683.990 2068.660 ;
        RECT 1415.950 2068.460 1416.270 2068.520 ;
        RECT 1690.570 2068.460 1690.890 2068.520 ;
        RECT 1415.950 2068.320 1690.890 2068.460 ;
        RECT 1415.950 2068.260 1416.270 2068.320 ;
        RECT 1690.570 2068.260 1690.890 2068.320 ;
        RECT 1434.810 2068.120 1435.130 2068.180 ;
        RECT 1711.270 2068.120 1711.590 2068.180 ;
        RECT 1434.810 2067.980 1711.590 2068.120 ;
        RECT 1434.810 2067.920 1435.130 2067.980 ;
        RECT 1711.270 2067.920 1711.590 2067.980 ;
        RECT 1430.670 2067.780 1430.990 2067.840 ;
        RECT 1718.170 2067.780 1718.490 2067.840 ;
        RECT 1430.670 2067.640 1718.490 2067.780 ;
        RECT 1430.670 2067.580 1430.990 2067.640 ;
        RECT 1718.170 2067.580 1718.490 2067.640 ;
        RECT 1415.490 2067.440 1415.810 2067.500 ;
        RECT 1704.370 2067.440 1704.690 2067.500 ;
        RECT 1415.490 2067.300 1704.690 2067.440 ;
        RECT 1415.490 2067.240 1415.810 2067.300 ;
        RECT 1704.370 2067.240 1704.690 2067.300 ;
        RECT 1431.130 2067.100 1431.450 2067.160 ;
        RECT 1725.070 2067.100 1725.390 2067.160 ;
        RECT 1431.130 2066.960 1725.390 2067.100 ;
        RECT 1431.130 2066.900 1431.450 2066.960 ;
        RECT 1725.070 2066.900 1725.390 2066.960 ;
        RECT 1429.290 2066.760 1429.610 2066.820 ;
        RECT 1731.970 2066.760 1732.290 2066.820 ;
        RECT 1429.290 2066.620 1732.290 2066.760 ;
        RECT 1429.290 2066.560 1429.610 2066.620 ;
        RECT 1731.970 2066.560 1732.290 2066.620 ;
        RECT 1415.030 2066.420 1415.350 2066.480 ;
        RECT 1718.630 2066.420 1718.950 2066.480 ;
        RECT 1415.030 2066.280 1718.950 2066.420 ;
        RECT 1415.030 2066.220 1415.350 2066.280 ;
        RECT 1718.630 2066.220 1718.950 2066.280 ;
        RECT 1433.890 2066.080 1434.210 2066.140 ;
        RECT 1676.770 2066.080 1677.090 2066.140 ;
        RECT 1433.890 2065.940 1677.090 2066.080 ;
        RECT 1433.890 2065.880 1434.210 2065.940 ;
        RECT 1676.770 2065.880 1677.090 2065.940 ;
        RECT 1432.970 2065.740 1433.290 2065.800 ;
        RECT 1669.870 2065.740 1670.190 2065.800 ;
        RECT 1432.970 2065.600 1670.190 2065.740 ;
        RECT 1432.970 2065.540 1433.290 2065.600 ;
        RECT 1669.870 2065.540 1670.190 2065.600 ;
        RECT 1432.050 2065.400 1432.370 2065.460 ;
        RECT 1607.770 2065.400 1608.090 2065.460 ;
        RECT 1432.050 2065.260 1608.090 2065.400 ;
        RECT 1432.050 2065.200 1432.370 2065.260 ;
        RECT 1607.770 2065.200 1608.090 2065.260 ;
        RECT 1466.090 2065.060 1466.410 2065.120 ;
        RECT 1614.670 2065.060 1614.990 2065.120 ;
        RECT 1466.090 2064.920 1614.990 2065.060 ;
        RECT 1466.090 2064.860 1466.410 2064.920 ;
        RECT 1614.670 2064.860 1614.990 2064.920 ;
        RECT 1412.270 2063.360 1412.590 2063.420 ;
        RECT 1413.650 2063.360 1413.970 2063.420 ;
        RECT 1412.270 2063.220 1413.970 2063.360 ;
        RECT 1412.270 2063.160 1412.590 2063.220 ;
        RECT 1413.650 2063.160 1413.970 2063.220 ;
        RECT 1414.110 2063.020 1414.430 2063.080 ;
        RECT 2339.170 2063.020 2339.490 2063.080 ;
        RECT 1414.110 2062.880 2339.490 2063.020 ;
        RECT 1414.110 2062.820 1414.430 2062.880 ;
        RECT 2339.170 2062.820 2339.490 2062.880 ;
        RECT 1426.990 2062.680 1427.310 2062.740 ;
        RECT 2193.350 2062.680 2193.670 2062.740 ;
        RECT 1426.990 2062.540 2193.670 2062.680 ;
        RECT 1426.990 2062.480 1427.310 2062.540 ;
        RECT 2193.350 2062.480 2193.670 2062.540 ;
        RECT 1423.310 2062.340 1423.630 2062.400 ;
        RECT 2190.590 2062.340 2190.910 2062.400 ;
        RECT 1423.310 2062.200 2190.910 2062.340 ;
        RECT 1423.310 2062.140 1423.630 2062.200 ;
        RECT 2190.590 2062.140 2190.910 2062.200 ;
        RECT 1423.770 2062.000 1424.090 2062.060 ;
        RECT 2191.510 2062.000 2191.830 2062.060 ;
        RECT 1423.770 2061.860 2191.830 2062.000 ;
        RECT 1423.770 2061.800 1424.090 2061.860 ;
        RECT 2191.510 2061.800 2191.830 2061.860 ;
        RECT 1424.230 2061.660 1424.550 2061.720 ;
        RECT 2191.970 2061.660 2192.290 2061.720 ;
        RECT 1424.230 2061.520 2192.290 2061.660 ;
        RECT 1424.230 2061.460 1424.550 2061.520 ;
        RECT 2191.970 2061.460 2192.290 2061.520 ;
        RECT 1422.850 2061.320 1423.170 2061.380 ;
        RECT 2191.050 2061.320 2191.370 2061.380 ;
        RECT 1422.850 2061.180 2191.370 2061.320 ;
        RECT 1422.850 2061.120 1423.170 2061.180 ;
        RECT 2191.050 2061.120 2191.370 2061.180 ;
        RECT 1426.530 2060.980 1426.850 2061.040 ;
        RECT 2228.770 2060.980 2229.090 2061.040 ;
        RECT 1426.530 2060.840 2229.090 2060.980 ;
        RECT 1426.530 2060.780 1426.850 2060.840 ;
        RECT 2228.770 2060.780 2229.090 2060.840 ;
        RECT 1426.070 2060.640 1426.390 2060.700 ;
        RECT 2256.370 2060.640 2256.690 2060.700 ;
        RECT 1426.070 2060.500 2256.690 2060.640 ;
        RECT 1426.070 2060.440 1426.390 2060.500 ;
        RECT 2256.370 2060.440 2256.690 2060.500 ;
        RECT 1409.970 2060.300 1410.290 2060.360 ;
        RECT 2242.570 2060.300 2242.890 2060.360 ;
        RECT 1409.970 2060.160 2242.890 2060.300 ;
        RECT 1409.970 2060.100 1410.290 2060.160 ;
        RECT 2242.570 2060.100 2242.890 2060.160 ;
        RECT 1438.950 2059.960 1439.270 2060.020 ;
        RECT 2300.990 2059.960 2301.310 2060.020 ;
        RECT 1438.950 2059.820 2301.310 2059.960 ;
        RECT 1438.950 2059.760 1439.270 2059.820 ;
        RECT 2300.990 2059.760 2301.310 2059.820 ;
        RECT 1421.010 2059.620 1421.330 2059.680 ;
        RECT 2294.090 2059.620 2294.410 2059.680 ;
        RECT 1421.010 2059.480 2294.410 2059.620 ;
        RECT 1421.010 2059.420 1421.330 2059.480 ;
        RECT 2294.090 2059.420 2294.410 2059.480 ;
        RECT 1427.450 2059.280 1427.770 2059.340 ;
        RECT 2192.430 2059.280 2192.750 2059.340 ;
        RECT 1427.450 2059.140 2192.750 2059.280 ;
        RECT 1427.450 2059.080 1427.770 2059.140 ;
        RECT 2192.430 2059.080 2192.750 2059.140 ;
        RECT 1427.910 2058.940 1428.230 2059.000 ;
        RECT 2192.890 2058.940 2193.210 2059.000 ;
        RECT 1427.910 2058.800 2193.210 2058.940 ;
        RECT 1427.910 2058.740 1428.230 2058.800 ;
        RECT 2192.890 2058.740 2193.210 2058.800 ;
        RECT 1460.110 2058.600 1460.430 2058.660 ;
        RECT 1601.330 2058.600 1601.650 2058.660 ;
        RECT 1460.110 2058.460 1601.650 2058.600 ;
        RECT 1460.110 2058.400 1460.430 2058.460 ;
        RECT 1601.330 2058.400 1601.650 2058.460 ;
        RECT 1493.690 2058.260 1494.010 2058.320 ;
        RECT 1580.170 2058.260 1580.490 2058.320 ;
        RECT 1493.690 2058.120 1580.490 2058.260 ;
        RECT 1493.690 2058.060 1494.010 2058.120 ;
        RECT 1580.170 2058.060 1580.490 2058.120 ;
        RECT 1409.065 2056.560 1409.355 2056.605 ;
        RECT 1409.970 2056.560 1410.290 2056.620 ;
        RECT 1409.065 2056.420 1410.290 2056.560 ;
        RECT 1409.065 2056.375 1409.355 2056.420 ;
        RECT 1409.970 2056.360 1410.290 2056.420 ;
        RECT 1409.970 2054.520 1410.290 2054.580 ;
        RECT 2273.390 2054.520 2273.710 2054.580 ;
        RECT 1409.970 2054.380 2273.710 2054.520 ;
        RECT 1409.970 2054.320 1410.290 2054.380 ;
        RECT 2273.390 2054.320 2273.710 2054.380 ;
        RECT 1412.270 2054.180 1412.590 2054.240 ;
        RECT 2277.070 2054.180 2277.390 2054.240 ;
        RECT 1412.270 2054.040 2277.390 2054.180 ;
        RECT 1412.270 2053.980 1412.590 2054.040 ;
        RECT 2277.070 2053.980 2277.390 2054.040 ;
        RECT 1414.110 2053.840 1414.430 2053.900 ;
        RECT 2283.970 2053.840 2284.290 2053.900 ;
        RECT 1414.110 2053.700 2284.290 2053.840 ;
        RECT 1414.110 2053.640 1414.430 2053.700 ;
        RECT 2283.970 2053.640 2284.290 2053.700 ;
        RECT 1410.430 2053.500 1410.750 2053.560 ;
        RECT 2290.870 2053.500 2291.190 2053.560 ;
        RECT 1410.430 2053.360 2291.190 2053.500 ;
        RECT 1410.430 2053.300 1410.750 2053.360 ;
        RECT 2290.870 2053.300 2291.190 2053.360 ;
        RECT 1413.190 2053.160 1413.510 2053.220 ;
        RECT 2304.670 2053.160 2304.990 2053.220 ;
        RECT 1413.190 2053.020 2304.990 2053.160 ;
        RECT 1413.190 2052.960 1413.510 2053.020 ;
        RECT 2304.670 2052.960 2304.990 2053.020 ;
        RECT 1409.510 2052.820 1409.830 2052.880 ;
        RECT 2311.570 2052.820 2311.890 2052.880 ;
        RECT 1409.510 2052.680 2311.890 2052.820 ;
        RECT 1409.510 2052.620 1409.830 2052.680 ;
        RECT 2311.570 2052.620 2311.890 2052.680 ;
        RECT 1409.050 2046.020 1409.370 2046.080 ;
        RECT 1408.855 2045.880 1409.370 2046.020 ;
        RECT 1409.050 2045.820 1409.370 2045.880 ;
        RECT 1409.510 2034.460 1409.830 2034.520 ;
        RECT 1414.110 2034.460 1414.430 2034.520 ;
        RECT 1409.510 2034.320 1414.430 2034.460 ;
        RECT 1409.510 2034.260 1409.830 2034.320 ;
        RECT 1414.110 2034.260 1414.430 2034.320 ;
        RECT 1414.110 2029.020 1414.430 2029.080 ;
        RECT 1435.730 2029.020 1436.050 2029.080 ;
        RECT 1414.110 2028.880 1436.050 2029.020 ;
        RECT 1414.110 2028.820 1414.430 2028.880 ;
        RECT 1435.730 2028.820 1436.050 2028.880 ;
        RECT 1412.270 2028.340 1412.590 2028.400 ;
        RECT 1414.110 2028.340 1414.430 2028.400 ;
        RECT 1412.270 2028.200 1414.430 2028.340 ;
        RECT 1412.270 2028.140 1412.590 2028.200 ;
        RECT 1414.110 2028.140 1414.430 2028.200 ;
        RECT 1409.050 2027.660 1409.370 2027.720 ;
        RECT 1412.270 2027.660 1412.590 2027.720 ;
        RECT 1409.050 2027.520 1412.590 2027.660 ;
        RECT 1409.050 2027.460 1409.370 2027.520 ;
        RECT 1412.270 2027.460 1412.590 2027.520 ;
        RECT 1409.970 2025.620 1410.290 2025.680 ;
        RECT 1413.190 2025.620 1413.510 2025.680 ;
        RECT 1409.970 2025.480 1413.510 2025.620 ;
        RECT 1409.970 2025.420 1410.290 2025.480 ;
        RECT 1413.190 2025.420 1413.510 2025.480 ;
        RECT 1409.050 2021.540 1409.370 2021.600 ;
        RECT 1421.930 2021.540 1422.250 2021.600 ;
        RECT 1409.050 2021.400 1422.250 2021.540 ;
        RECT 1409.050 2021.340 1409.370 2021.400 ;
        RECT 1421.930 2021.340 1422.250 2021.400 ;
        RECT 1413.190 2014.740 1413.510 2014.800 ;
        RECT 1414.570 2014.740 1414.890 2014.800 ;
        RECT 1413.190 2014.600 1414.890 2014.740 ;
        RECT 1413.190 2014.540 1413.510 2014.600 ;
        RECT 1414.570 2014.540 1414.890 2014.600 ;
        RECT 1414.110 1996.040 1414.430 1996.100 ;
        RECT 1436.190 1996.040 1436.510 1996.100 ;
        RECT 1414.110 1995.900 1436.510 1996.040 ;
        RECT 1414.110 1995.840 1414.430 1995.900 ;
        RECT 1436.190 1995.840 1436.510 1995.900 ;
        RECT 1414.110 1989.580 1414.430 1989.640 ;
        RECT 1436.650 1989.580 1436.970 1989.640 ;
        RECT 1414.110 1989.440 1436.970 1989.580 ;
        RECT 1414.110 1989.380 1414.430 1989.440 ;
        RECT 1436.650 1989.380 1436.970 1989.440 ;
        RECT 1414.110 1984.480 1414.430 1984.540 ;
        RECT 1437.110 1984.480 1437.430 1984.540 ;
        RECT 1414.110 1984.340 1437.430 1984.480 ;
        RECT 1414.110 1984.280 1414.430 1984.340 ;
        RECT 1437.110 1984.280 1437.430 1984.340 ;
        RECT 1414.110 1981.420 1414.430 1981.480 ;
        RECT 1437.570 1981.420 1437.890 1981.480 ;
        RECT 1414.110 1981.280 1437.890 1981.420 ;
        RECT 1414.110 1981.220 1414.430 1981.280 ;
        RECT 1437.570 1981.220 1437.890 1981.280 ;
        RECT 1414.110 1973.940 1414.430 1974.000 ;
        RECT 1438.030 1973.940 1438.350 1974.000 ;
        RECT 1414.110 1973.800 1438.350 1973.940 ;
        RECT 1414.110 1973.740 1414.430 1973.800 ;
        RECT 1438.030 1973.740 1438.350 1973.800 ;
        RECT 1414.110 1969.520 1414.430 1969.580 ;
        RECT 1441.710 1969.520 1442.030 1969.580 ;
        RECT 1414.110 1969.380 1442.030 1969.520 ;
        RECT 1414.110 1969.320 1414.430 1969.380 ;
        RECT 1441.710 1969.320 1442.030 1969.380 ;
        RECT 1409.510 1962.380 1409.830 1962.440 ;
        RECT 1441.250 1962.380 1441.570 1962.440 ;
        RECT 1409.510 1962.240 1441.570 1962.380 ;
        RECT 1409.510 1962.180 1409.830 1962.240 ;
        RECT 1441.250 1962.180 1441.570 1962.240 ;
        RECT 1414.110 1961.700 1414.430 1961.760 ;
        RECT 1440.790 1961.700 1441.110 1961.760 ;
        RECT 1414.110 1961.560 1441.110 1961.700 ;
        RECT 1414.110 1961.500 1414.430 1961.560 ;
        RECT 1440.790 1961.500 1441.110 1961.560 ;
        RECT 1410.430 1956.600 1410.750 1956.660 ;
        RECT 1428.370 1956.600 1428.690 1956.660 ;
        RECT 1410.430 1956.460 1428.690 1956.600 ;
        RECT 1410.430 1956.400 1410.750 1956.460 ;
        RECT 1428.370 1956.400 1428.690 1956.460 ;
        RECT 1413.650 1951.500 1413.970 1951.560 ;
        RECT 1428.830 1951.500 1429.150 1951.560 ;
        RECT 1413.650 1951.360 1429.150 1951.500 ;
        RECT 1413.650 1951.300 1413.970 1951.360 ;
        RECT 1428.830 1951.300 1429.150 1951.360 ;
        RECT 1413.650 1945.380 1413.970 1945.440 ;
        RECT 1429.750 1945.380 1430.070 1945.440 ;
        RECT 1413.650 1945.240 1430.070 1945.380 ;
        RECT 1413.650 1945.180 1413.970 1945.240 ;
        RECT 1429.750 1945.180 1430.070 1945.240 ;
        RECT 1413.650 1943.000 1413.970 1943.060 ;
        RECT 1430.210 1943.000 1430.530 1943.060 ;
        RECT 1413.650 1942.860 1430.530 1943.000 ;
        RECT 1413.650 1942.800 1413.970 1942.860 ;
        RECT 1430.210 1942.800 1430.530 1942.860 ;
        RECT 1413.650 1936.540 1413.970 1936.600 ;
        RECT 1429.290 1936.540 1429.610 1936.600 ;
        RECT 1413.650 1936.400 1429.610 1936.540 ;
        RECT 1413.650 1936.340 1413.970 1936.400 ;
        RECT 1429.290 1936.340 1429.610 1936.400 ;
        RECT 1413.650 1930.420 1413.970 1930.480 ;
        RECT 1431.130 1930.420 1431.450 1930.480 ;
        RECT 1413.650 1930.280 1431.450 1930.420 ;
        RECT 1413.650 1930.220 1413.970 1930.280 ;
        RECT 1431.130 1930.220 1431.450 1930.280 ;
        RECT 1413.650 1926.680 1413.970 1926.740 ;
        RECT 1430.670 1926.680 1430.990 1926.740 ;
        RECT 1413.650 1926.540 1430.990 1926.680 ;
        RECT 1413.650 1926.480 1413.970 1926.540 ;
        RECT 1430.670 1926.480 1430.990 1926.540 ;
        RECT 1414.110 1915.460 1414.430 1915.520 ;
        RECT 1434.810 1915.460 1435.130 1915.520 ;
        RECT 1414.110 1915.320 1435.130 1915.460 ;
        RECT 1414.110 1915.260 1414.430 1915.320 ;
        RECT 1434.810 1915.260 1435.130 1915.320 ;
        RECT 1414.110 1906.620 1414.430 1906.680 ;
        RECT 1434.350 1906.620 1434.670 1906.680 ;
        RECT 1414.110 1906.480 1434.670 1906.620 ;
        RECT 1414.110 1906.420 1414.430 1906.480 ;
        RECT 1434.350 1906.420 1434.670 1906.480 ;
        RECT 1408.590 1895.400 1408.910 1895.460 ;
        RECT 1416.410 1895.400 1416.730 1895.460 ;
        RECT 1408.590 1895.260 1416.730 1895.400 ;
        RECT 1408.590 1895.200 1408.910 1895.260 ;
        RECT 1416.410 1895.200 1416.730 1895.260 ;
        RECT 1414.110 1890.300 1414.430 1890.360 ;
        RECT 1433.430 1890.300 1433.750 1890.360 ;
        RECT 1414.110 1890.160 1433.750 1890.300 ;
        RECT 1414.110 1890.100 1414.430 1890.160 ;
        RECT 1433.430 1890.100 1433.750 1890.160 ;
        RECT 1414.110 1885.880 1414.430 1885.940 ;
        RECT 1433.890 1885.880 1434.210 1885.940 ;
        RECT 1414.110 1885.740 1434.210 1885.880 ;
        RECT 1414.110 1885.680 1414.430 1885.740 ;
        RECT 1433.890 1885.680 1434.210 1885.740 ;
        RECT 1414.110 1881.800 1414.430 1881.860 ;
        RECT 1432.970 1881.800 1433.290 1881.860 ;
        RECT 1414.110 1881.660 1433.290 1881.800 ;
        RECT 1414.110 1881.600 1414.430 1881.660 ;
        RECT 1432.970 1881.600 1433.290 1881.660 ;
        RECT 1414.110 1872.620 1414.430 1872.680 ;
        RECT 1440.330 1872.620 1440.650 1872.680 ;
        RECT 1414.110 1872.480 1440.650 1872.620 ;
        RECT 1414.110 1872.420 1414.430 1872.480 ;
        RECT 1440.330 1872.420 1440.650 1872.480 ;
        RECT 1410.430 1869.900 1410.750 1869.960 ;
        RECT 1413.190 1869.900 1413.510 1869.960 ;
        RECT 1410.430 1869.760 1413.510 1869.900 ;
        RECT 1410.430 1869.700 1410.750 1869.760 ;
        RECT 1413.190 1869.700 1413.510 1869.760 ;
        RECT 1413.650 1869.900 1413.970 1869.960 ;
        RECT 1494.610 1869.900 1494.930 1869.960 ;
        RECT 1413.650 1869.760 1494.930 1869.900 ;
        RECT 1413.650 1869.700 1413.970 1869.760 ;
        RECT 1494.610 1869.700 1494.930 1869.760 ;
        RECT 1414.110 1865.820 1414.430 1865.880 ;
        RECT 1439.410 1865.820 1439.730 1865.880 ;
        RECT 1414.110 1865.680 1439.730 1865.820 ;
        RECT 1414.110 1865.620 1414.430 1865.680 ;
        RECT 1439.410 1865.620 1439.730 1865.680 ;
        RECT 1414.110 1858.340 1414.430 1858.400 ;
        RECT 1439.870 1858.340 1440.190 1858.400 ;
        RECT 1414.110 1858.200 1440.190 1858.340 ;
        RECT 1414.110 1858.140 1414.430 1858.200 ;
        RECT 1439.870 1858.140 1440.190 1858.200 ;
        RECT 1414.110 1855.960 1414.430 1856.020 ;
        RECT 1549.810 1855.960 1550.130 1856.020 ;
        RECT 1414.110 1855.820 1550.130 1855.960 ;
        RECT 1414.110 1855.760 1414.430 1855.820 ;
        RECT 1549.810 1855.760 1550.130 1855.820 ;
        RECT 1413.650 1855.620 1413.970 1855.680 ;
        RECT 1549.350 1855.620 1549.670 1855.680 ;
        RECT 1413.650 1855.480 1549.670 1855.620 ;
        RECT 1413.650 1855.420 1413.970 1855.480 ;
        RECT 1549.350 1855.420 1549.670 1855.480 ;
        RECT 1414.110 1849.160 1414.430 1849.220 ;
        RECT 1548.890 1849.160 1549.210 1849.220 ;
        RECT 1414.110 1849.020 1549.210 1849.160 ;
        RECT 1414.110 1848.960 1414.430 1849.020 ;
        RECT 1548.890 1848.960 1549.210 1849.020 ;
        RECT 1414.110 1841.000 1414.430 1841.060 ;
        RECT 1432.510 1841.000 1432.830 1841.060 ;
        RECT 1414.110 1840.860 1432.830 1841.000 ;
        RECT 1414.110 1840.800 1414.430 1840.860 ;
        RECT 1432.510 1840.800 1432.830 1840.860 ;
        RECT 1414.110 1835.220 1414.430 1835.280 ;
        RECT 1466.090 1835.220 1466.410 1835.280 ;
        RECT 1414.110 1835.080 1466.410 1835.220 ;
        RECT 1414.110 1835.020 1414.430 1835.080 ;
        RECT 1466.090 1835.020 1466.410 1835.080 ;
        RECT 1414.110 1831.140 1414.430 1831.200 ;
        RECT 1432.050 1831.140 1432.370 1831.200 ;
        RECT 1414.110 1831.000 1432.370 1831.140 ;
        RECT 1414.110 1830.940 1414.430 1831.000 ;
        RECT 1432.050 1830.940 1432.370 1831.000 ;
        RECT 1408.590 1827.060 1408.910 1827.120 ;
        RECT 1420.550 1827.060 1420.870 1827.120 ;
        RECT 1408.590 1826.920 1420.870 1827.060 ;
        RECT 1408.590 1826.860 1408.910 1826.920 ;
        RECT 1420.550 1826.860 1420.870 1826.920 ;
        RECT 1410.430 1821.960 1410.750 1822.020 ;
        RECT 1413.190 1821.960 1413.510 1822.020 ;
        RECT 1410.430 1821.820 1413.510 1821.960 ;
        RECT 1410.430 1821.760 1410.750 1821.820 ;
        RECT 1413.190 1821.760 1413.510 1821.820 ;
        RECT 1408.590 1819.580 1408.910 1819.640 ;
        RECT 1416.870 1819.580 1417.190 1819.640 ;
        RECT 1408.590 1819.440 1417.190 1819.580 ;
        RECT 1408.590 1819.380 1408.910 1819.440 ;
        RECT 1416.870 1819.380 1417.190 1819.440 ;
        RECT 1408.590 1814.140 1408.910 1814.200 ;
        RECT 1419.630 1814.140 1419.950 1814.200 ;
        RECT 1408.590 1814.000 1419.950 1814.140 ;
        RECT 1408.590 1813.940 1408.910 1814.000 ;
        RECT 1419.630 1813.940 1419.950 1814.000 ;
        RECT 1408.590 1809.380 1408.910 1809.440 ;
        RECT 1420.090 1809.380 1420.410 1809.440 ;
        RECT 1408.590 1809.240 1420.410 1809.380 ;
        RECT 1408.590 1809.180 1408.910 1809.240 ;
        RECT 1420.090 1809.180 1420.410 1809.240 ;
        RECT 1414.110 1807.680 1414.430 1807.740 ;
        RECT 1494.150 1807.680 1494.470 1807.740 ;
        RECT 1414.110 1807.540 1494.470 1807.680 ;
        RECT 1414.110 1807.480 1414.430 1807.540 ;
        RECT 1494.150 1807.480 1494.470 1807.540 ;
        RECT 1409.050 1799.860 1409.370 1799.920 ;
        RECT 1422.390 1799.860 1422.710 1799.920 ;
        RECT 1409.050 1799.720 1422.710 1799.860 ;
        RECT 1409.050 1799.660 1409.370 1799.720 ;
        RECT 1422.390 1799.660 1422.710 1799.720 ;
        RECT 1408.590 1799.180 1408.910 1799.240 ;
        RECT 1417.330 1799.180 1417.650 1799.240 ;
        RECT 1408.590 1799.040 1417.650 1799.180 ;
        RECT 1408.590 1798.980 1408.910 1799.040 ;
        RECT 1417.330 1798.980 1417.650 1799.040 ;
        RECT 1414.110 1783.200 1414.430 1783.260 ;
        RECT 1438.950 1783.200 1439.270 1783.260 ;
        RECT 1414.110 1783.060 1439.270 1783.200 ;
        RECT 1414.110 1783.000 1414.430 1783.060 ;
        RECT 1438.950 1783.000 1439.270 1783.060 ;
        RECT 1408.590 1778.780 1408.910 1778.840 ;
        RECT 1419.170 1778.780 1419.490 1778.840 ;
        RECT 1408.590 1778.640 1419.490 1778.780 ;
        RECT 1408.590 1778.580 1408.910 1778.640 ;
        RECT 1419.170 1778.580 1419.490 1778.640 ;
        RECT 1408.590 1778.100 1408.910 1778.160 ;
        RECT 1421.010 1778.100 1421.330 1778.160 ;
        RECT 1408.590 1777.960 1421.330 1778.100 ;
        RECT 1408.590 1777.900 1408.910 1777.960 ;
        RECT 1421.010 1777.900 1421.330 1777.960 ;
        RECT 1408.590 1769.600 1408.910 1769.660 ;
        RECT 1418.710 1769.600 1419.030 1769.660 ;
        RECT 1408.590 1769.460 1419.030 1769.600 ;
        RECT 1408.590 1769.400 1408.910 1769.460 ;
        RECT 1418.710 1769.400 1419.030 1769.460 ;
        RECT 1408.590 1765.180 1408.910 1765.240 ;
        RECT 1418.250 1765.180 1418.570 1765.240 ;
        RECT 1408.590 1765.040 1418.570 1765.180 ;
        RECT 1408.590 1764.980 1408.910 1765.040 ;
        RECT 1418.250 1764.980 1418.570 1765.040 ;
        RECT 1408.590 1756.680 1408.910 1756.740 ;
        RECT 1417.790 1756.680 1418.110 1756.740 ;
        RECT 1408.590 1756.540 1418.110 1756.680 ;
        RECT 1408.590 1756.480 1408.910 1756.540 ;
        RECT 1417.790 1756.480 1418.110 1756.540 ;
        RECT 1414.110 1745.460 1414.430 1745.520 ;
        RECT 1472.990 1745.460 1473.310 1745.520 ;
        RECT 1414.110 1745.320 1473.310 1745.460 ;
        RECT 1414.110 1745.260 1414.430 1745.320 ;
        RECT 1472.990 1745.260 1473.310 1745.320 ;
        RECT 1414.110 1738.660 1414.430 1738.720 ;
        RECT 1459.190 1738.660 1459.510 1738.720 ;
        RECT 1414.110 1738.520 1459.510 1738.660 ;
        RECT 1414.110 1738.460 1414.430 1738.520 ;
        RECT 1459.190 1738.460 1459.510 1738.520 ;
        RECT 1409.970 1738.320 1410.290 1738.380 ;
        RECT 1452.290 1738.320 1452.610 1738.380 ;
        RECT 1409.970 1738.180 1452.610 1738.320 ;
        RECT 1409.970 1738.120 1410.290 1738.180 ;
        RECT 1452.290 1738.120 1452.610 1738.180 ;
        RECT 1414.110 1729.140 1414.430 1729.200 ;
        RECT 1438.490 1729.140 1438.810 1729.200 ;
        RECT 1414.110 1729.000 1438.810 1729.140 ;
        RECT 1414.110 1728.940 1414.430 1729.000 ;
        RECT 1438.490 1728.940 1438.810 1729.000 ;
        RECT 1413.650 1723.700 1413.970 1723.760 ;
        RECT 1431.590 1723.700 1431.910 1723.760 ;
        RECT 1413.650 1723.560 1431.910 1723.700 ;
        RECT 1413.650 1723.500 1413.970 1723.560 ;
        RECT 1431.590 1723.500 1431.910 1723.560 ;
        RECT 1409.970 1717.920 1410.290 1717.980 ;
        RECT 1473.450 1717.920 1473.770 1717.980 ;
        RECT 1409.970 1717.780 1473.770 1717.920 ;
        RECT 1409.970 1717.720 1410.290 1717.780 ;
        RECT 1473.450 1717.720 1473.770 1717.780 ;
        RECT 1410.430 1717.580 1410.750 1717.640 ;
        RECT 1424.690 1717.580 1425.010 1717.640 ;
        RECT 1410.430 1717.440 1425.010 1717.580 ;
        RECT 1410.430 1717.380 1410.750 1717.440 ;
        RECT 1424.690 1717.380 1425.010 1717.440 ;
        RECT 1414.110 1711.120 1414.430 1711.180 ;
        RECT 1493.690 1711.120 1494.010 1711.180 ;
        RECT 1414.110 1710.980 1494.010 1711.120 ;
        RECT 1414.110 1710.920 1414.430 1710.980 ;
        RECT 1493.690 1710.920 1494.010 1710.980 ;
        RECT 1409.510 1703.300 1409.830 1703.360 ;
        RECT 1423.310 1703.300 1423.630 1703.360 ;
        RECT 1409.510 1703.160 1423.630 1703.300 ;
        RECT 1409.510 1703.100 1409.830 1703.160 ;
        RECT 1423.310 1703.100 1423.630 1703.160 ;
        RECT 1409.050 1699.560 1409.370 1699.620 ;
        RECT 1422.850 1699.560 1423.170 1699.620 ;
        RECT 1409.050 1699.420 1423.170 1699.560 ;
        RECT 1409.050 1699.360 1409.370 1699.420 ;
        RECT 1422.850 1699.360 1423.170 1699.420 ;
        RECT 1409.510 1694.800 1409.830 1694.860 ;
        RECT 1423.770 1694.800 1424.090 1694.860 ;
        RECT 1409.510 1694.660 1424.090 1694.800 ;
        RECT 1409.510 1694.600 1409.830 1694.660 ;
        RECT 1423.770 1694.600 1424.090 1694.660 ;
        RECT 1409.510 1688.340 1409.830 1688.400 ;
        RECT 1424.230 1688.340 1424.550 1688.400 ;
        RECT 1409.510 1688.200 1424.550 1688.340 ;
        RECT 1409.510 1688.140 1409.830 1688.200 ;
        RECT 1424.230 1688.140 1424.550 1688.200 ;
        RECT 1411.810 1682.900 1412.130 1682.960 ;
        RECT 1427.450 1682.900 1427.770 1682.960 ;
        RECT 1411.810 1682.760 1427.770 1682.900 ;
        RECT 1411.810 1682.700 1412.130 1682.760 ;
        RECT 1427.450 1682.700 1427.770 1682.760 ;
        RECT 1411.810 1678.140 1412.130 1678.200 ;
        RECT 1427.910 1678.140 1428.230 1678.200 ;
        RECT 1411.810 1678.000 1428.230 1678.140 ;
        RECT 1411.810 1677.940 1412.130 1678.000 ;
        RECT 1427.910 1677.940 1428.230 1678.000 ;
        RECT 1410.430 1673.040 1410.750 1673.100 ;
        RECT 1426.990 1673.040 1427.310 1673.100 ;
        RECT 1410.430 1672.900 1427.310 1673.040 ;
        RECT 1410.430 1672.840 1410.750 1672.900 ;
        RECT 1426.990 1672.840 1427.310 1672.900 ;
        RECT 1411.810 1669.640 1412.130 1669.700 ;
        RECT 1459.650 1669.640 1459.970 1669.700 ;
        RECT 1411.810 1669.500 1459.970 1669.640 ;
        RECT 1411.810 1669.440 1412.130 1669.500 ;
        RECT 1459.650 1669.440 1459.970 1669.500 ;
        RECT 1409.510 1668.620 1409.830 1668.680 ;
        RECT 1426.530 1668.620 1426.850 1668.680 ;
        RECT 1409.510 1668.480 1426.850 1668.620 ;
        RECT 1409.510 1668.420 1409.830 1668.480 ;
        RECT 1426.530 1668.420 1426.850 1668.480 ;
        RECT 1414.110 1656.040 1414.430 1656.100 ;
        RECT 1460.110 1656.040 1460.430 1656.100 ;
        RECT 1414.110 1655.900 1460.430 1656.040 ;
        RECT 1414.110 1655.840 1414.430 1655.900 ;
        RECT 1460.110 1655.840 1460.430 1655.900 ;
        RECT 1410.430 1648.220 1410.750 1648.280 ;
        RECT 1425.610 1648.220 1425.930 1648.280 ;
        RECT 1410.430 1648.080 1425.930 1648.220 ;
        RECT 1410.430 1648.020 1410.750 1648.080 ;
        RECT 1425.610 1648.020 1425.930 1648.080 ;
        RECT 1409.510 1647.540 1409.830 1647.600 ;
        RECT 1425.150 1647.540 1425.470 1647.600 ;
        RECT 1409.510 1647.400 1425.470 1647.540 ;
        RECT 1409.510 1647.340 1409.830 1647.400 ;
        RECT 1425.150 1647.340 1425.470 1647.400 ;
        RECT 1410.430 1635.300 1410.750 1635.360 ;
        RECT 1426.070 1635.300 1426.390 1635.360 ;
        RECT 1410.430 1635.160 1426.390 1635.300 ;
        RECT 1410.430 1635.100 1410.750 1635.160 ;
        RECT 1426.070 1635.100 1426.390 1635.160 ;
      LAYER met1 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
        RECT 1550.000 407.860 2647.420 1489.320 ;
      LAYER via ;
        RECT 1890.700 3266.760 1890.960 3267.020 ;
        RECT 1917.840 3266.760 1918.100 3267.020 ;
        RECT 2542.060 3266.760 2542.320 3267.020 ;
        RECT 1890.700 3264.380 1890.960 3264.640 ;
        RECT 1917.840 3264.380 1918.100 3264.640 ;
        RECT 2542.060 3264.040 2542.320 3264.300 ;
        RECT 2566.900 3264.040 2567.160 3264.300 ;
        RECT 646.400 3263.700 646.660 3263.960 ;
        RECT 668.020 3263.700 668.280 3263.960 ;
        RECT 1293.160 3263.700 1293.420 3263.960 ;
        RECT 1317.540 3263.700 1317.800 3263.960 ;
        RECT 2594.500 3263.700 2594.760 3263.960 ;
        RECT 697.000 3263.020 697.260 3263.280 ;
        RECT 1332.260 3252.480 1332.520 3252.740 ;
        RECT 688.260 3251.800 688.520 3252.060 ;
        RECT 1414.140 3252.140 1414.400 3252.400 ;
        RECT 869.040 3251.800 869.300 3252.060 ;
        RECT 2582.080 3252.140 2582.340 3252.400 ;
        RECT 821.200 3251.120 821.460 3251.380 ;
        RECT 927.920 2898.200 928.180 2898.460 ;
        RECT 939.420 2898.200 939.680 2898.460 ;
        RECT 1332.260 3251.120 1332.520 3251.380 ;
        RECT 1407.700 3250.780 1407.960 3251.040 ;
        RECT 1414.140 3250.780 1414.400 3251.040 ;
        RECT 1473.020 3229.360 1473.280 3229.620 ;
        RECT 1536.960 3229.360 1537.220 3229.620 ;
        RECT 1459.220 3222.220 1459.480 3222.480 ;
        RECT 1535.580 3222.220 1535.840 3222.480 ;
        RECT 1452.320 3215.420 1452.580 3215.680 ;
        RECT 1535.580 3215.420 1535.840 3215.680 ;
        RECT 1438.520 3208.620 1438.780 3208.880 ;
        RECT 1538.340 3208.620 1538.600 3208.880 ;
        RECT 1431.620 3201.480 1431.880 3201.740 ;
        RECT 1538.340 3201.480 1538.600 3201.740 ;
        RECT 1424.720 3194.680 1424.980 3194.940 ;
        RECT 1533.280 3194.680 1533.540 3194.940 ;
        RECT 1473.480 3187.880 1473.740 3188.140 ;
        RECT 1534.200 3187.880 1534.460 3188.140 ;
        RECT 1352.040 2901.260 1352.300 2901.520 ;
        RECT 1397.580 2901.260 1397.840 2901.520 ;
        RECT 1459.680 2898.200 1459.940 2898.460 ;
        RECT 1538.340 2898.200 1538.600 2898.460 ;
        RECT 1935.780 3251.120 1936.040 3251.380 ;
        RECT 1732.920 2794.840 1733.180 2795.100 ;
        RECT 386.960 2794.160 387.220 2794.420 ;
        RECT 432.040 2794.160 432.300 2794.420 ;
        RECT 433.420 2794.160 433.680 2794.420 ;
        RECT 482.640 2794.160 482.900 2794.420 ;
        RECT 500.580 2794.160 500.840 2794.420 ;
        RECT 648.240 2794.160 648.500 2794.420 ;
        RECT 1053.040 2794.160 1053.300 2794.420 ;
        RECT 1418.740 2794.160 1419.000 2794.420 ;
        RECT 462.400 2793.820 462.660 2794.080 ;
        RECT 503.800 2793.820 504.060 2794.080 ;
        RECT 375.000 2793.480 375.260 2793.740 ;
        RECT 421.000 2793.480 421.260 2793.740 ;
        RECT 466.540 2793.480 466.800 2793.740 ;
        RECT 513.920 2793.820 514.180 2794.080 ;
        RECT 676.300 2793.820 676.560 2794.080 ;
        RECT 1419.200 2793.820 1419.460 2794.080 ;
        RECT 2415.100 2794.160 2415.360 2794.420 ;
        RECT 526.800 2793.480 527.060 2793.740 ;
        RECT 697.000 2793.480 697.260 2793.740 ;
        RECT 700.220 2793.480 700.480 2793.740 ;
        RECT 1001.060 2793.480 1001.320 2793.740 ;
        RECT 1090.300 2793.480 1090.560 2793.740 ;
        RECT 1094.440 2793.480 1094.700 2793.740 ;
        RECT 1139.980 2793.480 1140.240 2793.740 ;
        RECT 1186.900 2793.480 1187.160 2793.740 ;
        RECT 1642.760 2793.480 1643.020 2793.740 ;
        RECT 1687.840 2793.480 1688.100 2793.740 ;
        RECT 1689.220 2793.480 1689.480 2793.740 ;
        RECT 1723.720 2793.480 1723.980 2793.740 ;
        RECT 1766.500 2793.480 1766.760 2793.740 ;
        RECT 2245.820 2793.480 2246.080 2793.740 ;
        RECT 380.060 2793.140 380.320 2793.400 ;
        RECT 426.980 2793.140 427.240 2793.400 ;
        RECT 475.280 2793.140 475.540 2793.400 ;
        RECT 503.800 2793.140 504.060 2793.400 ;
        RECT 508.860 2793.140 509.120 2793.400 ;
        RECT 662.500 2793.140 662.760 2793.400 ;
        RECT 686.420 2793.140 686.680 2793.400 ;
        RECT 986.800 2793.140 987.060 2793.400 ;
        RECT 1083.400 2793.140 1083.660 2793.400 ;
        RECT 1129.400 2793.140 1129.660 2793.400 ;
        RECT 1173.100 2793.140 1173.360 2793.400 ;
        RECT 1780.300 2793.140 1780.560 2793.400 ;
        RECT 2284.460 2793.820 2284.720 2794.080 ;
        RECT 2301.020 2793.820 2301.280 2794.080 ;
        RECT 2304.240 2793.820 2304.500 2794.080 ;
        RECT 2347.480 2793.820 2347.740 2794.080 ;
        RECT 2385.660 2793.820 2385.920 2794.080 ;
        RECT 2428.900 2793.820 2429.160 2794.080 ;
        RECT 2308.840 2793.480 2309.100 2793.740 ;
        RECT 2356.680 2793.480 2356.940 2793.740 ;
        RECT 2402.680 2793.480 2402.940 2793.740 ;
        RECT 2298.260 2793.140 2298.520 2793.400 ;
        RECT 2343.800 2793.140 2344.060 2793.400 ;
        RECT 2391.640 2793.140 2391.900 2793.400 ;
        RECT 2435.800 2793.140 2436.060 2793.400 ;
        RECT 409.960 2792.800 410.220 2793.060 ;
        RECT 455.500 2792.800 455.760 2793.060 ;
        RECT 537.380 2792.800 537.640 2793.060 ;
        RECT 865.820 2792.800 866.080 2793.060 ;
        RECT 1122.040 2792.800 1122.300 2793.060 ;
        RECT 1166.200 2792.800 1166.460 2793.060 ;
        RECT 1677.260 2792.800 1677.520 2793.060 ;
        RECT 1723.720 2792.800 1723.980 2793.060 ;
        RECT 1741.200 2792.800 1741.460 2793.060 ;
        RECT 1787.200 2792.800 1787.460 2793.060 ;
        RECT 2273.420 2792.800 2273.680 2793.060 ;
        RECT 2321.720 2792.800 2321.980 2793.060 ;
        RECT 2367.260 2792.800 2367.520 2793.060 ;
        RECT 2415.100 2792.800 2415.360 2793.060 ;
        RECT 397.080 2792.460 397.340 2792.720 ;
        RECT 444.460 2792.460 444.720 2792.720 ;
        RECT 492.760 2792.460 493.020 2792.720 ;
        RECT 539.220 2792.460 539.480 2792.720 ;
        RECT 544.280 2792.460 544.540 2792.720 ;
        RECT 872.720 2792.460 872.980 2792.720 ;
        RECT 1042.460 2792.460 1042.720 2792.720 ;
        RECT 1087.540 2792.460 1087.800 2792.720 ;
        RECT 1135.840 2792.460 1136.100 2792.720 ;
        RECT 1180.000 2792.460 1180.260 2792.720 ;
        RECT 392.480 2792.120 392.740 2792.380 ;
        RECT 439.400 2792.120 439.660 2792.380 ;
        RECT 524.040 2792.120 524.300 2792.380 ;
        RECT 858.920 2792.120 859.180 2792.380 ;
        RECT 1055.800 2792.120 1056.060 2792.380 ;
        RECT 1059.020 2792.120 1059.280 2792.380 ;
        RECT 1105.480 2792.120 1105.740 2792.380 ;
        RECT 1152.400 2792.120 1152.660 2792.380 ;
        RECT 1420.580 2792.120 1420.840 2792.380 ;
        RECT 1652.880 2792.460 1653.140 2792.720 ;
        RECT 368.560 2791.780 368.820 2792.040 ;
        RECT 362.120 2791.100 362.380 2791.360 ;
        RECT 433.420 2791.780 433.680 2792.040 ;
        RECT 478.500 2791.780 478.760 2792.040 ;
        RECT 510.240 2791.780 510.500 2792.040 ;
        RECT 852.020 2791.780 852.280 2792.040 ;
        RECT 1100.880 2791.780 1101.140 2792.040 ;
        RECT 1146.420 2791.780 1146.680 2792.040 ;
        RECT 1549.380 2791.780 1549.640 2792.040 ;
        RECT 1596.300 2791.780 1596.560 2792.040 ;
        RECT 1690.600 2792.460 1690.860 2792.720 ;
        RECT 1695.200 2792.460 1695.460 2792.720 ;
        RECT 2268.360 2792.460 2268.620 2792.720 ;
        RECT 2315.280 2792.460 2315.540 2792.720 ;
        RECT 2361.280 2792.460 2361.540 2792.720 ;
        RECT 2408.200 2792.460 2408.460 2792.720 ;
        RECT 1662.540 2792.120 1662.800 2792.380 ;
        RECT 1706.240 2792.120 1706.500 2792.380 ;
        RECT 1752.700 2792.120 1752.960 2792.380 ;
        RECT 2266.520 2792.120 2266.780 2792.380 ;
        RECT 2284.460 2792.120 2284.720 2792.380 ;
        RECT 2333.680 2792.120 2333.940 2792.380 ;
        RECT 2340.120 2792.120 2340.380 2792.380 ;
        RECT 2347.480 2792.120 2347.740 2792.380 ;
        RECT 2394.860 2792.120 2395.120 2792.380 ;
        RECT 1699.340 2791.780 1699.600 2792.040 ;
        RECT 403.980 2791.440 404.240 2791.700 ;
        RECT 450.440 2791.440 450.700 2791.700 ;
        RECT 501.040 2791.440 501.300 2791.700 ;
        RECT 501.960 2791.440 502.220 2791.700 ;
        RECT 845.120 2791.440 845.380 2791.700 ;
        RECT 414.560 2791.100 414.820 2791.360 ;
        RECT 462.400 2791.100 462.660 2791.360 ;
        RECT 489.080 2791.100 489.340 2791.360 ;
        RECT 838.220 2791.100 838.480 2791.360 ;
        RECT 371.320 2790.760 371.580 2791.020 ;
        RECT 745.300 2790.760 745.560 2791.020 ;
        RECT 1019.000 2790.760 1019.260 2791.020 ;
        RECT 1065.460 2791.440 1065.720 2791.700 ;
        RECT 1111.460 2791.440 1111.720 2791.700 ;
        RECT 1159.300 2791.440 1159.560 2791.700 ;
        RECT 1682.320 2791.440 1682.580 2791.700 ;
        RECT 1728.780 2791.440 1729.040 2791.700 ;
        RECT 2326.780 2791.780 2327.040 2792.040 ;
        RECT 2374.160 2791.780 2374.420 2792.040 ;
        RECT 2415.100 2791.780 2415.360 2792.040 ;
        RECT 1747.640 2791.440 1747.900 2791.700 ;
        RECT 1794.100 2791.440 1794.360 2791.700 ;
        RECT 2090.800 2791.440 2091.060 2791.700 ;
        RECT 2279.860 2791.440 2280.120 2791.700 ;
        RECT 2301.480 2791.440 2301.740 2791.700 ;
        RECT 2435.800 2791.440 2436.060 2791.700 ;
        RECT 1034.640 2791.100 1034.900 2791.360 ;
        RECT 1076.500 2791.100 1076.760 2791.360 ;
        RECT 1122.040 2791.100 1122.300 2791.360 ;
        RECT 1146.420 2791.100 1146.680 2791.360 ;
        RECT 1193.800 2791.100 1194.060 2791.360 ;
        RECT 1411.380 2791.100 1411.640 2791.360 ;
        RECT 1587.100 2791.100 1587.360 2791.360 ;
        RECT 1069.600 2790.760 1069.860 2791.020 ;
        RECT 1118.360 2790.760 1118.620 2791.020 ;
        RECT 1159.300 2790.760 1159.560 2791.020 ;
        RECT 1425.180 2790.760 1425.440 2791.020 ;
        RECT 1600.900 2790.760 1601.160 2791.020 ;
        RECT 384.660 2790.420 384.920 2790.680 ;
        RECT 766.000 2790.420 766.260 2790.680 ;
        RECT 1411.840 2790.420 1412.100 2790.680 ;
        RECT 1613.320 2790.420 1613.580 2790.680 ;
        RECT 1659.320 2790.760 1659.580 2791.020 ;
        RECT 1662.540 2790.760 1662.800 2791.020 ;
        RECT 1624.820 2790.420 1625.080 2790.680 ;
        RECT 1670.360 2791.100 1670.620 2791.360 ;
        RECT 1718.200 2791.100 1718.460 2791.360 ;
        RECT 1724.640 2791.100 1724.900 2791.360 ;
        RECT 1773.400 2791.100 1773.660 2791.360 ;
        RECT 2266.980 2791.100 2267.240 2791.360 ;
        RECT 2428.900 2791.100 2429.160 2791.360 ;
        RECT 1669.440 2790.760 1669.700 2791.020 ;
        RECT 1712.680 2790.760 1712.940 2791.020 ;
        RECT 1759.600 2790.760 1759.860 2791.020 ;
        RECT 1797.320 2790.760 1797.580 2791.020 ;
        RECT 2387.500 2790.760 2387.760 2791.020 ;
        RECT 2394.860 2790.760 2395.120 2791.020 ;
        RECT 2442.700 2790.760 2442.960 2791.020 ;
        RECT 1724.640 2790.420 1724.900 2790.680 ;
        RECT 1760.060 2790.420 1760.320 2790.680 ;
        RECT 1783.520 2790.420 1783.780 2790.680 ;
        RECT 2373.700 2790.420 2373.960 2790.680 ;
        RECT 2377.380 2790.420 2377.640 2790.680 ;
        RECT 2422.000 2790.420 2422.260 2790.680 ;
        RECT 396.620 2790.080 396.880 2790.340 ;
        RECT 786.700 2790.080 786.960 2790.340 ;
        RECT 1420.120 2790.080 1420.380 2790.340 ;
        RECT 1636.780 2790.080 1637.040 2790.340 ;
        RECT 1741.200 2790.080 1741.460 2790.340 ;
        RECT 1790.420 2790.080 1790.680 2790.340 ;
        RECT 2380.600 2790.080 2380.860 2790.340 ;
        RECT 406.280 2789.740 406.540 2790.000 ;
        RECT 807.400 2789.740 807.660 2790.000 ;
        RECT 1419.660 2789.740 1419.920 2790.000 ;
        RECT 1642.760 2789.740 1643.020 2790.000 ;
        RECT 1797.780 2789.740 1798.040 2790.000 ;
        RECT 2394.400 2789.740 2394.660 2790.000 ;
        RECT 484.940 2789.400 485.200 2789.660 ;
        RECT 534.620 2789.400 534.880 2789.660 ;
        RECT 539.220 2789.400 539.480 2789.660 ;
        RECT 717.700 2789.400 717.960 2789.660 ;
        RECT 1549.840 2789.400 1550.100 2789.660 ;
        RECT 1642.300 2789.400 1642.560 2789.660 ;
        RECT 1645.520 2789.400 1645.780 2789.660 ;
        RECT 1648.280 2789.400 1648.540 2789.660 ;
        RECT 1690.600 2789.400 1690.860 2789.660 ;
        RECT 1762.820 2789.400 1763.080 2789.660 ;
        RECT 2380.600 2789.400 2380.860 2789.660 ;
        RECT 418.700 2789.060 418.960 2789.320 ;
        RECT 828.100 2789.060 828.360 2789.320 ;
        RECT 1010.720 2789.060 1010.980 2789.320 ;
        RECT 1055.800 2789.060 1056.060 2789.320 ;
        RECT 1410.920 2789.060 1411.180 2789.320 ;
        RECT 413.640 2788.720 413.900 2788.980 ;
        RECT 465.620 2788.720 465.880 2788.980 ;
        RECT 475.280 2788.720 475.540 2788.980 ;
        RECT 520.820 2788.720 521.080 2788.980 ;
        RECT 627.540 2788.720 627.800 2788.980 ;
        RECT 1042.460 2788.720 1042.720 2788.980 ;
        RECT 1417.820 2788.720 1418.080 2788.980 ;
        RECT 399.840 2788.380 400.100 2788.640 ;
        RECT 444.920 2788.380 445.180 2788.640 ;
        RECT 606.840 2788.380 607.100 2788.640 ;
        RECT 1034.640 2788.380 1034.900 2788.640 ;
        RECT 1045.220 2788.380 1045.480 2788.640 ;
        RECT 1090.300 2788.380 1090.560 2788.640 ;
        RECT 1418.280 2788.380 1418.540 2788.640 ;
        RECT 2218.220 2789.060 2218.480 2789.320 ;
        RECT 2402.680 2789.060 2402.940 2789.320 ;
        RECT 2235.700 2788.720 2235.960 2788.980 ;
        RECT 2238.920 2788.720 2239.180 2788.980 ;
        RECT 378.680 2788.040 378.940 2788.300 ;
        RECT 424.220 2788.040 424.480 2788.300 ;
        RECT 455.500 2788.040 455.760 2788.300 ;
        RECT 500.120 2788.040 500.380 2788.300 ;
        RECT 501.040 2788.040 501.300 2788.300 ;
        RECT 541.520 2788.040 541.780 2788.300 ;
        RECT 586.140 2788.040 586.400 2788.300 ;
        RECT 1019.000 2788.040 1019.260 2788.300 ;
        RECT 1024.520 2788.040 1024.780 2788.300 ;
        RECT 1069.600 2788.040 1069.860 2788.300 ;
        RECT 1617.920 2788.040 1618.180 2788.300 ;
        RECT 1669.440 2788.040 1669.700 2788.300 ;
        RECT 390.640 2787.700 390.900 2787.960 ;
        RECT 431.120 2787.700 431.380 2787.960 ;
        RECT 479.420 2787.700 479.680 2787.960 ;
        RECT 1007.500 2787.700 1007.760 2787.960 ;
        RECT 1038.320 2787.700 1038.580 2787.960 ;
        RECT 1083.400 2787.700 1083.660 2787.960 ;
        RECT 1548.920 2787.700 1549.180 2787.960 ;
        RECT 1628.500 2787.700 1628.760 2787.960 ;
        RECT 1631.720 2787.700 1631.980 2787.960 ;
        RECT 1677.260 2787.700 1677.520 2787.960 ;
        RECT 1828.140 2788.040 1828.400 2788.300 ;
        RECT 1869.540 2788.040 1869.800 2788.300 ;
        RECT 2408.200 2788.720 2408.460 2788.980 ;
        RECT 2415.100 2788.380 2415.360 2788.640 ;
        RECT 2090.800 2788.040 2091.060 2788.300 ;
        RECT 2232.020 2788.040 2232.280 2788.300 ;
        RECT 2294.120 2788.040 2294.380 2788.300 ;
        RECT 2333.680 2788.040 2333.940 2788.300 ;
        RECT 2377.380 2788.040 2377.640 2788.300 ;
        RECT 2252.720 2787.700 2252.980 2787.960 ;
        RECT 2422.000 2787.700 2422.260 2787.960 ;
        RECT 365.340 2731.600 365.600 2731.860 ;
        RECT 740.700 2731.600 740.960 2731.860 ;
        RECT 427.440 2731.260 427.700 2731.520 ;
        RECT 844.200 2731.260 844.460 2731.520 ;
        RECT 433.880 2730.920 434.140 2731.180 ;
        RECT 854.780 2730.920 855.040 2731.180 ;
        RECT 434.340 2730.580 434.600 2730.840 ;
        RECT 865.360 2730.580 865.620 2730.840 ;
        RECT 441.240 2730.240 441.500 2730.500 ;
        RECT 875.480 2730.240 875.740 2730.500 ;
        RECT 455.040 2729.900 455.300 2730.160 ;
        RECT 896.180 2729.900 896.440 2730.160 ;
        RECT 448.140 2729.560 448.400 2729.820 ;
        RECT 886.060 2729.560 886.320 2729.820 ;
        RECT 461.940 2729.220 462.200 2729.480 ;
        RECT 906.760 2729.220 907.020 2729.480 ;
        RECT 468.840 2728.880 469.100 2729.140 ;
        RECT 916.880 2728.880 917.140 2729.140 ;
        RECT 468.380 2728.540 468.640 2728.800 ;
        RECT 927.460 2728.540 927.720 2728.800 ;
        RECT 288.980 2725.140 289.240 2725.400 ;
        RECT 553.940 2725.140 554.200 2725.400 ;
        RECT 289.440 2724.800 289.700 2725.060 ;
        RECT 564.060 2724.800 564.320 2725.060 ;
        RECT 475.740 2724.460 476.000 2724.720 ;
        RECT 937.580 2724.460 937.840 2724.720 ;
        RECT 481.260 2724.120 481.520 2724.380 ;
        RECT 941.720 2724.120 941.980 2724.380 ;
        RECT 470.680 2723.780 470.940 2724.040 ;
        RECT 942.180 2723.780 942.440 2724.040 ;
        RECT 460.560 2723.440 460.820 2723.700 ;
        RECT 942.640 2723.440 942.900 2723.700 ;
        RECT 449.980 2723.100 450.240 2723.360 ;
        RECT 943.100 2723.100 943.360 2723.360 ;
        RECT 439.860 2722.760 440.120 2723.020 ;
        RECT 943.560 2722.760 943.820 2723.020 ;
        RECT 429.280 2722.420 429.540 2722.680 ;
        RECT 944.020 2722.420 944.280 2722.680 ;
        RECT 419.160 2722.080 419.420 2722.340 ;
        RECT 944.480 2722.080 944.740 2722.340 ;
        RECT 408.580 2721.740 408.840 2722.000 ;
        RECT 979.900 2721.740 980.160 2722.000 ;
        RECT 288.520 2721.400 288.780 2721.660 ;
        RECT 543.360 2721.400 543.620 2721.660 ;
        RECT 288.060 2721.060 288.320 2721.320 ;
        RECT 533.240 2721.060 533.500 2721.320 ;
        RECT 287.600 2720.720 287.860 2720.980 ;
        RECT 522.660 2720.720 522.920 2720.980 ;
        RECT 287.140 2720.380 287.400 2720.640 ;
        RECT 512.540 2720.380 512.800 2720.640 ;
        RECT 358.440 2718.340 358.700 2718.600 ;
        RECT 377.300 2718.340 377.560 2718.600 ;
        RECT 636.740 2718.340 637.000 2718.600 ;
        RECT 1045.220 2718.340 1045.480 2718.600 ;
        RECT 1145.040 2718.340 1145.300 2718.600 ;
        RECT 1300.980 2718.340 1301.240 2718.600 ;
        RECT 616.040 2718.000 616.300 2718.260 ;
        RECT 1038.320 2718.000 1038.580 2718.260 ;
        RECT 1138.140 2718.000 1138.400 2718.260 ;
        RECT 1290.400 2718.000 1290.660 2718.260 ;
        RECT 351.080 2717.660 351.340 2717.920 ;
        RECT 356.600 2717.660 356.860 2717.920 ;
        RECT 595.340 2717.660 595.600 2717.920 ;
        RECT 1024.520 2717.660 1024.780 2717.920 ;
        RECT 1041.540 2717.660 1041.800 2717.920 ;
        RECT 1114.220 2717.660 1114.480 2717.920 ;
        RECT 1158.840 2717.660 1159.100 2717.920 ;
        RECT 1321.680 2717.660 1321.940 2717.920 ;
        RECT 574.640 2717.320 574.900 2717.580 ;
        RECT 1010.720 2717.320 1010.980 2717.580 ;
        RECT 1048.440 2717.320 1048.700 2717.580 ;
        RECT 1124.340 2717.320 1124.600 2717.580 ;
        RECT 1151.940 2717.320 1152.200 2717.580 ;
        RECT 1311.100 2717.320 1311.360 2717.580 ;
        RECT 500.580 2716.980 500.840 2717.240 ;
        RECT 948.160 2716.980 948.420 2717.240 ;
        RECT 1055.340 2716.980 1055.600 2717.240 ;
        RECT 1134.920 2716.980 1135.180 2717.240 ;
        RECT 1165.740 2716.980 1166.000 2717.240 ;
        RECT 1332.260 2716.980 1332.520 2717.240 ;
        RECT 315.200 2716.640 315.460 2716.900 ;
        RECT 410.420 2716.640 410.680 2716.900 ;
        RECT 496.440 2716.640 496.700 2716.900 ;
        RECT 968.860 2716.640 969.120 2716.900 ;
        RECT 1062.240 2716.640 1062.500 2716.900 ;
        RECT 1155.620 2716.640 1155.880 2716.900 ;
        RECT 1165.280 2716.640 1165.540 2716.900 ;
        RECT 1342.380 2716.640 1342.640 2716.900 ;
        RECT 286.220 2716.300 286.480 2716.560 ;
        RECT 398.460 2716.300 398.720 2716.560 ;
        RECT 509.780 2716.300 510.040 2716.560 ;
        RECT 989.560 2716.300 989.820 2716.560 ;
        RECT 1076.040 2716.300 1076.300 2716.560 ;
        RECT 1176.320 2716.300 1176.580 2716.560 ;
        RECT 1179.540 2716.300 1179.800 2716.560 ;
        RECT 1363.080 2716.300 1363.340 2716.560 ;
        RECT 335.900 2715.960 336.160 2716.220 ;
        RECT 479.420 2715.960 479.680 2716.220 ;
        RECT 517.140 2715.960 517.400 2716.220 ;
        RECT 1010.260 2715.960 1010.520 2716.220 ;
        RECT 1054.880 2715.960 1055.140 2716.220 ;
        RECT 1145.500 2715.960 1145.760 2716.220 ;
        RECT 1172.640 2715.960 1172.900 2716.220 ;
        RECT 1352.960 2715.960 1353.220 2716.220 ;
        RECT 337.740 2715.620 338.000 2715.880 ;
        RECT 491.840 2715.620 492.100 2715.880 ;
        RECT 530.940 2715.620 531.200 2715.880 ;
        RECT 1030.960 2715.620 1031.220 2715.880 ;
        RECT 1069.140 2715.620 1069.400 2715.880 ;
        RECT 1166.200 2715.620 1166.460 2715.880 ;
        RECT 1186.440 2715.620 1186.700 2715.880 ;
        RECT 1373.660 2715.620 1373.920 2715.880 ;
        RECT 286.680 2715.280 286.940 2715.540 ;
        RECT 501.960 2715.280 502.220 2715.540 ;
        RECT 551.640 2715.280 551.900 2715.540 ;
        RECT 1062.240 2715.280 1062.500 2715.540 ;
        RECT 1082.940 2715.280 1083.200 2715.540 ;
        RECT 1186.900 2715.280 1187.160 2715.540 ;
        RECT 1193.340 2715.280 1193.600 2715.540 ;
        RECT 1383.780 2715.280 1384.040 2715.540 ;
        RECT 387.880 2714.940 388.140 2715.200 ;
        RECT 927.920 2714.940 928.180 2715.200 ;
        RECT 1013.940 2714.940 1014.200 2715.200 ;
        RECT 1072.820 2714.940 1073.080 2715.200 ;
        RECT 1089.380 2714.940 1089.640 2715.200 ;
        RECT 1197.020 2714.940 1197.280 2715.200 ;
        RECT 1200.240 2714.940 1200.500 2715.200 ;
        RECT 1394.360 2714.940 1394.620 2715.200 ;
        RECT 325.780 2714.600 326.040 2714.860 ;
        RECT 700.220 2714.600 700.480 2714.860 ;
        RECT 872.720 2714.600 872.980 2714.860 ;
        RECT 1052.120 2714.600 1052.380 2714.860 ;
        RECT 1103.640 2714.600 1103.900 2714.860 ;
        RECT 444.920 2714.260 445.180 2714.520 ;
        RECT 802.800 2714.260 803.060 2714.520 ;
        RECT 865.820 2714.260 866.080 2714.520 ;
        RECT 1041.540 2714.260 1041.800 2714.520 ;
        RECT 351.540 2713.920 351.800 2714.180 ;
        RECT 367.180 2713.920 367.440 2714.180 ;
        RECT 465.620 2713.920 465.880 2714.180 ;
        RECT 823.500 2713.920 823.760 2714.180 ;
        RECT 858.920 2713.920 859.180 2714.180 ;
        RECT 1020.840 2713.920 1021.100 2714.180 ;
        RECT 1034.640 2713.920 1034.900 2714.180 ;
        RECT 1103.640 2713.920 1103.900 2714.180 ;
        RECT 431.120 2713.580 431.380 2713.840 ;
        RECT 782.100 2713.580 782.360 2713.840 ;
        RECT 852.020 2713.580 852.280 2713.840 ;
        RECT 1000.140 2713.580 1000.400 2713.840 ;
        RECT 1027.740 2713.580 1028.000 2713.840 ;
        RECT 1093.520 2713.580 1093.780 2713.840 ;
        RECT 424.220 2713.240 424.480 2713.500 ;
        RECT 761.400 2713.240 761.660 2713.500 ;
        RECT 845.120 2713.240 845.380 2713.500 ;
        RECT 979.440 2713.240 979.700 2713.500 ;
        RECT 1021.300 2713.240 1021.560 2713.500 ;
        RECT 1082.940 2713.240 1083.200 2713.500 ;
        RECT 1131.240 2714.600 1131.500 2714.860 ;
        RECT 1280.280 2714.600 1280.540 2714.860 ;
        RECT 1130.780 2714.260 1131.040 2714.520 ;
        RECT 1269.700 2714.260 1269.960 2714.520 ;
        RECT 1117.440 2713.920 1117.700 2714.180 ;
        RECT 1249.000 2713.920 1249.260 2714.180 ;
        RECT 1123.420 2713.580 1123.680 2713.840 ;
        RECT 1259.580 2713.580 1259.840 2713.840 ;
        RECT 1228.300 2713.240 1228.560 2713.500 ;
        RECT 541.520 2712.900 541.780 2713.160 ;
        RECT 730.120 2712.900 730.380 2713.160 ;
        RECT 838.220 2712.900 838.480 2713.160 ;
        RECT 958.740 2712.900 959.000 2713.160 ;
        RECT 1110.540 2712.900 1110.800 2713.160 ;
        RECT 1238.880 2712.900 1239.140 2713.160 ;
        RECT 534.620 2712.560 534.880 2712.820 ;
        RECT 709.420 2712.560 709.680 2712.820 ;
        RECT 1089.840 2712.560 1090.100 2712.820 ;
        RECT 1207.600 2712.560 1207.860 2712.820 ;
        RECT 520.820 2712.220 521.080 2712.480 ;
        RECT 688.720 2712.220 688.980 2712.480 ;
        RECT 1096.740 2712.220 1097.000 2712.480 ;
        RECT 1217.720 2712.220 1217.980 2712.480 ;
        RECT 500.120 2711.880 500.380 2712.140 ;
        RECT 657.440 2711.880 657.700 2712.140 ;
        RECT 1410.460 2152.580 1410.720 2152.840 ;
        RECT 2307.920 2152.580 2308.180 2152.840 ;
        RECT 1414.140 2145.440 1414.400 2145.700 ;
        RECT 2301.480 2145.440 2301.740 2145.700 ;
        RECT 1414.140 2138.640 1414.400 2138.900 ;
        RECT 2266.980 2138.640 2267.240 2138.900 ;
        RECT 1413.680 2138.300 1413.940 2138.560 ;
        RECT 2252.720 2138.300 2252.980 2138.560 ;
        RECT 1410.460 2131.840 1410.720 2132.100 ;
        RECT 2245.820 2131.840 2246.080 2132.100 ;
        RECT 1414.140 2125.040 1414.400 2125.300 ;
        RECT 2238.920 2125.040 2239.180 2125.300 ;
        RECT 1414.140 2117.900 1414.400 2118.160 ;
        RECT 2232.020 2117.900 2232.280 2118.160 ;
        RECT 1410.460 2117.560 1410.720 2117.820 ;
        RECT 2218.220 2117.560 2218.480 2117.820 ;
        RECT 1414.140 2111.100 1414.400 2111.360 ;
        RECT 1797.780 2111.100 1798.040 2111.360 ;
        RECT 1414.140 2104.300 1414.400 2104.560 ;
        RECT 1797.320 2104.300 1797.580 2104.560 ;
        RECT 1414.140 2097.160 1414.400 2097.420 ;
        RECT 1790.420 2097.160 1790.680 2097.420 ;
        RECT 1410.460 2096.820 1410.720 2097.080 ;
        RECT 1762.820 2096.820 1763.080 2097.080 ;
        RECT 1409.540 2090.360 1409.800 2090.620 ;
        RECT 1783.520 2090.360 1783.780 2090.620 ;
        RECT 1425.640 2087.640 1425.900 2087.900 ;
        RECT 1594.000 2087.640 1594.260 2087.900 ;
        RECT 1422.420 2087.300 1422.680 2087.560 ;
        RECT 1617.920 2087.300 1618.180 2087.560 ;
        RECT 1416.900 2086.960 1417.160 2087.220 ;
        RECT 1645.520 2086.960 1645.780 2087.220 ;
        RECT 1414.140 2083.560 1414.400 2083.820 ;
        RECT 2366.800 2083.560 2367.060 2083.820 ;
        RECT 1436.680 2083.220 1436.940 2083.480 ;
        RECT 2263.300 2083.220 2263.560 2083.480 ;
        RECT 1436.220 2082.880 1436.480 2083.140 ;
        RECT 2263.760 2082.880 2264.020 2083.140 ;
        RECT 1412.760 2082.540 1413.020 2082.800 ;
        RECT 2266.520 2082.540 2266.780 2082.800 ;
        RECT 1412.300 2082.200 1412.560 2082.460 ;
        RECT 2270.200 2082.200 2270.460 2082.460 ;
        RECT 1435.760 2081.860 1436.020 2082.120 ;
        RECT 2305.160 2081.860 2305.420 2082.120 ;
        RECT 1421.960 2081.520 1422.220 2081.780 ;
        RECT 2297.800 2081.520 2298.060 2081.780 ;
        RECT 1414.600 2081.180 1414.860 2081.440 ;
        RECT 2318.500 2081.180 2318.760 2081.440 ;
        RECT 1409.540 2080.840 1409.800 2081.100 ;
        RECT 2325.400 2080.840 2325.660 2081.100 ;
        RECT 1408.620 2080.500 1408.880 2080.760 ;
        RECT 2332.300 2080.500 2332.560 2080.760 ;
        RECT 1409.080 2080.160 1409.340 2080.420 ;
        RECT 2339.660 2080.160 2339.920 2080.420 ;
        RECT 1440.360 2079.820 1440.620 2080.080 ;
        RECT 1663.000 2079.820 1663.260 2080.080 ;
        RECT 1439.440 2079.480 1439.700 2079.740 ;
        RECT 1656.100 2079.480 1656.360 2079.740 ;
        RECT 1417.360 2079.140 1417.620 2079.400 ;
        RECT 1624.820 2079.140 1625.080 2079.400 ;
        RECT 1494.180 2078.800 1494.440 2079.060 ;
        RECT 1631.720 2078.800 1631.980 2079.060 ;
        RECT 1414.140 2076.760 1414.400 2077.020 ;
        RECT 2359.900 2076.760 2360.160 2077.020 ;
        RECT 1413.680 2076.420 1413.940 2076.680 ;
        RECT 2353.000 2076.420 2353.260 2076.680 ;
        RECT 1429.780 2076.080 1430.040 2076.340 ;
        RECT 1745.800 2076.080 1746.060 2076.340 ;
        RECT 1440.820 2075.740 1441.080 2076.000 ;
        RECT 1760.520 2075.740 1760.780 2076.000 ;
        RECT 1428.860 2075.400 1429.120 2075.660 ;
        RECT 1752.700 2075.400 1752.960 2075.660 ;
        RECT 1441.280 2075.060 1441.540 2075.320 ;
        RECT 1766.500 2075.060 1766.760 2075.320 ;
        RECT 1441.740 2074.720 1442.000 2074.980 ;
        RECT 1773.860 2074.720 1774.120 2074.980 ;
        RECT 1428.400 2074.380 1428.660 2074.640 ;
        RECT 1760.060 2074.380 1760.320 2074.640 ;
        RECT 1438.060 2074.040 1438.320 2074.300 ;
        RECT 1780.300 2074.040 1780.560 2074.300 ;
        RECT 1437.600 2073.700 1437.860 2073.960 ;
        RECT 1787.200 2073.700 1787.460 2073.960 ;
        RECT 1437.140 2073.360 1437.400 2073.620 ;
        RECT 1794.560 2073.360 1794.820 2073.620 ;
        RECT 1430.240 2073.020 1430.500 2073.280 ;
        RECT 1738.900 2073.020 1739.160 2073.280 ;
        RECT 1439.900 2072.680 1440.160 2072.940 ;
        RECT 1649.200 2072.680 1649.460 2072.940 ;
        RECT 1432.540 2072.340 1432.800 2072.600 ;
        RECT 1621.600 2072.340 1621.860 2072.600 ;
        RECT 1494.640 2072.000 1494.900 2072.260 ;
        RECT 1649.660 2072.000 1649.920 2072.260 ;
        RECT 1414.140 2069.620 1414.400 2069.880 ;
        RECT 2346.100 2069.620 2346.360 2069.880 ;
        RECT 1433.460 2069.280 1433.720 2069.540 ;
        RECT 1684.160 2069.280 1684.420 2069.540 ;
        RECT 1434.380 2068.940 1434.640 2069.200 ;
        RECT 1697.500 2068.940 1697.760 2069.200 ;
        RECT 1416.440 2068.600 1416.700 2068.860 ;
        RECT 1683.700 2068.600 1683.960 2068.860 ;
        RECT 1415.980 2068.260 1416.240 2068.520 ;
        RECT 1690.600 2068.260 1690.860 2068.520 ;
        RECT 1434.840 2067.920 1435.100 2068.180 ;
        RECT 1711.300 2067.920 1711.560 2068.180 ;
        RECT 1430.700 2067.580 1430.960 2067.840 ;
        RECT 1718.200 2067.580 1718.460 2067.840 ;
        RECT 1415.520 2067.240 1415.780 2067.500 ;
        RECT 1704.400 2067.240 1704.660 2067.500 ;
        RECT 1431.160 2066.900 1431.420 2067.160 ;
        RECT 1725.100 2066.900 1725.360 2067.160 ;
        RECT 1429.320 2066.560 1429.580 2066.820 ;
        RECT 1732.000 2066.560 1732.260 2066.820 ;
        RECT 1415.060 2066.220 1415.320 2066.480 ;
        RECT 1718.660 2066.220 1718.920 2066.480 ;
        RECT 1433.920 2065.880 1434.180 2066.140 ;
        RECT 1676.800 2065.880 1677.060 2066.140 ;
        RECT 1433.000 2065.540 1433.260 2065.800 ;
        RECT 1669.900 2065.540 1670.160 2065.800 ;
        RECT 1432.080 2065.200 1432.340 2065.460 ;
        RECT 1607.800 2065.200 1608.060 2065.460 ;
        RECT 1466.120 2064.860 1466.380 2065.120 ;
        RECT 1614.700 2064.860 1614.960 2065.120 ;
        RECT 1412.300 2063.160 1412.560 2063.420 ;
        RECT 1413.680 2063.160 1413.940 2063.420 ;
        RECT 1414.140 2062.820 1414.400 2063.080 ;
        RECT 2339.200 2062.820 2339.460 2063.080 ;
        RECT 1427.020 2062.480 1427.280 2062.740 ;
        RECT 2193.380 2062.480 2193.640 2062.740 ;
        RECT 1423.340 2062.140 1423.600 2062.400 ;
        RECT 2190.620 2062.140 2190.880 2062.400 ;
        RECT 1423.800 2061.800 1424.060 2062.060 ;
        RECT 2191.540 2061.800 2191.800 2062.060 ;
        RECT 1424.260 2061.460 1424.520 2061.720 ;
        RECT 2192.000 2061.460 2192.260 2061.720 ;
        RECT 1422.880 2061.120 1423.140 2061.380 ;
        RECT 2191.080 2061.120 2191.340 2061.380 ;
        RECT 1426.560 2060.780 1426.820 2061.040 ;
        RECT 2228.800 2060.780 2229.060 2061.040 ;
        RECT 1426.100 2060.440 1426.360 2060.700 ;
        RECT 2256.400 2060.440 2256.660 2060.700 ;
        RECT 1410.000 2060.100 1410.260 2060.360 ;
        RECT 2242.600 2060.100 2242.860 2060.360 ;
        RECT 1438.980 2059.760 1439.240 2060.020 ;
        RECT 2301.020 2059.760 2301.280 2060.020 ;
        RECT 1421.040 2059.420 1421.300 2059.680 ;
        RECT 2294.120 2059.420 2294.380 2059.680 ;
        RECT 1427.480 2059.080 1427.740 2059.340 ;
        RECT 2192.460 2059.080 2192.720 2059.340 ;
        RECT 1427.940 2058.740 1428.200 2059.000 ;
        RECT 2192.920 2058.740 2193.180 2059.000 ;
        RECT 1460.140 2058.400 1460.400 2058.660 ;
        RECT 1601.360 2058.400 1601.620 2058.660 ;
        RECT 1493.720 2058.060 1493.980 2058.320 ;
        RECT 1580.200 2058.060 1580.460 2058.320 ;
        RECT 1410.000 2056.360 1410.260 2056.620 ;
        RECT 1410.000 2054.320 1410.260 2054.580 ;
        RECT 2273.420 2054.320 2273.680 2054.580 ;
        RECT 1412.300 2053.980 1412.560 2054.240 ;
        RECT 2277.100 2053.980 2277.360 2054.240 ;
        RECT 1414.140 2053.640 1414.400 2053.900 ;
        RECT 2284.000 2053.640 2284.260 2053.900 ;
        RECT 1410.460 2053.300 1410.720 2053.560 ;
        RECT 2290.900 2053.300 2291.160 2053.560 ;
        RECT 1413.220 2052.960 1413.480 2053.220 ;
        RECT 2304.700 2052.960 2304.960 2053.220 ;
        RECT 1409.540 2052.620 1409.800 2052.880 ;
        RECT 2311.600 2052.620 2311.860 2052.880 ;
        RECT 1409.080 2045.820 1409.340 2046.080 ;
        RECT 1409.540 2034.260 1409.800 2034.520 ;
        RECT 1414.140 2034.260 1414.400 2034.520 ;
        RECT 1414.140 2028.820 1414.400 2029.080 ;
        RECT 1435.760 2028.820 1436.020 2029.080 ;
        RECT 1412.300 2028.140 1412.560 2028.400 ;
        RECT 1414.140 2028.140 1414.400 2028.400 ;
        RECT 1409.080 2027.460 1409.340 2027.720 ;
        RECT 1412.300 2027.460 1412.560 2027.720 ;
        RECT 1410.000 2025.420 1410.260 2025.680 ;
        RECT 1413.220 2025.420 1413.480 2025.680 ;
        RECT 1409.080 2021.340 1409.340 2021.600 ;
        RECT 1421.960 2021.340 1422.220 2021.600 ;
        RECT 1413.220 2014.540 1413.480 2014.800 ;
        RECT 1414.600 2014.540 1414.860 2014.800 ;
        RECT 1414.140 1995.840 1414.400 1996.100 ;
        RECT 1436.220 1995.840 1436.480 1996.100 ;
        RECT 1414.140 1989.380 1414.400 1989.640 ;
        RECT 1436.680 1989.380 1436.940 1989.640 ;
        RECT 1414.140 1984.280 1414.400 1984.540 ;
        RECT 1437.140 1984.280 1437.400 1984.540 ;
        RECT 1414.140 1981.220 1414.400 1981.480 ;
        RECT 1437.600 1981.220 1437.860 1981.480 ;
        RECT 1414.140 1973.740 1414.400 1974.000 ;
        RECT 1438.060 1973.740 1438.320 1974.000 ;
        RECT 1414.140 1969.320 1414.400 1969.580 ;
        RECT 1441.740 1969.320 1442.000 1969.580 ;
        RECT 1409.540 1962.180 1409.800 1962.440 ;
        RECT 1441.280 1962.180 1441.540 1962.440 ;
        RECT 1414.140 1961.500 1414.400 1961.760 ;
        RECT 1440.820 1961.500 1441.080 1961.760 ;
        RECT 1410.460 1956.400 1410.720 1956.660 ;
        RECT 1428.400 1956.400 1428.660 1956.660 ;
        RECT 1413.680 1951.300 1413.940 1951.560 ;
        RECT 1428.860 1951.300 1429.120 1951.560 ;
        RECT 1413.680 1945.180 1413.940 1945.440 ;
        RECT 1429.780 1945.180 1430.040 1945.440 ;
        RECT 1413.680 1942.800 1413.940 1943.060 ;
        RECT 1430.240 1942.800 1430.500 1943.060 ;
        RECT 1413.680 1936.340 1413.940 1936.600 ;
        RECT 1429.320 1936.340 1429.580 1936.600 ;
        RECT 1413.680 1930.220 1413.940 1930.480 ;
        RECT 1431.160 1930.220 1431.420 1930.480 ;
        RECT 1413.680 1926.480 1413.940 1926.740 ;
        RECT 1430.700 1926.480 1430.960 1926.740 ;
        RECT 1414.140 1915.260 1414.400 1915.520 ;
        RECT 1434.840 1915.260 1435.100 1915.520 ;
        RECT 1414.140 1906.420 1414.400 1906.680 ;
        RECT 1434.380 1906.420 1434.640 1906.680 ;
        RECT 1408.620 1895.200 1408.880 1895.460 ;
        RECT 1416.440 1895.200 1416.700 1895.460 ;
        RECT 1414.140 1890.100 1414.400 1890.360 ;
        RECT 1433.460 1890.100 1433.720 1890.360 ;
        RECT 1414.140 1885.680 1414.400 1885.940 ;
        RECT 1433.920 1885.680 1434.180 1885.940 ;
        RECT 1414.140 1881.600 1414.400 1881.860 ;
        RECT 1433.000 1881.600 1433.260 1881.860 ;
        RECT 1414.140 1872.420 1414.400 1872.680 ;
        RECT 1440.360 1872.420 1440.620 1872.680 ;
        RECT 1410.460 1869.700 1410.720 1869.960 ;
        RECT 1413.220 1869.700 1413.480 1869.960 ;
        RECT 1413.680 1869.700 1413.940 1869.960 ;
        RECT 1494.640 1869.700 1494.900 1869.960 ;
        RECT 1414.140 1865.620 1414.400 1865.880 ;
        RECT 1439.440 1865.620 1439.700 1865.880 ;
        RECT 1414.140 1858.140 1414.400 1858.400 ;
        RECT 1439.900 1858.140 1440.160 1858.400 ;
        RECT 1414.140 1855.760 1414.400 1856.020 ;
        RECT 1549.840 1855.760 1550.100 1856.020 ;
        RECT 1413.680 1855.420 1413.940 1855.680 ;
        RECT 1549.380 1855.420 1549.640 1855.680 ;
        RECT 1414.140 1848.960 1414.400 1849.220 ;
        RECT 1548.920 1848.960 1549.180 1849.220 ;
        RECT 1414.140 1840.800 1414.400 1841.060 ;
        RECT 1432.540 1840.800 1432.800 1841.060 ;
        RECT 1414.140 1835.020 1414.400 1835.280 ;
        RECT 1466.120 1835.020 1466.380 1835.280 ;
        RECT 1414.140 1830.940 1414.400 1831.200 ;
        RECT 1432.080 1830.940 1432.340 1831.200 ;
        RECT 1408.620 1826.860 1408.880 1827.120 ;
        RECT 1420.580 1826.860 1420.840 1827.120 ;
        RECT 1410.460 1821.760 1410.720 1822.020 ;
        RECT 1413.220 1821.760 1413.480 1822.020 ;
        RECT 1408.620 1819.380 1408.880 1819.640 ;
        RECT 1416.900 1819.380 1417.160 1819.640 ;
        RECT 1408.620 1813.940 1408.880 1814.200 ;
        RECT 1419.660 1813.940 1419.920 1814.200 ;
        RECT 1408.620 1809.180 1408.880 1809.440 ;
        RECT 1420.120 1809.180 1420.380 1809.440 ;
        RECT 1414.140 1807.480 1414.400 1807.740 ;
        RECT 1494.180 1807.480 1494.440 1807.740 ;
        RECT 1409.080 1799.660 1409.340 1799.920 ;
        RECT 1422.420 1799.660 1422.680 1799.920 ;
        RECT 1408.620 1798.980 1408.880 1799.240 ;
        RECT 1417.360 1798.980 1417.620 1799.240 ;
        RECT 1414.140 1783.000 1414.400 1783.260 ;
        RECT 1438.980 1783.000 1439.240 1783.260 ;
        RECT 1408.620 1778.580 1408.880 1778.840 ;
        RECT 1419.200 1778.580 1419.460 1778.840 ;
        RECT 1408.620 1777.900 1408.880 1778.160 ;
        RECT 1421.040 1777.900 1421.300 1778.160 ;
        RECT 1408.620 1769.400 1408.880 1769.660 ;
        RECT 1418.740 1769.400 1419.000 1769.660 ;
        RECT 1408.620 1764.980 1408.880 1765.240 ;
        RECT 1418.280 1764.980 1418.540 1765.240 ;
        RECT 1408.620 1756.480 1408.880 1756.740 ;
        RECT 1417.820 1756.480 1418.080 1756.740 ;
        RECT 1414.140 1745.260 1414.400 1745.520 ;
        RECT 1473.020 1745.260 1473.280 1745.520 ;
        RECT 1414.140 1738.460 1414.400 1738.720 ;
        RECT 1459.220 1738.460 1459.480 1738.720 ;
        RECT 1410.000 1738.120 1410.260 1738.380 ;
        RECT 1452.320 1738.120 1452.580 1738.380 ;
        RECT 1414.140 1728.940 1414.400 1729.200 ;
        RECT 1438.520 1728.940 1438.780 1729.200 ;
        RECT 1413.680 1723.500 1413.940 1723.760 ;
        RECT 1431.620 1723.500 1431.880 1723.760 ;
        RECT 1410.000 1717.720 1410.260 1717.980 ;
        RECT 1473.480 1717.720 1473.740 1717.980 ;
        RECT 1410.460 1717.380 1410.720 1717.640 ;
        RECT 1424.720 1717.380 1424.980 1717.640 ;
        RECT 1414.140 1710.920 1414.400 1711.180 ;
        RECT 1493.720 1710.920 1493.980 1711.180 ;
        RECT 1409.540 1703.100 1409.800 1703.360 ;
        RECT 1423.340 1703.100 1423.600 1703.360 ;
        RECT 1409.080 1699.360 1409.340 1699.620 ;
        RECT 1422.880 1699.360 1423.140 1699.620 ;
        RECT 1409.540 1694.600 1409.800 1694.860 ;
        RECT 1423.800 1694.600 1424.060 1694.860 ;
        RECT 1409.540 1688.140 1409.800 1688.400 ;
        RECT 1424.260 1688.140 1424.520 1688.400 ;
        RECT 1411.840 1682.700 1412.100 1682.960 ;
        RECT 1427.480 1682.700 1427.740 1682.960 ;
        RECT 1411.840 1677.940 1412.100 1678.200 ;
        RECT 1427.940 1677.940 1428.200 1678.200 ;
        RECT 1410.460 1672.840 1410.720 1673.100 ;
        RECT 1427.020 1672.840 1427.280 1673.100 ;
        RECT 1411.840 1669.440 1412.100 1669.700 ;
        RECT 1459.680 1669.440 1459.940 1669.700 ;
        RECT 1409.540 1668.420 1409.800 1668.680 ;
        RECT 1426.560 1668.420 1426.820 1668.680 ;
        RECT 1414.140 1655.840 1414.400 1656.100 ;
        RECT 1460.140 1655.840 1460.400 1656.100 ;
        RECT 1410.460 1648.020 1410.720 1648.280 ;
        RECT 1425.640 1648.020 1425.900 1648.280 ;
        RECT 1409.540 1647.340 1409.800 1647.600 ;
        RECT 1425.180 1647.340 1425.440 1647.600 ;
        RECT 1410.460 1635.100 1410.720 1635.360 ;
        RECT 1426.100 1635.100 1426.360 1635.360 ;
      LAYER met2 ;
        RECT 1890.700 3266.730 1890.960 3267.050 ;
        RECT 1917.840 3266.730 1918.100 3267.050 ;
        RECT 2542.060 3266.730 2542.320 3267.050 ;
        RECT 1890.760 3264.670 1890.900 3266.730 ;
        RECT 1917.900 3264.670 1918.040 3266.730 ;
        RECT 1890.700 3264.525 1890.960 3264.670 ;
        RECT 1917.840 3264.525 1918.100 3264.670 ;
        RECT 2542.120 3264.525 2542.260 3266.730 ;
        RECT 646.390 3264.155 646.670 3264.525 ;
        RECT 668.010 3264.155 668.290 3264.525 ;
        RECT 1293.150 3264.155 1293.430 3264.525 ;
        RECT 1890.690 3264.155 1890.970 3264.525 ;
        RECT 1917.830 3264.155 1918.110 3264.525 ;
        RECT 2542.050 3264.155 2542.330 3264.525 ;
        RECT 2566.890 3264.155 2567.170 3264.525 ;
        RECT 646.460 3263.990 646.600 3264.155 ;
        RECT 668.080 3263.990 668.220 3264.155 ;
        RECT 1293.220 3263.990 1293.360 3264.155 ;
        RECT 1917.900 3264.025 1918.040 3264.155 ;
        RECT 2542.060 3264.010 2542.320 3264.155 ;
        RECT 2566.900 3264.010 2567.160 3264.155 ;
        RECT 646.400 3263.670 646.660 3263.990 ;
        RECT 668.020 3263.670 668.280 3263.990 ;
        RECT 1293.160 3263.670 1293.420 3263.990 ;
        RECT 1317.540 3263.670 1317.800 3263.990 ;
        RECT 2542.120 3263.855 2542.260 3264.010 ;
        RECT 2594.500 3263.670 2594.760 3263.990 ;
        RECT 697.000 3262.990 697.260 3263.310 ;
        RECT 688.260 3251.770 688.520 3252.090 ;
        RECT 289.430 3230.155 289.710 3230.525 ;
        RECT 288.970 3224.715 289.250 3225.085 ;
        RECT 288.510 3215.875 288.790 3216.245 ;
        RECT 288.050 3209.755 288.330 3210.125 ;
        RECT 287.590 3201.595 287.870 3201.965 ;
        RECT 287.130 3196.155 287.410 3196.525 ;
        RECT 286.670 3187.995 286.950 3188.365 ;
        RECT 286.210 2898.315 286.490 2898.685 ;
        RECT 286.280 2716.590 286.420 2898.315 ;
        RECT 286.220 2716.270 286.480 2716.590 ;
        RECT 286.740 2715.570 286.880 3187.995 ;
        RECT 287.200 2720.670 287.340 3196.155 ;
        RECT 287.660 2721.010 287.800 3201.595 ;
        RECT 288.120 2721.350 288.260 3209.755 ;
        RECT 288.580 2721.690 288.720 3215.875 ;
        RECT 289.040 2725.430 289.180 3224.715 ;
        RECT 288.980 2725.110 289.240 2725.430 ;
        RECT 289.500 2725.090 289.640 3230.155 ;
      LAYER met2 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met2 ;
        RECT 688.320 3248.600 688.460 3251.770 ;
        RECT 688.250 3248.230 688.530 3248.600 ;
        RECT 697.060 2948.325 697.200 3262.990 ;
        RECT 1317.600 3258.405 1317.740 3263.670 ;
        RECT 1317.530 3258.035 1317.810 3258.405 ;
        RECT 1332.260 3252.450 1332.520 3252.770 ;
        RECT 869.040 3251.770 869.300 3252.090 ;
        RECT 869.100 3251.605 869.240 3251.770 ;
        RECT 821.190 3251.235 821.470 3251.605 ;
        RECT 869.030 3251.235 869.310 3251.605 ;
        RECT 1332.320 3251.410 1332.460 3252.450 ;
        RECT 1414.140 3252.110 1414.400 3252.430 ;
        RECT 2582.080 3252.110 2582.340 3252.430 ;
        RECT 821.200 3251.090 821.460 3251.235 ;
        RECT 941.710 3230.155 941.990 3230.525 ;
        RECT 696.990 2947.955 697.270 2948.325 ;
        RECT 927.920 2898.170 928.180 2898.490 ;
        RECT 939.410 2898.315 939.690 2898.685 ;
        RECT 939.420 2898.170 939.680 2898.315 ;
        RECT 337.730 2794.275 338.010 2794.645 ;
        RECT 344.630 2794.275 344.910 2794.645 ;
        RECT 351.530 2794.275 351.810 2794.645 ;
        RECT 358.430 2794.275 358.710 2794.645 ;
        RECT 362.110 2794.275 362.390 2794.645 ;
        RECT 365.330 2794.275 365.610 2794.645 ;
        RECT 368.550 2794.275 368.830 2794.645 ;
        RECT 371.310 2794.275 371.590 2794.645 ;
        RECT 374.990 2794.275 375.270 2794.645 ;
        RECT 378.670 2794.275 378.950 2794.645 ;
        RECT 380.050 2794.275 380.330 2794.645 ;
        RECT 384.650 2794.275 384.930 2794.645 ;
        RECT 386.950 2794.275 387.230 2794.645 ;
        RECT 390.630 2794.275 390.910 2794.645 ;
        RECT 392.470 2794.275 392.750 2794.645 ;
        RECT 396.610 2794.275 396.890 2794.645 ;
        RECT 399.830 2794.275 400.110 2794.645 ;
        RECT 403.970 2794.275 404.250 2794.645 ;
        RECT 406.270 2794.275 406.550 2794.645 ;
        RECT 409.950 2794.275 410.230 2794.645 ;
        RECT 413.630 2794.275 413.910 2794.645 ;
        RECT 414.550 2794.275 414.830 2794.645 ;
        RECT 418.690 2794.275 418.970 2794.645 ;
        RECT 420.990 2794.275 421.270 2794.645 ;
        RECT 427.430 2794.275 427.710 2794.645 ;
        RECT 432.030 2794.275 432.310 2794.645 ;
        RECT 289.440 2724.770 289.700 2725.090 ;
        RECT 288.520 2721.370 288.780 2721.690 ;
        RECT 288.060 2721.030 288.320 2721.350 ;
        RECT 287.600 2720.690 287.860 2721.010 ;
        RECT 287.140 2720.350 287.400 2720.670 ;
        RECT 315.200 2716.610 315.460 2716.930 ;
        RECT 286.680 2715.250 286.940 2715.570 ;
        RECT 305.070 2714.715 305.350 2715.085 ;
        RECT 305.140 2700.000 305.280 2714.715 ;
        RECT 315.260 2700.000 315.400 2716.610 ;
        RECT 335.900 2715.930 336.160 2716.250 ;
        RECT 325.780 2714.570 326.040 2714.890 ;
        RECT 325.840 2700.000 325.980 2714.570 ;
        RECT 335.960 2700.000 336.100 2715.930 ;
        RECT 337.800 2715.910 337.940 2794.275 ;
        RECT 337.740 2715.590 338.000 2715.910 ;
        RECT 344.700 2712.250 344.840 2794.275 ;
        RECT 351.070 2792.235 351.350 2792.605 ;
        RECT 351.140 2717.950 351.280 2792.235 ;
        RECT 351.080 2717.630 351.340 2717.950 ;
        RECT 351.600 2714.210 351.740 2794.275 ;
        RECT 358.500 2718.630 358.640 2794.275 ;
        RECT 362.180 2791.390 362.320 2794.275 ;
        RECT 362.120 2791.070 362.380 2791.390 ;
        RECT 365.400 2731.890 365.540 2794.275 ;
        RECT 368.620 2792.070 368.760 2794.275 ;
        RECT 368.560 2791.750 368.820 2792.070 ;
        RECT 371.380 2791.050 371.520 2794.275 ;
        RECT 375.060 2793.770 375.200 2794.275 ;
        RECT 375.000 2793.450 375.260 2793.770 ;
        RECT 371.320 2790.730 371.580 2791.050 ;
        RECT 378.740 2788.330 378.880 2794.275 ;
        RECT 380.120 2793.430 380.260 2794.275 ;
        RECT 380.060 2793.110 380.320 2793.430 ;
        RECT 384.720 2790.710 384.860 2794.275 ;
        RECT 386.960 2794.130 387.220 2794.275 ;
        RECT 384.660 2790.390 384.920 2790.710 ;
        RECT 378.680 2788.010 378.940 2788.330 ;
        RECT 390.700 2787.990 390.840 2794.275 ;
        RECT 392.540 2792.410 392.680 2794.275 ;
        RECT 392.480 2792.090 392.740 2792.410 ;
        RECT 396.680 2790.370 396.820 2794.275 ;
        RECT 397.070 2793.595 397.350 2793.965 ;
        RECT 397.140 2792.750 397.280 2793.595 ;
        RECT 397.080 2792.430 397.340 2792.750 ;
        RECT 396.620 2790.050 396.880 2790.370 ;
        RECT 399.900 2788.670 400.040 2794.275 ;
        RECT 404.040 2791.730 404.180 2794.275 ;
        RECT 403.980 2791.410 404.240 2791.730 ;
        RECT 406.340 2790.030 406.480 2794.275 ;
        RECT 410.020 2793.090 410.160 2794.275 ;
        RECT 409.960 2792.770 410.220 2793.090 ;
        RECT 410.410 2790.875 410.690 2791.245 ;
        RECT 406.280 2789.710 406.540 2790.030 ;
        RECT 399.840 2788.350 400.100 2788.670 ;
        RECT 390.640 2787.670 390.900 2787.990 ;
        RECT 365.340 2731.570 365.600 2731.890 ;
        RECT 408.580 2721.710 408.840 2722.030 ;
        RECT 358.440 2718.310 358.700 2718.630 ;
        RECT 377.300 2718.310 377.560 2718.630 ;
        RECT 356.600 2717.630 356.860 2717.950 ;
        RECT 351.540 2713.890 351.800 2714.210 ;
        RECT 344.700 2712.110 345.300 2712.250 ;
        RECT 345.160 2700.010 345.300 2712.110 ;
        RECT 345.160 2700.000 346.610 2700.010 ;
        RECT 356.660 2700.000 356.800 2717.630 ;
        RECT 367.180 2713.890 367.440 2714.210 ;
        RECT 367.240 2700.000 367.380 2713.890 ;
        RECT 377.360 2700.000 377.500 2718.310 ;
        RECT 398.460 2716.270 398.720 2716.590 ;
        RECT 387.880 2714.910 388.140 2715.230 ;
        RECT 387.940 2700.000 388.080 2714.910 ;
        RECT 398.520 2700.000 398.660 2716.270 ;
        RECT 408.640 2700.000 408.780 2721.710 ;
        RECT 410.480 2716.930 410.620 2790.875 ;
        RECT 413.700 2789.010 413.840 2794.275 ;
        RECT 414.620 2791.390 414.760 2794.275 ;
        RECT 414.560 2791.070 414.820 2791.390 ;
        RECT 418.760 2789.350 418.900 2794.275 ;
        RECT 421.060 2793.770 421.200 2794.275 ;
        RECT 421.000 2793.450 421.260 2793.770 ;
        RECT 426.970 2793.595 427.250 2793.965 ;
        RECT 427.040 2793.430 427.180 2793.595 ;
        RECT 426.980 2793.110 427.240 2793.430 ;
        RECT 418.700 2789.030 418.960 2789.350 ;
        RECT 413.640 2788.690 413.900 2789.010 ;
        RECT 424.220 2788.010 424.480 2788.330 ;
        RECT 419.160 2722.050 419.420 2722.370 ;
        RECT 410.420 2716.610 410.680 2716.930 ;
        RECT 419.220 2700.000 419.360 2722.050 ;
        RECT 424.280 2713.530 424.420 2788.010 ;
        RECT 427.500 2731.550 427.640 2794.275 ;
        RECT 432.040 2794.130 432.300 2794.275 ;
        RECT 433.420 2794.130 433.680 2794.450 ;
        RECT 434.330 2794.275 434.610 2794.645 ;
        RECT 439.390 2794.275 439.670 2794.645 ;
        RECT 441.230 2794.275 441.510 2794.645 ;
        RECT 444.450 2794.275 444.730 2794.645 ;
        RECT 448.130 2794.275 448.410 2794.645 ;
        RECT 450.430 2794.275 450.710 2794.645 ;
        RECT 455.030 2794.275 455.310 2794.645 ;
        RECT 461.930 2794.275 462.210 2794.645 ;
        RECT 466.530 2794.275 466.810 2794.645 ;
        RECT 468.370 2794.275 468.650 2794.645 ;
        RECT 475.730 2794.275 476.010 2794.645 ;
        RECT 478.490 2794.275 478.770 2794.645 ;
        RECT 482.630 2794.275 482.910 2794.645 ;
        RECT 484.930 2794.275 485.210 2794.645 ;
        RECT 489.070 2794.275 489.350 2794.645 ;
        RECT 492.750 2794.275 493.030 2794.645 ;
        RECT 496.430 2794.275 496.710 2794.645 ;
        RECT 433.480 2792.070 433.620 2794.130 ;
        RECT 433.870 2793.595 434.150 2793.965 ;
        RECT 433.420 2791.750 433.680 2792.070 ;
        RECT 431.120 2787.670 431.380 2787.990 ;
        RECT 427.440 2731.230 427.700 2731.550 ;
        RECT 429.280 2722.390 429.540 2722.710 ;
        RECT 424.220 2713.210 424.480 2713.530 ;
        RECT 429.340 2700.000 429.480 2722.390 ;
        RECT 431.180 2713.870 431.320 2787.670 ;
        RECT 433.940 2731.210 434.080 2793.595 ;
        RECT 433.880 2730.890 434.140 2731.210 ;
        RECT 434.400 2730.870 434.540 2794.275 ;
        RECT 439.460 2792.410 439.600 2794.275 ;
        RECT 439.400 2792.090 439.660 2792.410 ;
        RECT 434.340 2730.550 434.600 2730.870 ;
        RECT 441.300 2730.530 441.440 2794.275 ;
        RECT 444.520 2792.750 444.660 2794.275 ;
        RECT 444.460 2792.430 444.720 2792.750 ;
        RECT 444.920 2788.350 445.180 2788.670 ;
        RECT 441.240 2730.210 441.500 2730.530 ;
        RECT 439.860 2722.730 440.120 2723.050 ;
        RECT 431.120 2713.550 431.380 2713.870 ;
        RECT 439.920 2700.000 440.060 2722.730 ;
        RECT 444.980 2714.550 445.120 2788.350 ;
        RECT 448.200 2729.850 448.340 2794.275 ;
        RECT 450.500 2791.730 450.640 2794.275 ;
        RECT 450.440 2791.410 450.700 2791.730 ;
        RECT 455.100 2730.190 455.240 2794.275 ;
        RECT 455.490 2793.595 455.770 2793.965 ;
        RECT 455.560 2793.090 455.700 2793.595 ;
        RECT 455.500 2792.770 455.760 2793.090 ;
        RECT 455.560 2788.330 455.700 2792.770 ;
        RECT 455.500 2788.010 455.760 2788.330 ;
        RECT 455.040 2729.870 455.300 2730.190 ;
        RECT 448.140 2729.530 448.400 2729.850 ;
        RECT 462.000 2729.510 462.140 2794.275 ;
        RECT 462.400 2793.965 462.660 2794.110 ;
        RECT 462.390 2793.595 462.670 2793.965 ;
        RECT 466.600 2793.770 466.740 2794.275 ;
        RECT 462.460 2791.390 462.600 2793.595 ;
        RECT 466.540 2793.450 466.800 2793.770 ;
        RECT 462.400 2791.070 462.660 2791.390 ;
        RECT 465.620 2788.690 465.880 2789.010 ;
        RECT 461.940 2729.190 462.200 2729.510 ;
        RECT 460.560 2723.410 460.820 2723.730 ;
        RECT 449.980 2723.070 450.240 2723.390 ;
        RECT 444.920 2714.230 445.180 2714.550 ;
        RECT 450.040 2700.000 450.180 2723.070 ;
        RECT 460.620 2700.000 460.760 2723.410 ;
        RECT 465.680 2714.210 465.820 2788.690 ;
        RECT 468.440 2728.830 468.580 2794.275 ;
        RECT 468.830 2793.595 469.110 2793.965 ;
        RECT 475.270 2793.595 475.550 2793.965 ;
        RECT 468.900 2729.170 469.040 2793.595 ;
        RECT 475.340 2793.430 475.480 2793.595 ;
        RECT 475.280 2793.110 475.540 2793.430 ;
        RECT 475.340 2789.010 475.480 2793.110 ;
        RECT 475.280 2788.690 475.540 2789.010 ;
        RECT 468.840 2728.850 469.100 2729.170 ;
        RECT 468.380 2728.510 468.640 2728.830 ;
        RECT 475.800 2724.750 475.940 2794.275 ;
        RECT 478.560 2792.070 478.700 2794.275 ;
        RECT 482.640 2794.130 482.900 2794.275 ;
        RECT 478.500 2791.750 478.760 2792.070 ;
        RECT 485.000 2789.690 485.140 2794.275 ;
        RECT 489.140 2791.390 489.280 2794.275 ;
        RECT 492.820 2792.750 492.960 2794.275 ;
        RECT 492.760 2792.430 493.020 2792.750 ;
        RECT 489.080 2791.070 489.340 2791.390 ;
        RECT 484.940 2789.370 485.200 2789.690 ;
        RECT 479.420 2787.670 479.680 2787.990 ;
        RECT 475.740 2724.430 476.000 2724.750 ;
        RECT 470.680 2723.750 470.940 2724.070 ;
        RECT 465.620 2713.890 465.880 2714.210 ;
        RECT 470.740 2700.000 470.880 2723.750 ;
        RECT 479.480 2716.250 479.620 2787.670 ;
        RECT 481.260 2724.090 481.520 2724.410 ;
        RECT 479.420 2715.930 479.680 2716.250 ;
        RECT 481.320 2700.000 481.460 2724.090 ;
        RECT 496.500 2716.930 496.640 2794.275 ;
        RECT 500.580 2794.130 500.840 2794.450 ;
        RECT 501.950 2794.275 502.230 2794.645 ;
        RECT 509.770 2794.275 510.050 2794.645 ;
        RECT 513.910 2794.275 514.190 2794.645 ;
        RECT 517.130 2794.275 517.410 2794.645 ;
        RECT 524.030 2794.275 524.310 2794.645 ;
        RECT 526.790 2794.275 527.070 2794.645 ;
        RECT 530.930 2794.275 531.210 2794.645 ;
        RECT 537.370 2794.275 537.650 2794.645 ;
        RECT 539.210 2794.275 539.490 2794.645 ;
        RECT 544.270 2794.275 544.550 2794.645 ;
        RECT 551.630 2794.275 551.910 2794.645 ;
        RECT 500.110 2792.915 500.390 2793.285 ;
        RECT 500.180 2788.330 500.320 2792.915 ;
        RECT 500.120 2788.010 500.380 2788.330 ;
        RECT 496.440 2716.610 496.700 2716.930 ;
        RECT 491.840 2715.590 492.100 2715.910 ;
        RECT 491.900 2700.000 492.040 2715.590 ;
        RECT 500.180 2712.170 500.320 2788.010 ;
        RECT 500.640 2717.270 500.780 2794.130 ;
        RECT 501.030 2793.595 501.310 2793.965 ;
        RECT 501.100 2791.730 501.240 2793.595 ;
        RECT 502.020 2791.730 502.160 2794.275 ;
        RECT 503.800 2793.790 504.060 2794.110 ;
        RECT 503.860 2793.430 504.000 2793.790 ;
        RECT 508.850 2793.595 509.130 2793.965 ;
        RECT 508.920 2793.430 509.060 2793.595 ;
        RECT 503.800 2793.110 504.060 2793.430 ;
        RECT 508.860 2793.110 509.120 2793.430 ;
        RECT 501.040 2791.410 501.300 2791.730 ;
        RECT 501.960 2791.410 502.220 2791.730 ;
        RECT 501.100 2788.330 501.240 2791.410 ;
        RECT 501.040 2788.010 501.300 2788.330 ;
        RECT 500.580 2716.950 500.840 2717.270 ;
        RECT 509.840 2716.590 509.980 2794.275 ;
        RECT 513.980 2794.110 514.120 2794.275 ;
        RECT 510.230 2793.595 510.510 2793.965 ;
        RECT 513.920 2793.790 514.180 2794.110 ;
        RECT 510.300 2792.070 510.440 2793.595 ;
        RECT 510.240 2791.750 510.500 2792.070 ;
        RECT 512.540 2720.350 512.800 2720.670 ;
        RECT 509.780 2716.270 510.040 2716.590 ;
        RECT 501.960 2715.250 502.220 2715.570 ;
        RECT 500.120 2711.850 500.380 2712.170 ;
        RECT 502.020 2700.000 502.160 2715.250 ;
        RECT 512.600 2700.000 512.740 2720.350 ;
        RECT 517.200 2716.250 517.340 2794.275 ;
        RECT 520.810 2792.915 521.090 2793.285 ;
        RECT 520.880 2789.010 521.020 2792.915 ;
        RECT 524.100 2792.410 524.240 2794.275 ;
        RECT 526.860 2793.770 527.000 2794.275 ;
        RECT 526.800 2793.450 527.060 2793.770 ;
        RECT 524.040 2792.090 524.300 2792.410 ;
        RECT 520.820 2788.690 521.080 2789.010 ;
        RECT 517.140 2715.930 517.400 2716.250 ;
        RECT 520.880 2712.510 521.020 2788.690 ;
        RECT 522.660 2720.690 522.920 2721.010 ;
        RECT 520.820 2712.190 521.080 2712.510 ;
        RECT 522.720 2700.000 522.860 2720.690 ;
        RECT 531.000 2715.910 531.140 2794.275 ;
        RECT 534.610 2793.595 534.890 2793.965 ;
        RECT 534.680 2789.690 534.820 2793.595 ;
        RECT 537.440 2793.090 537.580 2794.275 ;
        RECT 537.380 2792.770 537.640 2793.090 ;
        RECT 539.280 2792.750 539.420 2794.275 ;
        RECT 541.510 2792.915 541.790 2793.285 ;
        RECT 539.220 2792.430 539.480 2792.750 ;
        RECT 539.280 2789.690 539.420 2792.430 ;
        RECT 534.620 2789.370 534.880 2789.690 ;
        RECT 539.220 2789.370 539.480 2789.690 ;
        RECT 533.240 2721.030 533.500 2721.350 ;
        RECT 530.940 2715.590 531.200 2715.910 ;
        RECT 533.300 2700.000 533.440 2721.030 ;
        RECT 534.680 2712.850 534.820 2789.370 ;
        RECT 541.580 2788.330 541.720 2792.915 ;
        RECT 544.340 2792.750 544.480 2794.275 ;
        RECT 544.280 2792.430 544.540 2792.750 ;
        RECT 541.520 2788.010 541.780 2788.330 ;
        RECT 541.580 2713.190 541.720 2788.010 ;
        RECT 543.360 2721.370 543.620 2721.690 ;
        RECT 541.520 2712.870 541.780 2713.190 ;
        RECT 534.620 2712.530 534.880 2712.850 ;
        RECT 543.420 2700.000 543.560 2721.370 ;
        RECT 551.700 2715.570 551.840 2794.275 ;
        RECT 648.240 2794.130 648.500 2794.450 ;
        RECT 627.540 2788.690 627.800 2789.010 ;
        RECT 606.840 2788.350 607.100 2788.670 ;
        RECT 586.140 2788.010 586.400 2788.330 ;
        RECT 553.940 2725.110 554.200 2725.430 ;
        RECT 551.640 2715.250 551.900 2715.570 ;
        RECT 554.000 2700.000 554.140 2725.110 ;
        RECT 564.060 2724.770 564.320 2725.090 ;
        RECT 564.120 2700.000 564.260 2724.770 ;
        RECT 574.640 2717.290 574.900 2717.610 ;
        RECT 574.700 2700.000 574.840 2717.290 ;
        RECT 586.200 2700.010 586.340 2788.010 ;
        RECT 595.340 2717.630 595.600 2717.950 ;
        RECT 585.350 2700.000 586.340 2700.010 ;
        RECT 595.400 2700.000 595.540 2717.630 ;
        RECT 606.900 2700.010 607.040 2788.350 ;
        RECT 616.040 2717.970 616.300 2718.290 ;
        RECT 606.050 2700.000 607.040 2700.010 ;
        RECT 616.100 2700.000 616.240 2717.970 ;
        RECT 627.600 2700.010 627.740 2788.690 ;
        RECT 636.740 2718.310 637.000 2718.630 ;
        RECT 626.750 2700.000 627.740 2700.010 ;
        RECT 636.800 2700.000 636.940 2718.310 ;
        RECT 648.300 2700.010 648.440 2794.130 ;
        RECT 676.300 2793.790 676.560 2794.110 ;
        RECT 662.500 2793.110 662.760 2793.430 ;
        RECT 657.440 2711.850 657.700 2712.170 ;
        RECT 647.450 2700.000 648.440 2700.010 ;
        RECT 657.500 2700.000 657.640 2711.850 ;
      LAYER met2 ;
        RECT 300.030 2695.720 304.800 2697.365 ;
      LAYER met2 ;
        RECT 305.080 2696.000 305.360 2700.000 ;
      LAYER met2 ;
        RECT 305.640 2695.720 314.920 2697.365 ;
      LAYER met2 ;
        RECT 315.200 2696.000 315.480 2700.000 ;
      LAYER met2 ;
        RECT 315.760 2695.720 325.500 2697.365 ;
      LAYER met2 ;
        RECT 325.780 2696.000 326.060 2700.000 ;
      LAYER met2 ;
        RECT 326.340 2695.720 335.620 2697.365 ;
      LAYER met2 ;
        RECT 335.900 2696.000 336.180 2700.000 ;
        RECT 345.160 2699.870 346.760 2700.000 ;
      LAYER met2 ;
        RECT 336.460 2695.720 346.200 2697.365 ;
      LAYER met2 ;
        RECT 346.480 2696.000 346.760 2699.870 ;
      LAYER met2 ;
        RECT 347.040 2695.720 356.320 2697.365 ;
      LAYER met2 ;
        RECT 356.600 2696.000 356.880 2700.000 ;
      LAYER met2 ;
        RECT 357.160 2695.720 366.900 2697.365 ;
      LAYER met2 ;
        RECT 367.180 2696.000 367.460 2700.000 ;
      LAYER met2 ;
        RECT 367.740 2695.720 377.020 2697.365 ;
      LAYER met2 ;
        RECT 377.300 2696.000 377.580 2700.000 ;
      LAYER met2 ;
        RECT 377.860 2695.720 387.600 2697.365 ;
      LAYER met2 ;
        RECT 387.880 2696.000 388.160 2700.000 ;
      LAYER met2 ;
        RECT 388.440 2695.720 398.180 2697.365 ;
      LAYER met2 ;
        RECT 398.460 2696.000 398.740 2700.000 ;
      LAYER met2 ;
        RECT 399.020 2695.720 408.300 2697.365 ;
      LAYER met2 ;
        RECT 408.580 2696.000 408.860 2700.000 ;
      LAYER met2 ;
        RECT 409.140 2695.720 418.880 2697.365 ;
      LAYER met2 ;
        RECT 419.160 2696.000 419.440 2700.000 ;
      LAYER met2 ;
        RECT 419.720 2695.720 429.000 2697.365 ;
      LAYER met2 ;
        RECT 429.280 2696.000 429.560 2700.000 ;
      LAYER met2 ;
        RECT 429.840 2695.720 439.580 2697.365 ;
      LAYER met2 ;
        RECT 439.860 2696.000 440.140 2700.000 ;
      LAYER met2 ;
        RECT 440.420 2695.720 449.700 2697.365 ;
      LAYER met2 ;
        RECT 449.980 2696.000 450.260 2700.000 ;
      LAYER met2 ;
        RECT 450.540 2695.720 460.280 2697.365 ;
      LAYER met2 ;
        RECT 460.560 2696.000 460.840 2700.000 ;
      LAYER met2 ;
        RECT 461.120 2695.720 470.400 2697.365 ;
      LAYER met2 ;
        RECT 470.680 2696.000 470.960 2700.000 ;
      LAYER met2 ;
        RECT 471.240 2695.720 480.980 2697.365 ;
      LAYER met2 ;
        RECT 481.260 2696.000 481.540 2700.000 ;
      LAYER met2 ;
        RECT 481.820 2695.720 491.560 2697.365 ;
      LAYER met2 ;
        RECT 491.840 2696.000 492.120 2700.000 ;
      LAYER met2 ;
        RECT 492.400 2695.720 501.680 2697.365 ;
      LAYER met2 ;
        RECT 501.960 2696.000 502.240 2700.000 ;
      LAYER met2 ;
        RECT 502.520 2695.720 512.260 2697.365 ;
      LAYER met2 ;
        RECT 512.540 2696.000 512.820 2700.000 ;
      LAYER met2 ;
        RECT 513.100 2695.720 522.380 2697.365 ;
      LAYER met2 ;
        RECT 522.660 2696.000 522.940 2700.000 ;
      LAYER met2 ;
        RECT 523.220 2695.720 532.960 2697.365 ;
      LAYER met2 ;
        RECT 533.240 2696.000 533.520 2700.000 ;
      LAYER met2 ;
        RECT 533.800 2695.720 543.080 2697.365 ;
      LAYER met2 ;
        RECT 543.360 2696.000 543.640 2700.000 ;
      LAYER met2 ;
        RECT 543.920 2695.720 553.660 2697.365 ;
      LAYER met2 ;
        RECT 553.940 2696.000 554.220 2700.000 ;
      LAYER met2 ;
        RECT 554.500 2695.720 563.780 2697.365 ;
      LAYER met2 ;
        RECT 564.060 2696.000 564.340 2700.000 ;
      LAYER met2 ;
        RECT 564.620 2695.720 574.360 2697.365 ;
      LAYER met2 ;
        RECT 574.640 2696.000 574.920 2700.000 ;
        RECT 585.220 2699.870 586.340 2700.000 ;
      LAYER met2 ;
        RECT 575.200 2695.720 584.940 2697.365 ;
      LAYER met2 ;
        RECT 585.220 2696.000 585.500 2699.870 ;
      LAYER met2 ;
        RECT 585.780 2695.720 595.060 2697.365 ;
      LAYER met2 ;
        RECT 595.340 2696.000 595.620 2700.000 ;
        RECT 605.920 2699.870 607.040 2700.000 ;
      LAYER met2 ;
        RECT 595.900 2695.720 605.640 2697.365 ;
      LAYER met2 ;
        RECT 605.920 2696.000 606.200 2699.870 ;
      LAYER met2 ;
        RECT 606.480 2695.720 615.760 2697.365 ;
      LAYER met2 ;
        RECT 616.040 2696.000 616.320 2700.000 ;
        RECT 626.620 2699.870 627.740 2700.000 ;
      LAYER met2 ;
        RECT 616.600 2695.720 626.340 2697.365 ;
      LAYER met2 ;
        RECT 626.620 2696.000 626.900 2699.870 ;
      LAYER met2 ;
        RECT 627.180 2695.720 636.460 2697.365 ;
      LAYER met2 ;
        RECT 636.740 2696.000 637.020 2700.000 ;
        RECT 647.320 2699.870 648.440 2700.000 ;
      LAYER met2 ;
        RECT 637.300 2695.720 647.040 2697.365 ;
      LAYER met2 ;
        RECT 647.320 2696.000 647.600 2699.870 ;
      LAYER met2 ;
        RECT 647.880 2695.720 657.160 2697.365 ;
      LAYER met2 ;
        RECT 657.440 2696.000 657.720 2700.000 ;
        RECT 662.560 2699.330 662.700 2793.110 ;
        RECT 668.020 2699.330 668.300 2700.000 ;
        RECT 662.560 2699.190 668.300 2699.330 ;
        RECT 676.360 2699.330 676.500 2793.790 ;
        RECT 697.000 2793.450 697.260 2793.770 ;
        RECT 700.220 2793.450 700.480 2793.770 ;
        RECT 686.420 2793.110 686.680 2793.430 ;
        RECT 686.480 2715.085 686.620 2793.110 ;
        RECT 686.410 2714.715 686.690 2715.085 ;
        RECT 688.720 2712.190 688.980 2712.510 ;
        RECT 688.780 2700.000 688.920 2712.190 ;
        RECT 697.060 2700.010 697.200 2793.450 ;
        RECT 700.280 2714.890 700.420 2793.450 ;
        RECT 865.820 2792.770 866.080 2793.090 ;
        RECT 858.920 2792.090 859.180 2792.410 ;
        RECT 852.020 2791.750 852.280 2792.070 ;
        RECT 845.120 2791.410 845.380 2791.730 ;
        RECT 838.220 2791.070 838.480 2791.390 ;
        RECT 745.300 2790.730 745.560 2791.050 ;
        RECT 717.700 2789.370 717.960 2789.690 ;
        RECT 700.220 2714.570 700.480 2714.890 ;
        RECT 709.420 2712.530 709.680 2712.850 ;
        RECT 697.060 2700.000 699.430 2700.010 ;
        RECT 709.480 2700.000 709.620 2712.530 ;
        RECT 678.600 2699.330 678.880 2700.000 ;
        RECT 676.360 2699.190 678.880 2699.330 ;
      LAYER met2 ;
        RECT 658.000 2695.720 667.740 2697.365 ;
      LAYER met2 ;
        RECT 668.020 2696.000 668.300 2699.190 ;
      LAYER met2 ;
        RECT 668.580 2695.720 678.320 2697.365 ;
      LAYER met2 ;
        RECT 678.600 2696.000 678.880 2699.190 ;
      LAYER met2 ;
        RECT 679.160 2695.720 688.440 2697.365 ;
      LAYER met2 ;
        RECT 688.720 2696.000 689.000 2700.000 ;
        RECT 697.060 2699.870 699.580 2700.000 ;
      LAYER met2 ;
        RECT 689.280 2695.720 699.020 2697.365 ;
      LAYER met2 ;
        RECT 699.300 2696.000 699.580 2699.870 ;
      LAYER met2 ;
        RECT 699.860 2695.720 709.140 2697.365 ;
      LAYER met2 ;
        RECT 709.420 2696.000 709.700 2700.000 ;
        RECT 717.760 2699.330 717.900 2789.370 ;
        RECT 740.700 2731.570 740.960 2731.890 ;
        RECT 730.120 2712.870 730.380 2713.190 ;
        RECT 730.180 2700.000 730.320 2712.870 ;
        RECT 740.760 2700.000 740.900 2731.570 ;
        RECT 720.000 2699.330 720.280 2700.000 ;
        RECT 717.760 2699.190 720.280 2699.330 ;
      LAYER met2 ;
        RECT 709.980 2695.720 719.720 2697.365 ;
      LAYER met2 ;
        RECT 720.000 2696.000 720.280 2699.190 ;
      LAYER met2 ;
        RECT 720.560 2695.720 729.840 2697.365 ;
      LAYER met2 ;
        RECT 730.120 2696.000 730.400 2700.000 ;
      LAYER met2 ;
        RECT 730.680 2695.720 740.420 2697.365 ;
      LAYER met2 ;
        RECT 740.700 2696.000 740.980 2700.000 ;
        RECT 745.360 2699.330 745.500 2790.730 ;
        RECT 766.000 2790.390 766.260 2790.710 ;
        RECT 761.400 2713.210 761.660 2713.530 ;
        RECT 761.460 2700.000 761.600 2713.210 ;
        RECT 766.060 2700.690 766.200 2790.390 ;
        RECT 786.700 2790.050 786.960 2790.370 ;
        RECT 782.100 2713.550 782.360 2713.870 ;
        RECT 766.060 2700.550 769.420 2700.690 ;
        RECT 750.820 2699.330 751.100 2700.000 ;
        RECT 745.360 2699.190 751.100 2699.330 ;
      LAYER met2 ;
        RECT 741.260 2695.720 750.540 2697.365 ;
      LAYER met2 ;
        RECT 750.820 2696.000 751.100 2699.190 ;
      LAYER met2 ;
        RECT 751.380 2695.720 761.120 2697.365 ;
      LAYER met2 ;
        RECT 761.400 2696.000 761.680 2700.000 ;
        RECT 769.280 2699.330 769.420 2700.550 ;
        RECT 782.160 2700.000 782.300 2713.550 ;
        RECT 771.980 2699.330 772.260 2700.000 ;
        RECT 769.280 2699.190 772.260 2699.330 ;
      LAYER met2 ;
        RECT 761.960 2695.720 771.700 2697.365 ;
      LAYER met2 ;
        RECT 771.980 2696.000 772.260 2699.190 ;
      LAYER met2 ;
        RECT 772.540 2695.720 781.820 2697.365 ;
      LAYER met2 ;
        RECT 782.100 2696.000 782.380 2700.000 ;
        RECT 786.760 2699.330 786.900 2790.050 ;
        RECT 807.400 2789.710 807.660 2790.030 ;
        RECT 802.800 2714.230 803.060 2714.550 ;
        RECT 802.860 2700.000 803.000 2714.230 ;
        RECT 807.460 2700.690 807.600 2789.710 ;
        RECT 828.100 2789.030 828.360 2789.350 ;
        RECT 823.500 2713.890 823.760 2714.210 ;
        RECT 807.460 2700.550 811.740 2700.690 ;
        RECT 811.600 2700.010 811.740 2700.550 ;
        RECT 811.600 2700.000 813.510 2700.010 ;
        RECT 823.560 2700.000 823.700 2713.890 ;
        RECT 828.160 2700.690 828.300 2789.030 ;
        RECT 838.280 2713.190 838.420 2791.070 ;
        RECT 844.200 2731.230 844.460 2731.550 ;
        RECT 838.220 2712.870 838.480 2713.190 ;
        RECT 828.160 2700.550 832.900 2700.690 ;
        RECT 832.760 2700.010 832.900 2700.550 ;
        RECT 832.760 2700.000 834.210 2700.010 ;
        RECT 844.260 2700.000 844.400 2731.230 ;
        RECT 845.180 2713.530 845.320 2791.410 ;
        RECT 852.080 2713.870 852.220 2791.750 ;
        RECT 854.780 2730.890 855.040 2731.210 ;
        RECT 852.020 2713.550 852.280 2713.870 ;
        RECT 845.120 2713.210 845.380 2713.530 ;
        RECT 854.840 2700.000 854.980 2730.890 ;
        RECT 858.980 2714.210 859.120 2792.090 ;
        RECT 865.360 2730.550 865.620 2730.870 ;
        RECT 858.920 2713.890 859.180 2714.210 ;
        RECT 865.420 2700.000 865.560 2730.550 ;
        RECT 865.880 2714.550 866.020 2792.770 ;
        RECT 872.720 2792.430 872.980 2792.750 ;
        RECT 872.780 2714.890 872.920 2792.430 ;
        RECT 875.480 2730.210 875.740 2730.530 ;
        RECT 872.720 2714.570 872.980 2714.890 ;
        RECT 865.820 2714.230 866.080 2714.550 ;
        RECT 875.540 2700.000 875.680 2730.210 ;
        RECT 896.180 2729.870 896.440 2730.190 ;
        RECT 886.060 2729.530 886.320 2729.850 ;
        RECT 886.120 2700.000 886.260 2729.530 ;
        RECT 896.240 2700.000 896.380 2729.870 ;
        RECT 906.760 2729.190 907.020 2729.510 ;
        RECT 906.820 2700.000 906.960 2729.190 ;
        RECT 916.880 2728.850 917.140 2729.170 ;
        RECT 916.940 2700.000 917.080 2728.850 ;
        RECT 927.460 2728.510 927.720 2728.830 ;
        RECT 927.520 2700.000 927.660 2728.510 ;
        RECT 927.980 2715.230 928.120 2898.170 ;
        RECT 937.580 2724.430 937.840 2724.750 ;
        RECT 927.920 2714.910 928.180 2715.230 ;
        RECT 937.640 2700.000 937.780 2724.430 ;
        RECT 941.780 2724.410 941.920 3230.155 ;
        RECT 942.170 3224.715 942.450 3225.085 ;
        RECT 941.720 2724.090 941.980 2724.410 ;
        RECT 942.240 2724.070 942.380 3224.715 ;
        RECT 942.630 3215.875 942.910 3216.245 ;
        RECT 942.180 2723.750 942.440 2724.070 ;
        RECT 942.700 2723.730 942.840 3215.875 ;
        RECT 943.090 3209.755 943.370 3210.125 ;
        RECT 942.640 2723.410 942.900 2723.730 ;
        RECT 943.160 2723.390 943.300 3209.755 ;
        RECT 943.550 3201.595 943.830 3201.965 ;
        RECT 943.100 2723.070 943.360 2723.390 ;
        RECT 943.620 2723.050 943.760 3201.595 ;
        RECT 944.010 3196.155 944.290 3196.525 ;
        RECT 943.560 2722.730 943.820 2723.050 ;
        RECT 944.080 2722.710 944.220 3196.155 ;
        RECT 944.470 3187.995 944.750 3188.365 ;
        RECT 944.020 2722.390 944.280 2722.710 ;
        RECT 944.540 2722.370 944.680 3187.995 ;
      LAYER met2 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met2 ;
        RECT 1332.260 3251.090 1332.520 3251.410 ;
        RECT 1332.320 3249.565 1332.460 3251.090 ;
        RECT 1414.200 3251.070 1414.340 3252.110 ;
        RECT 1407.700 3250.750 1407.960 3251.070 ;
        RECT 1414.140 3250.750 1414.400 3251.070 ;
        RECT 1332.250 3249.195 1332.530 3249.565 ;
        RECT 1345.590 2946.595 1345.870 2946.965 ;
        RECT 1345.660 2936.085 1345.800 2946.595 ;
        RECT 1345.590 2935.715 1345.870 2936.085 ;
        RECT 1352.030 2901.715 1352.310 2902.085 ;
        RECT 1352.100 2901.550 1352.240 2901.715 ;
        RECT 1352.040 2901.230 1352.300 2901.550 ;
        RECT 1397.580 2901.230 1397.840 2901.550 ;
        RECT 1054.870 2799.715 1055.150 2800.085 ;
        RECT 1053.030 2795.635 1053.310 2796.005 ;
        RECT 979.890 2794.275 980.170 2794.645 ;
        RECT 1013.930 2794.275 1014.210 2794.645 ;
        RECT 1018.990 2794.275 1019.270 2794.645 ;
        RECT 1020.830 2794.275 1021.110 2794.645 ;
        RECT 1027.730 2794.275 1028.010 2794.645 ;
        RECT 1034.630 2794.275 1034.910 2794.645 ;
        RECT 1042.450 2794.275 1042.730 2794.645 ;
        RECT 1053.100 2794.450 1053.240 2795.635 ;
        RECT 944.480 2722.050 944.740 2722.370 ;
        RECT 979.960 2722.030 980.100 2794.275 ;
        RECT 986.790 2793.595 987.070 2793.965 ;
        RECT 1001.050 2793.595 1001.330 2793.965 ;
        RECT 986.860 2793.430 987.000 2793.595 ;
        RECT 1001.060 2793.450 1001.320 2793.595 ;
        RECT 986.800 2793.110 987.060 2793.430 ;
        RECT 1010.710 2792.915 1010.990 2793.285 ;
        RECT 1010.780 2789.350 1010.920 2792.915 ;
        RECT 1010.720 2789.030 1010.980 2789.350 ;
        RECT 1007.490 2788.155 1007.770 2788.525 ;
        RECT 1007.560 2787.990 1007.700 2788.155 ;
        RECT 1007.500 2787.670 1007.760 2787.990 ;
        RECT 979.900 2721.710 980.160 2722.030 ;
        RECT 1010.780 2717.610 1010.920 2789.030 ;
        RECT 1010.720 2717.290 1010.980 2717.610 ;
        RECT 948.160 2716.950 948.420 2717.270 ;
        RECT 948.220 2700.000 948.360 2716.950 ;
        RECT 968.860 2716.610 969.120 2716.930 ;
        RECT 958.740 2712.870 959.000 2713.190 ;
        RECT 958.800 2700.000 958.940 2712.870 ;
        RECT 968.920 2700.000 969.060 2716.610 ;
        RECT 989.560 2716.270 989.820 2716.590 ;
        RECT 979.440 2713.210 979.700 2713.530 ;
        RECT 979.500 2700.000 979.640 2713.210 ;
        RECT 989.620 2700.000 989.760 2716.270 ;
        RECT 1010.260 2715.930 1010.520 2716.250 ;
        RECT 1000.140 2713.550 1000.400 2713.870 ;
        RECT 1000.200 2700.000 1000.340 2713.550 ;
        RECT 1010.320 2700.000 1010.460 2715.930 ;
        RECT 1014.000 2715.230 1014.140 2794.275 ;
        RECT 1019.060 2791.050 1019.200 2794.275 ;
        RECT 1019.000 2790.730 1019.260 2791.050 ;
        RECT 1019.060 2788.330 1019.200 2790.730 ;
        RECT 1019.000 2788.010 1019.260 2788.330 ;
        RECT 1013.940 2714.910 1014.200 2715.230 ;
        RECT 1020.900 2714.970 1021.040 2794.275 ;
        RECT 1024.510 2792.915 1024.790 2793.285 ;
        RECT 1024.580 2788.330 1024.720 2792.915 ;
        RECT 1024.520 2788.010 1024.780 2788.330 ;
        RECT 1024.580 2717.950 1024.720 2788.010 ;
        RECT 1024.520 2717.630 1024.780 2717.950 ;
        RECT 1020.900 2714.830 1021.500 2714.970 ;
        RECT 1020.840 2713.890 1021.100 2714.210 ;
        RECT 1020.900 2700.000 1021.040 2713.890 ;
        RECT 1021.360 2713.530 1021.500 2714.830 ;
        RECT 1027.800 2713.870 1027.940 2794.275 ;
        RECT 1034.700 2791.390 1034.840 2794.275 ;
        RECT 1042.520 2792.750 1042.660 2794.275 ;
        RECT 1053.040 2794.130 1053.300 2794.450 ;
        RECT 1045.210 2792.915 1045.490 2793.285 ;
        RECT 1042.460 2792.430 1042.720 2792.750 ;
        RECT 1034.640 2791.070 1034.900 2791.390 ;
        RECT 1034.700 2788.670 1034.840 2791.070 ;
        RECT 1042.520 2789.010 1042.660 2792.430 ;
        RECT 1042.460 2788.690 1042.720 2789.010 ;
        RECT 1045.280 2788.670 1045.420 2792.915 ;
        RECT 1034.640 2788.350 1034.900 2788.670 ;
        RECT 1038.310 2788.155 1038.590 2788.525 ;
        RECT 1045.220 2788.350 1045.480 2788.670 ;
        RECT 1038.380 2787.990 1038.520 2788.155 ;
        RECT 1034.630 2787.475 1034.910 2787.845 ;
        RECT 1038.320 2787.670 1038.580 2787.990 ;
        RECT 1030.960 2715.590 1031.220 2715.910 ;
        RECT 1027.740 2713.550 1028.000 2713.870 ;
        RECT 1021.300 2713.210 1021.560 2713.530 ;
        RECT 1031.020 2700.000 1031.160 2715.590 ;
        RECT 1034.700 2714.210 1034.840 2787.475 ;
        RECT 1038.380 2718.290 1038.520 2787.670 ;
        RECT 1041.530 2787.475 1041.810 2787.845 ;
        RECT 1038.320 2717.970 1038.580 2718.290 ;
        RECT 1041.600 2717.950 1041.740 2787.475 ;
        RECT 1045.280 2718.630 1045.420 2788.350 ;
        RECT 1048.430 2787.475 1048.710 2787.845 ;
        RECT 1045.220 2718.310 1045.480 2718.630 ;
        RECT 1041.540 2717.630 1041.800 2717.950 ;
        RECT 1048.500 2717.610 1048.640 2787.475 ;
        RECT 1048.440 2717.290 1048.700 2717.610 ;
        RECT 1054.940 2716.250 1055.080 2799.715 ;
        RECT 1059.010 2794.275 1059.290 2794.645 ;
        RECT 1065.450 2794.275 1065.730 2794.645 ;
        RECT 1069.590 2794.275 1069.870 2794.645 ;
        RECT 1082.930 2794.275 1083.210 2794.645 ;
        RECT 1087.530 2794.275 1087.810 2794.645 ;
        RECT 1089.830 2794.275 1090.110 2794.645 ;
        RECT 1094.430 2794.275 1094.710 2794.645 ;
        RECT 1096.730 2794.275 1097.010 2794.645 ;
        RECT 1100.870 2794.275 1101.150 2794.645 ;
        RECT 1103.630 2794.275 1103.910 2794.645 ;
        RECT 1105.470 2794.275 1105.750 2794.645 ;
        RECT 1110.530 2794.275 1110.810 2794.645 ;
        RECT 1111.450 2794.275 1111.730 2794.645 ;
        RECT 1118.350 2794.275 1118.630 2794.645 ;
        RECT 1124.330 2794.275 1124.610 2794.645 ;
        RECT 1129.390 2794.275 1129.670 2794.645 ;
        RECT 1131.230 2794.275 1131.510 2794.645 ;
        RECT 1135.830 2794.275 1136.110 2794.645 ;
        RECT 1138.130 2794.275 1138.410 2794.645 ;
        RECT 1139.970 2794.275 1140.250 2794.645 ;
        RECT 1145.030 2794.275 1145.310 2794.645 ;
        RECT 1146.410 2794.275 1146.690 2794.645 ;
        RECT 1151.930 2794.275 1152.210 2794.645 ;
        RECT 1158.830 2794.275 1159.110 2794.645 ;
        RECT 1165.270 2794.275 1165.550 2794.645 ;
        RECT 1172.630 2794.275 1172.910 2794.645 ;
        RECT 1179.530 2794.275 1179.810 2794.645 ;
        RECT 1186.430 2794.275 1186.710 2794.645 ;
        RECT 1200.230 2794.275 1200.510 2794.645 ;
        RECT 1059.080 2792.410 1059.220 2794.275 ;
        RECT 1055.800 2792.090 1056.060 2792.410 ;
        RECT 1059.020 2792.090 1059.280 2792.410 ;
        RECT 1055.860 2789.350 1056.000 2792.090 ;
        RECT 1065.520 2791.730 1065.660 2794.275 ;
        RECT 1065.460 2791.410 1065.720 2791.730 ;
        RECT 1069.660 2791.050 1069.800 2794.275 ;
        RECT 1076.490 2793.595 1076.770 2793.965 ;
        RECT 1076.560 2791.390 1076.700 2793.595 ;
        RECT 1076.500 2791.070 1076.760 2791.390 ;
        RECT 1069.600 2790.730 1069.860 2791.050 ;
        RECT 1055.800 2789.030 1056.060 2789.350 ;
        RECT 1055.330 2788.155 1055.610 2788.525 ;
        RECT 1069.660 2788.330 1069.800 2790.730 ;
        RECT 1055.400 2717.270 1055.540 2788.155 ;
        RECT 1069.600 2788.010 1069.860 2788.330 ;
        RECT 1062.230 2787.475 1062.510 2787.845 ;
        RECT 1069.130 2787.475 1069.410 2787.845 ;
        RECT 1076.030 2787.475 1076.310 2787.845 ;
        RECT 1055.340 2716.950 1055.600 2717.270 ;
        RECT 1062.300 2716.930 1062.440 2787.475 ;
        RECT 1062.240 2716.610 1062.500 2716.930 ;
        RECT 1054.880 2715.930 1055.140 2716.250 ;
        RECT 1069.200 2715.910 1069.340 2787.475 ;
        RECT 1076.100 2716.590 1076.240 2787.475 ;
        RECT 1076.040 2716.270 1076.300 2716.590 ;
        RECT 1069.140 2715.590 1069.400 2715.910 ;
        RECT 1083.000 2715.570 1083.140 2794.275 ;
        RECT 1083.390 2793.595 1083.670 2793.965 ;
        RECT 1083.460 2793.430 1083.600 2793.595 ;
        RECT 1083.400 2793.110 1083.660 2793.430 ;
        RECT 1083.460 2787.990 1083.600 2793.110 ;
        RECT 1087.600 2792.750 1087.740 2794.275 ;
        RECT 1089.370 2793.595 1089.650 2793.965 ;
        RECT 1087.540 2792.430 1087.800 2792.750 ;
        RECT 1083.400 2787.670 1083.660 2787.990 ;
        RECT 1062.240 2715.250 1062.500 2715.570 ;
        RECT 1082.940 2715.250 1083.200 2715.570 ;
        RECT 1052.120 2714.570 1052.380 2714.890 ;
        RECT 1041.540 2714.230 1041.800 2714.550 ;
        RECT 1034.640 2713.890 1034.900 2714.210 ;
        RECT 1041.600 2700.000 1041.740 2714.230 ;
        RECT 1052.180 2700.000 1052.320 2714.570 ;
        RECT 1062.300 2700.000 1062.440 2715.250 ;
        RECT 1089.440 2715.230 1089.580 2793.595 ;
        RECT 1072.820 2714.910 1073.080 2715.230 ;
        RECT 1089.380 2714.910 1089.640 2715.230 ;
        RECT 1072.880 2700.000 1073.020 2714.910 ;
        RECT 1082.940 2713.210 1083.200 2713.530 ;
        RECT 1083.000 2700.000 1083.140 2713.210 ;
        RECT 1089.900 2712.850 1090.040 2794.275 ;
        RECT 1094.500 2793.770 1094.640 2794.275 ;
        RECT 1090.300 2793.450 1090.560 2793.770 ;
        RECT 1094.440 2793.450 1094.700 2793.770 ;
        RECT 1090.360 2788.670 1090.500 2793.450 ;
        RECT 1090.300 2788.350 1090.560 2788.670 ;
        RECT 1093.520 2713.550 1093.780 2713.870 ;
        RECT 1089.840 2712.530 1090.100 2712.850 ;
        RECT 1093.580 2700.000 1093.720 2713.550 ;
        RECT 1096.800 2712.510 1096.940 2794.275 ;
        RECT 1100.940 2792.070 1101.080 2794.275 ;
        RECT 1100.880 2791.750 1101.140 2792.070 ;
        RECT 1103.700 2714.890 1103.840 2794.275 ;
        RECT 1105.540 2792.410 1105.680 2794.275 ;
        RECT 1105.480 2792.090 1105.740 2792.410 ;
        RECT 1103.640 2714.570 1103.900 2714.890 ;
        RECT 1103.640 2713.890 1103.900 2714.210 ;
        RECT 1096.740 2712.190 1097.000 2712.510 ;
        RECT 1103.700 2700.000 1103.840 2713.890 ;
        RECT 1110.600 2713.190 1110.740 2794.275 ;
        RECT 1111.520 2791.730 1111.660 2794.275 ;
        RECT 1117.430 2792.235 1117.710 2792.605 ;
        RECT 1111.460 2791.410 1111.720 2791.730 ;
        RECT 1114.220 2717.630 1114.480 2717.950 ;
        RECT 1110.540 2712.870 1110.800 2713.190 ;
        RECT 1114.280 2700.000 1114.420 2717.630 ;
        RECT 1117.500 2714.210 1117.640 2792.235 ;
        RECT 1118.420 2791.050 1118.560 2794.275 ;
        RECT 1122.030 2793.595 1122.310 2793.965 ;
        RECT 1122.100 2793.090 1122.240 2793.595 ;
        RECT 1122.040 2792.770 1122.300 2793.090 ;
        RECT 1122.100 2791.390 1122.240 2792.770 ;
        RECT 1122.040 2791.070 1122.300 2791.390 ;
        RECT 1118.360 2790.730 1118.620 2791.050 ;
        RECT 1124.400 2726.530 1124.540 2794.275 ;
        RECT 1129.460 2793.430 1129.600 2794.275 ;
        RECT 1130.770 2793.595 1131.050 2793.965 ;
        RECT 1129.400 2793.110 1129.660 2793.430 ;
        RECT 1123.480 2726.390 1124.540 2726.530 ;
        RECT 1117.440 2713.890 1117.700 2714.210 ;
        RECT 1123.480 2713.870 1123.620 2726.390 ;
        RECT 1124.340 2717.290 1124.600 2717.610 ;
        RECT 1123.420 2713.550 1123.680 2713.870 ;
        RECT 1124.400 2700.000 1124.540 2717.290 ;
        RECT 1130.840 2714.550 1130.980 2793.595 ;
        RECT 1131.300 2714.890 1131.440 2794.275 ;
        RECT 1135.900 2792.750 1136.040 2794.275 ;
        RECT 1135.840 2792.430 1136.100 2792.750 ;
        RECT 1138.200 2718.290 1138.340 2794.275 ;
        RECT 1140.040 2793.770 1140.180 2794.275 ;
        RECT 1139.980 2793.450 1140.240 2793.770 ;
        RECT 1145.100 2718.630 1145.240 2794.275 ;
        RECT 1146.480 2792.070 1146.620 2794.275 ;
        RECT 1146.420 2791.750 1146.680 2792.070 ;
        RECT 1146.480 2791.390 1146.620 2791.750 ;
        RECT 1146.420 2791.070 1146.680 2791.390 ;
        RECT 1145.040 2718.310 1145.300 2718.630 ;
        RECT 1138.140 2717.970 1138.400 2718.290 ;
        RECT 1152.000 2717.610 1152.140 2794.275 ;
        RECT 1152.390 2792.235 1152.670 2792.605 ;
        RECT 1152.400 2792.090 1152.660 2792.235 ;
        RECT 1158.900 2717.950 1159.040 2794.275 ;
        RECT 1159.290 2791.555 1159.570 2791.925 ;
        RECT 1159.300 2791.410 1159.560 2791.555 ;
        RECT 1159.290 2790.875 1159.570 2791.245 ;
        RECT 1159.300 2790.730 1159.560 2790.875 ;
        RECT 1158.840 2717.630 1159.100 2717.950 ;
        RECT 1151.940 2717.290 1152.200 2717.610 ;
        RECT 1134.920 2716.950 1135.180 2717.270 ;
        RECT 1131.240 2714.570 1131.500 2714.890 ;
        RECT 1130.780 2714.230 1131.040 2714.550 ;
        RECT 1134.980 2700.000 1135.120 2716.950 ;
        RECT 1165.340 2716.930 1165.480 2794.275 ;
        RECT 1165.730 2793.595 1166.010 2793.965 ;
        RECT 1165.800 2717.270 1165.940 2793.595 ;
        RECT 1166.190 2792.915 1166.470 2793.285 ;
        RECT 1166.200 2792.770 1166.460 2792.915 ;
        RECT 1165.740 2716.950 1166.000 2717.270 ;
        RECT 1155.620 2716.610 1155.880 2716.930 ;
        RECT 1165.280 2716.610 1165.540 2716.930 ;
        RECT 1145.500 2715.930 1145.760 2716.250 ;
        RECT 1145.560 2700.000 1145.700 2715.930 ;
        RECT 1155.680 2700.000 1155.820 2716.610 ;
        RECT 1172.700 2716.250 1172.840 2794.275 ;
        RECT 1173.090 2793.595 1173.370 2793.965 ;
        RECT 1173.160 2793.430 1173.300 2793.595 ;
        RECT 1173.100 2793.110 1173.360 2793.430 ;
        RECT 1179.600 2716.590 1179.740 2794.275 ;
        RECT 1179.990 2793.595 1180.270 2793.965 ;
        RECT 1180.060 2792.750 1180.200 2793.595 ;
        RECT 1180.000 2792.430 1180.260 2792.750 ;
        RECT 1176.320 2716.270 1176.580 2716.590 ;
        RECT 1179.540 2716.270 1179.800 2716.590 ;
        RECT 1172.640 2715.930 1172.900 2716.250 ;
        RECT 1166.200 2715.590 1166.460 2715.910 ;
        RECT 1166.260 2700.000 1166.400 2715.590 ;
        RECT 1176.380 2700.000 1176.520 2716.270 ;
        RECT 1186.500 2715.910 1186.640 2794.275 ;
        RECT 1186.890 2793.595 1187.170 2793.965 ;
        RECT 1186.900 2793.450 1187.160 2793.595 ;
        RECT 1193.790 2791.555 1194.070 2791.925 ;
        RECT 1193.860 2791.390 1194.000 2791.555 ;
        RECT 1193.800 2791.070 1194.060 2791.390 ;
        RECT 1193.330 2790.195 1193.610 2790.565 ;
        RECT 1186.440 2715.590 1186.700 2715.910 ;
        RECT 1193.400 2715.570 1193.540 2790.195 ;
        RECT 1186.900 2715.250 1187.160 2715.570 ;
        RECT 1193.340 2715.250 1193.600 2715.570 ;
        RECT 1186.960 2700.000 1187.100 2715.250 ;
        RECT 1200.300 2715.230 1200.440 2794.275 ;
        RECT 1300.980 2718.310 1301.240 2718.630 ;
        RECT 1290.400 2717.970 1290.660 2718.290 ;
        RECT 1197.020 2714.910 1197.280 2715.230 ;
        RECT 1200.240 2714.910 1200.500 2715.230 ;
        RECT 1197.080 2700.000 1197.220 2714.910 ;
        RECT 1280.280 2714.570 1280.540 2714.890 ;
        RECT 1269.700 2714.230 1269.960 2714.550 ;
        RECT 1249.000 2713.890 1249.260 2714.210 ;
        RECT 1228.300 2713.210 1228.560 2713.530 ;
        RECT 1207.600 2712.530 1207.860 2712.850 ;
        RECT 1207.660 2700.000 1207.800 2712.530 ;
        RECT 1217.720 2712.190 1217.980 2712.510 ;
        RECT 1217.780 2700.000 1217.920 2712.190 ;
        RECT 1228.360 2700.000 1228.500 2713.210 ;
        RECT 1238.880 2712.870 1239.140 2713.190 ;
        RECT 1238.940 2700.000 1239.080 2712.870 ;
        RECT 1249.060 2700.000 1249.200 2713.890 ;
        RECT 1259.580 2713.550 1259.840 2713.870 ;
        RECT 1259.640 2700.000 1259.780 2713.550 ;
        RECT 1269.760 2700.000 1269.900 2714.230 ;
        RECT 1280.340 2700.000 1280.480 2714.570 ;
        RECT 1290.460 2700.000 1290.600 2717.970 ;
        RECT 1301.040 2700.000 1301.180 2718.310 ;
        RECT 1321.680 2717.630 1321.940 2717.950 ;
        RECT 1311.100 2717.290 1311.360 2717.610 ;
        RECT 1311.160 2700.000 1311.300 2717.290 ;
        RECT 1321.740 2700.000 1321.880 2717.630 ;
        RECT 1332.260 2716.950 1332.520 2717.270 ;
        RECT 1332.320 2700.000 1332.460 2716.950 ;
        RECT 1342.380 2716.610 1342.640 2716.930 ;
        RECT 1342.440 2700.000 1342.580 2716.610 ;
        RECT 1363.080 2716.270 1363.340 2716.590 ;
        RECT 1352.960 2715.930 1353.220 2716.250 ;
        RECT 1353.020 2700.000 1353.160 2715.930 ;
        RECT 1363.140 2700.000 1363.280 2716.270 ;
        RECT 1373.660 2715.590 1373.920 2715.910 ;
        RECT 1373.720 2700.000 1373.860 2715.590 ;
        RECT 1383.780 2715.250 1384.040 2715.570 ;
        RECT 1383.840 2700.000 1383.980 2715.250 ;
        RECT 1394.360 2714.910 1394.620 2715.230 ;
        RECT 1394.420 2700.000 1394.560 2714.910 ;
        RECT 792.680 2699.330 792.960 2700.000 ;
        RECT 786.760 2699.190 792.960 2699.330 ;
      LAYER met2 ;
        RECT 782.660 2695.720 792.400 2697.365 ;
      LAYER met2 ;
        RECT 792.680 2696.000 792.960 2699.190 ;
      LAYER met2 ;
        RECT 793.240 2695.720 802.520 2697.365 ;
      LAYER met2 ;
        RECT 802.800 2696.000 803.080 2700.000 ;
        RECT 811.600 2699.870 813.660 2700.000 ;
      LAYER met2 ;
        RECT 803.360 2695.720 813.100 2697.365 ;
      LAYER met2 ;
        RECT 813.380 2696.000 813.660 2699.870 ;
      LAYER met2 ;
        RECT 813.940 2695.720 823.220 2697.365 ;
      LAYER met2 ;
        RECT 823.500 2696.000 823.780 2700.000 ;
        RECT 832.760 2699.870 834.360 2700.000 ;
      LAYER met2 ;
        RECT 824.060 2695.720 833.800 2697.365 ;
      LAYER met2 ;
        RECT 834.080 2696.000 834.360 2699.870 ;
      LAYER met2 ;
        RECT 834.640 2695.720 843.920 2697.365 ;
      LAYER met2 ;
        RECT 844.200 2696.000 844.480 2700.000 ;
      LAYER met2 ;
        RECT 844.760 2695.720 854.500 2697.365 ;
      LAYER met2 ;
        RECT 854.780 2696.000 855.060 2700.000 ;
      LAYER met2 ;
        RECT 855.340 2695.720 865.080 2697.365 ;
      LAYER met2 ;
        RECT 865.360 2696.000 865.640 2700.000 ;
      LAYER met2 ;
        RECT 865.920 2695.720 875.200 2697.365 ;
      LAYER met2 ;
        RECT 875.480 2696.000 875.760 2700.000 ;
      LAYER met2 ;
        RECT 876.040 2695.720 885.780 2697.365 ;
      LAYER met2 ;
        RECT 886.060 2696.000 886.340 2700.000 ;
      LAYER met2 ;
        RECT 886.620 2695.720 895.900 2697.365 ;
      LAYER met2 ;
        RECT 896.180 2696.000 896.460 2700.000 ;
      LAYER met2 ;
        RECT 896.740 2695.720 906.480 2697.365 ;
      LAYER met2 ;
        RECT 906.760 2696.000 907.040 2700.000 ;
      LAYER met2 ;
        RECT 907.320 2695.720 916.600 2697.365 ;
      LAYER met2 ;
        RECT 916.880 2696.000 917.160 2700.000 ;
      LAYER met2 ;
        RECT 917.440 2695.720 927.180 2697.365 ;
      LAYER met2 ;
        RECT 927.460 2696.000 927.740 2700.000 ;
      LAYER met2 ;
        RECT 928.020 2695.720 937.300 2697.365 ;
      LAYER met2 ;
        RECT 937.580 2696.000 937.860 2700.000 ;
      LAYER met2 ;
        RECT 938.140 2695.720 947.880 2697.365 ;
      LAYER met2 ;
        RECT 948.160 2696.000 948.440 2700.000 ;
      LAYER met2 ;
        RECT 948.720 2695.720 958.460 2697.365 ;
      LAYER met2 ;
        RECT 958.740 2696.000 959.020 2700.000 ;
      LAYER met2 ;
        RECT 959.300 2695.720 968.580 2697.365 ;
      LAYER met2 ;
        RECT 968.860 2696.000 969.140 2700.000 ;
      LAYER met2 ;
        RECT 969.420 2695.720 979.160 2697.365 ;
      LAYER met2 ;
        RECT 979.440 2696.000 979.720 2700.000 ;
      LAYER met2 ;
        RECT 980.000 2695.720 989.280 2697.365 ;
      LAYER met2 ;
        RECT 989.560 2696.000 989.840 2700.000 ;
      LAYER met2 ;
        RECT 990.120 2695.720 999.860 2697.365 ;
      LAYER met2 ;
        RECT 1000.140 2696.000 1000.420 2700.000 ;
      LAYER met2 ;
        RECT 1000.700 2695.720 1009.980 2697.365 ;
      LAYER met2 ;
        RECT 1010.260 2696.000 1010.540 2700.000 ;
      LAYER met2 ;
        RECT 1010.820 2695.720 1020.560 2697.365 ;
      LAYER met2 ;
        RECT 1020.840 2696.000 1021.120 2700.000 ;
      LAYER met2 ;
        RECT 1021.400 2695.720 1030.680 2697.365 ;
      LAYER met2 ;
        RECT 1030.960 2696.000 1031.240 2700.000 ;
      LAYER met2 ;
        RECT 1031.520 2695.720 1041.260 2697.365 ;
      LAYER met2 ;
        RECT 1041.540 2696.000 1041.820 2700.000 ;
      LAYER met2 ;
        RECT 1042.100 2695.720 1051.840 2697.365 ;
      LAYER met2 ;
        RECT 1052.120 2696.000 1052.400 2700.000 ;
      LAYER met2 ;
        RECT 1052.680 2695.720 1061.960 2697.365 ;
      LAYER met2 ;
        RECT 1062.240 2696.000 1062.520 2700.000 ;
      LAYER met2 ;
        RECT 1062.800 2695.720 1072.540 2697.365 ;
      LAYER met2 ;
        RECT 1072.820 2696.000 1073.100 2700.000 ;
      LAYER met2 ;
        RECT 1073.380 2695.720 1082.660 2697.365 ;
      LAYER met2 ;
        RECT 1082.940 2696.000 1083.220 2700.000 ;
      LAYER met2 ;
        RECT 1083.500 2695.720 1093.240 2697.365 ;
      LAYER met2 ;
        RECT 1093.520 2696.000 1093.800 2700.000 ;
      LAYER met2 ;
        RECT 1094.080 2695.720 1103.360 2697.365 ;
      LAYER met2 ;
        RECT 1103.640 2696.000 1103.920 2700.000 ;
      LAYER met2 ;
        RECT 1104.200 2695.720 1113.940 2697.365 ;
      LAYER met2 ;
        RECT 1114.220 2696.000 1114.500 2700.000 ;
      LAYER met2 ;
        RECT 1114.780 2695.720 1124.060 2697.365 ;
      LAYER met2 ;
        RECT 1124.340 2696.000 1124.620 2700.000 ;
      LAYER met2 ;
        RECT 1124.900 2695.720 1134.640 2697.365 ;
      LAYER met2 ;
        RECT 1134.920 2696.000 1135.200 2700.000 ;
      LAYER met2 ;
        RECT 1135.480 2695.720 1145.220 2697.365 ;
      LAYER met2 ;
        RECT 1145.500 2696.000 1145.780 2700.000 ;
      LAYER met2 ;
        RECT 1146.060 2695.720 1155.340 2697.365 ;
      LAYER met2 ;
        RECT 1155.620 2696.000 1155.900 2700.000 ;
      LAYER met2 ;
        RECT 1156.180 2695.720 1165.920 2697.365 ;
      LAYER met2 ;
        RECT 1166.200 2696.000 1166.480 2700.000 ;
      LAYER met2 ;
        RECT 1166.760 2695.720 1176.040 2697.365 ;
      LAYER met2 ;
        RECT 1176.320 2696.000 1176.600 2700.000 ;
      LAYER met2 ;
        RECT 1176.880 2695.720 1186.620 2697.365 ;
      LAYER met2 ;
        RECT 1186.900 2696.000 1187.180 2700.000 ;
      LAYER met2 ;
        RECT 1187.460 2695.720 1196.740 2697.365 ;
      LAYER met2 ;
        RECT 1197.020 2696.000 1197.300 2700.000 ;
      LAYER met2 ;
        RECT 1197.580 2695.720 1207.320 2697.365 ;
      LAYER met2 ;
        RECT 1207.600 2696.000 1207.880 2700.000 ;
      LAYER met2 ;
        RECT 1208.160 2695.720 1217.440 2697.365 ;
      LAYER met2 ;
        RECT 1217.720 2696.000 1218.000 2700.000 ;
      LAYER met2 ;
        RECT 1218.280 2695.720 1228.020 2697.365 ;
      LAYER met2 ;
        RECT 1228.300 2696.000 1228.580 2700.000 ;
      LAYER met2 ;
        RECT 1228.860 2695.720 1238.600 2697.365 ;
      LAYER met2 ;
        RECT 1238.880 2696.000 1239.160 2700.000 ;
      LAYER met2 ;
        RECT 1239.440 2695.720 1248.720 2697.365 ;
      LAYER met2 ;
        RECT 1249.000 2696.000 1249.280 2700.000 ;
      LAYER met2 ;
        RECT 1249.560 2695.720 1259.300 2697.365 ;
      LAYER met2 ;
        RECT 1259.580 2696.000 1259.860 2700.000 ;
      LAYER met2 ;
        RECT 1260.140 2695.720 1269.420 2697.365 ;
      LAYER met2 ;
        RECT 1269.700 2696.000 1269.980 2700.000 ;
      LAYER met2 ;
        RECT 1270.260 2695.720 1280.000 2697.365 ;
      LAYER met2 ;
        RECT 1280.280 2696.000 1280.560 2700.000 ;
      LAYER met2 ;
        RECT 1280.840 2695.720 1290.120 2697.365 ;
      LAYER met2 ;
        RECT 1290.400 2696.000 1290.680 2700.000 ;
      LAYER met2 ;
        RECT 1290.960 2695.720 1300.700 2697.365 ;
      LAYER met2 ;
        RECT 1300.980 2696.000 1301.260 2700.000 ;
      LAYER met2 ;
        RECT 1301.540 2695.720 1310.820 2697.365 ;
      LAYER met2 ;
        RECT 1311.100 2696.000 1311.380 2700.000 ;
      LAYER met2 ;
        RECT 1311.660 2695.720 1321.400 2697.365 ;
      LAYER met2 ;
        RECT 1321.680 2696.000 1321.960 2700.000 ;
      LAYER met2 ;
        RECT 1322.240 2695.720 1331.980 2697.365 ;
      LAYER met2 ;
        RECT 1332.260 2696.000 1332.540 2700.000 ;
      LAYER met2 ;
        RECT 1332.820 2695.720 1342.100 2697.365 ;
      LAYER met2 ;
        RECT 1342.380 2696.000 1342.660 2700.000 ;
      LAYER met2 ;
        RECT 1342.940 2695.720 1352.680 2697.365 ;
      LAYER met2 ;
        RECT 1352.960 2696.000 1353.240 2700.000 ;
      LAYER met2 ;
        RECT 1353.520 2695.720 1362.800 2697.365 ;
      LAYER met2 ;
        RECT 1363.080 2696.000 1363.360 2700.000 ;
      LAYER met2 ;
        RECT 1363.640 2695.720 1373.380 2697.365 ;
      LAYER met2 ;
        RECT 1373.660 2696.000 1373.940 2700.000 ;
      LAYER met2 ;
        RECT 1374.220 2695.720 1383.500 2697.365 ;
      LAYER met2 ;
        RECT 1383.780 2696.000 1384.060 2700.000 ;
      LAYER met2 ;
        RECT 1384.340 2695.720 1394.080 2697.365 ;
      LAYER met2 ;
        RECT 1394.360 2696.000 1394.640 2700.000 ;
      LAYER met2 ;
        RECT 1394.920 2695.720 1397.390 2697.365 ;
        RECT 300.030 1604.280 1397.390 2695.720 ;
        RECT 300.030 1602.195 302.040 1604.280 ;
        RECT 302.880 1602.195 306.640 1604.280 ;
        RECT 307.480 1602.195 311.700 1604.280 ;
        RECT 312.540 1602.195 316.300 1604.280 ;
        RECT 317.140 1602.195 321.360 1604.280 ;
        RECT 322.200 1602.195 325.960 1604.280 ;
        RECT 326.800 1602.195 331.020 1604.280 ;
        RECT 331.860 1602.195 335.620 1604.280 ;
        RECT 336.460 1602.195 340.680 1604.280 ;
        RECT 341.520 1602.195 345.280 1604.280 ;
        RECT 346.120 1602.195 350.340 1604.280 ;
        RECT 351.180 1602.195 354.940 1604.280 ;
        RECT 355.780 1602.195 360.000 1604.280 ;
        RECT 360.840 1602.195 364.600 1604.280 ;
        RECT 365.440 1602.195 369.660 1604.280 ;
        RECT 370.500 1602.195 374.260 1604.280 ;
        RECT 375.100 1602.195 379.320 1604.280 ;
        RECT 380.160 1602.195 384.380 1604.280 ;
        RECT 385.220 1602.195 388.980 1604.280 ;
        RECT 389.820 1602.195 394.040 1604.280 ;
        RECT 394.880 1602.195 398.640 1604.280 ;
        RECT 399.480 1602.195 403.700 1604.280 ;
        RECT 404.540 1602.195 408.300 1604.280 ;
        RECT 409.140 1602.195 413.360 1604.280 ;
        RECT 414.200 1602.195 417.960 1604.280 ;
        RECT 418.800 1602.195 423.020 1604.280 ;
        RECT 423.860 1602.195 427.620 1604.280 ;
        RECT 428.460 1602.195 432.680 1604.280 ;
        RECT 433.520 1602.195 437.280 1604.280 ;
        RECT 438.120 1602.195 442.340 1604.280 ;
        RECT 443.180 1602.195 446.940 1604.280 ;
        RECT 447.780 1602.195 452.000 1604.280 ;
        RECT 452.840 1602.195 457.060 1604.280 ;
        RECT 457.900 1602.195 461.660 1604.280 ;
        RECT 462.500 1602.195 466.720 1604.280 ;
        RECT 467.560 1602.195 471.320 1604.280 ;
        RECT 472.160 1602.195 476.380 1604.280 ;
        RECT 477.220 1602.195 480.980 1604.280 ;
        RECT 481.820 1602.195 486.040 1604.280 ;
        RECT 486.880 1602.195 490.640 1604.280 ;
        RECT 491.480 1602.195 495.700 1604.280 ;
        RECT 496.540 1602.195 500.300 1604.280 ;
        RECT 501.140 1602.195 505.360 1604.280 ;
        RECT 506.200 1602.195 509.960 1604.280 ;
        RECT 510.800 1602.195 515.020 1604.280 ;
        RECT 515.860 1602.195 519.620 1604.280 ;
        RECT 520.460 1602.195 524.680 1604.280 ;
        RECT 525.520 1602.195 529.740 1604.280 ;
        RECT 530.580 1602.195 534.340 1604.280 ;
        RECT 535.180 1602.195 539.400 1604.280 ;
        RECT 540.240 1602.195 544.000 1604.280 ;
        RECT 544.840 1602.195 549.060 1604.280 ;
        RECT 549.900 1602.195 553.660 1604.280 ;
        RECT 554.500 1602.195 558.720 1604.280 ;
        RECT 559.560 1602.195 563.320 1604.280 ;
        RECT 564.160 1602.195 568.380 1604.280 ;
        RECT 569.220 1602.195 572.980 1604.280 ;
        RECT 573.820 1602.195 578.040 1604.280 ;
        RECT 578.880 1602.195 582.640 1604.280 ;
        RECT 583.480 1602.195 587.700 1604.280 ;
        RECT 588.540 1602.195 592.300 1604.280 ;
        RECT 593.140 1602.195 597.360 1604.280 ;
        RECT 598.200 1602.195 602.420 1604.280 ;
        RECT 603.260 1602.195 607.020 1604.280 ;
        RECT 607.860 1602.195 612.080 1604.280 ;
        RECT 612.920 1602.195 616.680 1604.280 ;
        RECT 617.520 1602.195 621.740 1604.280 ;
        RECT 622.580 1602.195 626.340 1604.280 ;
        RECT 627.180 1602.195 631.400 1604.280 ;
        RECT 632.240 1602.195 636.000 1604.280 ;
        RECT 636.840 1602.195 641.060 1604.280 ;
        RECT 641.900 1602.195 645.660 1604.280 ;
        RECT 646.500 1602.195 650.720 1604.280 ;
        RECT 651.560 1602.195 655.320 1604.280 ;
        RECT 656.160 1602.195 660.380 1604.280 ;
        RECT 661.220 1602.195 664.980 1604.280 ;
        RECT 665.820 1602.195 670.040 1604.280 ;
        RECT 670.880 1602.195 675.100 1604.280 ;
        RECT 675.940 1602.195 679.700 1604.280 ;
        RECT 680.540 1602.195 684.760 1604.280 ;
        RECT 685.600 1602.195 689.360 1604.280 ;
        RECT 690.200 1602.195 694.420 1604.280 ;
        RECT 695.260 1602.195 699.020 1604.280 ;
        RECT 699.860 1602.195 704.080 1604.280 ;
        RECT 704.920 1602.195 708.680 1604.280 ;
        RECT 709.520 1602.195 713.740 1604.280 ;
        RECT 714.580 1602.195 718.340 1604.280 ;
        RECT 719.180 1602.195 723.400 1604.280 ;
        RECT 724.240 1602.195 728.000 1604.280 ;
        RECT 728.840 1602.195 733.060 1604.280 ;
        RECT 733.900 1602.195 737.660 1604.280 ;
        RECT 738.500 1602.195 742.720 1604.280 ;
        RECT 743.560 1602.195 747.780 1604.280 ;
        RECT 748.620 1602.195 752.380 1604.280 ;
        RECT 753.220 1602.195 757.440 1604.280 ;
        RECT 758.280 1602.195 762.040 1604.280 ;
        RECT 762.880 1602.195 767.100 1604.280 ;
        RECT 767.940 1602.195 771.700 1604.280 ;
        RECT 772.540 1602.195 776.760 1604.280 ;
        RECT 777.600 1602.195 781.360 1604.280 ;
        RECT 782.200 1602.195 786.420 1604.280 ;
        RECT 787.260 1602.195 791.020 1604.280 ;
        RECT 791.860 1602.195 796.080 1604.280 ;
        RECT 796.920 1602.195 800.680 1604.280 ;
        RECT 801.520 1602.195 805.740 1604.280 ;
        RECT 806.580 1602.195 810.340 1604.280 ;
        RECT 811.180 1602.195 815.400 1604.280 ;
        RECT 816.240 1602.195 820.460 1604.280 ;
        RECT 821.300 1602.195 825.060 1604.280 ;
        RECT 825.900 1602.195 830.120 1604.280 ;
        RECT 830.960 1602.195 834.720 1604.280 ;
        RECT 835.560 1602.195 839.780 1604.280 ;
        RECT 840.620 1602.195 844.380 1604.280 ;
        RECT 845.220 1602.195 849.440 1604.280 ;
      LAYER met2 ;
        RECT 849.720 1600.000 850.000 1604.000 ;
      LAYER met2 ;
        RECT 850.280 1602.195 854.040 1604.280 ;
      LAYER met2 ;
        RECT 854.320 1600.000 854.600 1604.000 ;
      LAYER met2 ;
        RECT 854.880 1602.195 859.100 1604.280 ;
      LAYER met2 ;
        RECT 859.380 1600.000 859.660 1604.000 ;
      LAYER met2 ;
        RECT 859.940 1602.195 863.700 1604.280 ;
      LAYER met2 ;
        RECT 863.980 1600.000 864.260 1604.000 ;
      LAYER met2 ;
        RECT 864.540 1602.195 868.760 1604.280 ;
      LAYER met2 ;
        RECT 869.040 1600.000 869.320 1604.000 ;
      LAYER met2 ;
        RECT 869.600 1602.195 873.360 1604.280 ;
      LAYER met2 ;
        RECT 873.640 1600.000 873.920 1604.000 ;
      LAYER met2 ;
        RECT 874.200 1602.195 878.420 1604.280 ;
      LAYER met2 ;
        RECT 878.700 1600.000 878.980 1604.000 ;
      LAYER met2 ;
        RECT 879.260 1602.195 883.020 1604.280 ;
      LAYER met2 ;
        RECT 883.300 1600.000 883.580 1604.000 ;
      LAYER met2 ;
        RECT 883.860 1602.195 888.080 1604.280 ;
      LAYER met2 ;
        RECT 888.360 1600.000 888.640 1604.000 ;
      LAYER met2 ;
        RECT 888.920 1602.195 893.140 1604.280 ;
      LAYER met2 ;
        RECT 893.420 1600.000 893.700 1604.000 ;
      LAYER met2 ;
        RECT 893.980 1602.195 897.740 1604.280 ;
      LAYER met2 ;
        RECT 898.020 1600.000 898.300 1604.000 ;
      LAYER met2 ;
        RECT 898.580 1602.195 902.800 1604.280 ;
      LAYER met2 ;
        RECT 903.080 1600.000 903.360 1604.000 ;
      LAYER met2 ;
        RECT 903.640 1602.195 907.400 1604.280 ;
      LAYER met2 ;
        RECT 907.680 1600.000 907.960 1604.000 ;
      LAYER met2 ;
        RECT 908.240 1602.195 912.460 1604.280 ;
      LAYER met2 ;
        RECT 912.740 1600.000 913.020 1604.000 ;
      LAYER met2 ;
        RECT 913.300 1602.195 917.060 1604.280 ;
      LAYER met2 ;
        RECT 917.340 1600.000 917.620 1604.000 ;
      LAYER met2 ;
        RECT 917.900 1602.195 922.120 1604.280 ;
      LAYER met2 ;
        RECT 922.400 1600.000 922.680 1604.000 ;
      LAYER met2 ;
        RECT 922.960 1602.195 926.720 1604.280 ;
      LAYER met2 ;
        RECT 927.000 1600.000 927.280 1604.000 ;
      LAYER met2 ;
        RECT 927.560 1602.195 931.780 1604.280 ;
      LAYER met2 ;
        RECT 932.060 1600.000 932.340 1604.000 ;
      LAYER met2 ;
        RECT 932.620 1602.195 936.380 1604.280 ;
      LAYER met2 ;
        RECT 936.660 1600.000 936.940 1604.000 ;
      LAYER met2 ;
        RECT 937.220 1602.195 941.440 1604.280 ;
      LAYER met2 ;
        RECT 941.720 1600.000 942.000 1604.000 ;
      LAYER met2 ;
        RECT 942.280 1602.195 946.040 1604.280 ;
      LAYER met2 ;
        RECT 946.320 1600.000 946.600 1604.000 ;
      LAYER met2 ;
        RECT 946.880 1602.195 951.100 1604.280 ;
      LAYER met2 ;
        RECT 951.380 1600.000 951.660 1604.000 ;
      LAYER met2 ;
        RECT 951.940 1602.195 955.700 1604.280 ;
      LAYER met2 ;
        RECT 955.980 1600.000 956.260 1604.000 ;
      LAYER met2 ;
        RECT 956.540 1602.195 960.760 1604.280 ;
      LAYER met2 ;
        RECT 961.040 1600.000 961.320 1604.000 ;
      LAYER met2 ;
        RECT 961.600 1602.195 965.820 1604.280 ;
      LAYER met2 ;
        RECT 966.100 1600.000 966.380 1604.000 ;
      LAYER met2 ;
        RECT 966.660 1602.195 970.420 1604.280 ;
      LAYER met2 ;
        RECT 970.700 1600.000 970.980 1604.000 ;
      LAYER met2 ;
        RECT 971.260 1602.195 975.480 1604.280 ;
      LAYER met2 ;
        RECT 975.760 1600.000 976.040 1604.000 ;
      LAYER met2 ;
        RECT 976.320 1602.195 980.080 1604.280 ;
      LAYER met2 ;
        RECT 980.360 1600.000 980.640 1604.000 ;
      LAYER met2 ;
        RECT 980.920 1602.195 985.140 1604.280 ;
      LAYER met2 ;
        RECT 985.420 1600.000 985.700 1604.000 ;
      LAYER met2 ;
        RECT 985.980 1602.195 989.740 1604.280 ;
      LAYER met2 ;
        RECT 990.020 1600.000 990.300 1604.000 ;
      LAYER met2 ;
        RECT 990.580 1602.195 994.800 1604.280 ;
      LAYER met2 ;
        RECT 995.080 1600.000 995.360 1604.000 ;
      LAYER met2 ;
        RECT 995.640 1602.195 999.400 1604.280 ;
      LAYER met2 ;
        RECT 999.680 1600.000 999.960 1604.000 ;
      LAYER met2 ;
        RECT 1000.240 1602.195 1004.460 1604.280 ;
      LAYER met2 ;
        RECT 1004.740 1600.000 1005.020 1604.000 ;
      LAYER met2 ;
        RECT 1005.300 1602.195 1009.060 1604.280 ;
      LAYER met2 ;
        RECT 1009.340 1600.000 1009.620 1604.000 ;
      LAYER met2 ;
        RECT 1009.900 1602.195 1014.120 1604.280 ;
      LAYER met2 ;
        RECT 1014.400 1600.000 1014.680 1604.000 ;
      LAYER met2 ;
        RECT 1014.960 1602.195 1018.720 1604.280 ;
      LAYER met2 ;
        RECT 1019.000 1600.000 1019.280 1604.000 ;
      LAYER met2 ;
        RECT 1019.560 1602.195 1023.780 1604.280 ;
      LAYER met2 ;
        RECT 1024.060 1600.000 1024.340 1604.000 ;
      LAYER met2 ;
        RECT 1024.620 1602.195 1028.380 1604.280 ;
      LAYER met2 ;
        RECT 1028.660 1600.000 1028.940 1604.000 ;
      LAYER met2 ;
        RECT 1029.220 1602.195 1033.440 1604.280 ;
      LAYER met2 ;
        RECT 1033.720 1600.000 1034.000 1604.000 ;
      LAYER met2 ;
        RECT 1034.280 1602.195 1038.500 1604.280 ;
      LAYER met2 ;
        RECT 1038.780 1600.000 1039.060 1604.000 ;
      LAYER met2 ;
        RECT 1039.340 1602.195 1043.100 1604.280 ;
      LAYER met2 ;
        RECT 1043.380 1600.000 1043.660 1604.000 ;
      LAYER met2 ;
        RECT 1043.940 1602.195 1048.160 1604.280 ;
      LAYER met2 ;
        RECT 1048.440 1600.000 1048.720 1604.000 ;
      LAYER met2 ;
        RECT 1049.000 1602.195 1052.760 1604.280 ;
      LAYER met2 ;
        RECT 1053.040 1600.000 1053.320 1604.000 ;
      LAYER met2 ;
        RECT 1053.600 1602.195 1057.820 1604.280 ;
      LAYER met2 ;
        RECT 1058.100 1600.000 1058.380 1604.000 ;
      LAYER met2 ;
        RECT 1058.660 1602.195 1062.420 1604.280 ;
      LAYER met2 ;
        RECT 1062.700 1600.000 1062.980 1604.000 ;
      LAYER met2 ;
        RECT 1063.260 1602.195 1067.480 1604.280 ;
      LAYER met2 ;
        RECT 1067.760 1600.000 1068.040 1604.000 ;
      LAYER met2 ;
        RECT 1068.320 1602.195 1072.080 1604.280 ;
      LAYER met2 ;
        RECT 1072.360 1600.000 1072.640 1604.000 ;
      LAYER met2 ;
        RECT 1072.920 1602.195 1077.140 1604.280 ;
      LAYER met2 ;
        RECT 1077.420 1600.000 1077.700 1604.000 ;
      LAYER met2 ;
        RECT 1077.980 1602.195 1081.740 1604.280 ;
      LAYER met2 ;
        RECT 1082.020 1600.000 1082.300 1604.000 ;
      LAYER met2 ;
        RECT 1082.580 1602.195 1086.800 1604.280 ;
      LAYER met2 ;
        RECT 1087.080 1600.000 1087.360 1604.000 ;
      LAYER met2 ;
        RECT 1087.640 1602.195 1091.400 1604.280 ;
      LAYER met2 ;
        RECT 1091.680 1600.000 1091.960 1604.000 ;
      LAYER met2 ;
        RECT 1092.240 1602.195 1096.460 1604.280 ;
      LAYER met2 ;
        RECT 1096.740 1600.000 1097.020 1604.000 ;
      LAYER met2 ;
        RECT 1097.300 1602.195 1101.060 1604.280 ;
      LAYER met2 ;
        RECT 1101.340 1600.000 1101.620 1604.000 ;
      LAYER met2 ;
        RECT 1101.900 1602.195 1106.120 1604.280 ;
      LAYER met2 ;
        RECT 1106.400 1600.000 1106.680 1604.000 ;
      LAYER met2 ;
        RECT 1106.960 1602.195 1111.180 1604.280 ;
      LAYER met2 ;
        RECT 1111.460 1600.000 1111.740 1604.000 ;
      LAYER met2 ;
        RECT 1112.020 1602.195 1115.780 1604.280 ;
      LAYER met2 ;
        RECT 1116.060 1600.000 1116.340 1604.000 ;
      LAYER met2 ;
        RECT 1116.620 1602.195 1120.840 1604.280 ;
      LAYER met2 ;
        RECT 1121.120 1600.000 1121.400 1604.000 ;
      LAYER met2 ;
        RECT 1121.680 1602.195 1125.440 1604.280 ;
      LAYER met2 ;
        RECT 1125.720 1600.000 1126.000 1604.000 ;
      LAYER met2 ;
        RECT 1126.280 1602.195 1130.500 1604.280 ;
      LAYER met2 ;
        RECT 1130.780 1600.000 1131.060 1604.000 ;
      LAYER met2 ;
        RECT 1131.340 1602.195 1135.100 1604.280 ;
      LAYER met2 ;
        RECT 1135.380 1600.000 1135.660 1604.000 ;
      LAYER met2 ;
        RECT 1135.940 1602.195 1140.160 1604.280 ;
      LAYER met2 ;
        RECT 1140.440 1600.000 1140.720 1604.000 ;
      LAYER met2 ;
        RECT 1141.000 1602.195 1144.760 1604.280 ;
      LAYER met2 ;
        RECT 1145.040 1600.000 1145.320 1604.000 ;
      LAYER met2 ;
        RECT 1145.600 1602.195 1149.820 1604.280 ;
      LAYER met2 ;
        RECT 1150.100 1600.000 1150.380 1604.000 ;
      LAYER met2 ;
        RECT 1150.660 1602.195 1154.420 1604.280 ;
      LAYER met2 ;
        RECT 1154.700 1600.000 1154.980 1604.000 ;
      LAYER met2 ;
        RECT 1155.260 1602.195 1159.480 1604.280 ;
      LAYER met2 ;
        RECT 1159.760 1600.000 1160.040 1604.000 ;
      LAYER met2 ;
        RECT 1160.320 1602.195 1164.080 1604.280 ;
      LAYER met2 ;
        RECT 1164.360 1600.000 1164.640 1604.000 ;
      LAYER met2 ;
        RECT 1164.920 1602.195 1169.140 1604.280 ;
      LAYER met2 ;
        RECT 1169.420 1600.000 1169.700 1604.000 ;
      LAYER met2 ;
        RECT 1169.980 1602.195 1173.740 1604.280 ;
      LAYER met2 ;
        RECT 1174.020 1600.000 1174.300 1604.000 ;
      LAYER met2 ;
        RECT 1174.580 1602.195 1178.800 1604.280 ;
      LAYER met2 ;
        RECT 1179.080 1600.000 1179.360 1604.000 ;
      LAYER met2 ;
        RECT 1179.640 1602.195 1183.860 1604.280 ;
      LAYER met2 ;
        RECT 1184.140 1600.000 1184.420 1604.000 ;
      LAYER met2 ;
        RECT 1184.700 1602.195 1188.460 1604.280 ;
      LAYER met2 ;
        RECT 1188.740 1600.000 1189.020 1604.000 ;
      LAYER met2 ;
        RECT 1189.300 1602.195 1193.520 1604.280 ;
      LAYER met2 ;
        RECT 1193.800 1600.000 1194.080 1604.000 ;
      LAYER met2 ;
        RECT 1194.360 1602.195 1198.120 1604.280 ;
      LAYER met2 ;
        RECT 1198.400 1600.000 1198.680 1604.000 ;
      LAYER met2 ;
        RECT 1198.960 1602.195 1203.180 1604.280 ;
      LAYER met2 ;
        RECT 1203.460 1600.000 1203.740 1604.000 ;
      LAYER met2 ;
        RECT 1204.020 1602.195 1207.780 1604.280 ;
      LAYER met2 ;
        RECT 1208.060 1600.000 1208.340 1604.000 ;
      LAYER met2 ;
        RECT 1208.620 1602.195 1212.840 1604.280 ;
      LAYER met2 ;
        RECT 1213.120 1600.000 1213.400 1604.000 ;
      LAYER met2 ;
        RECT 1213.680 1602.195 1217.440 1604.280 ;
      LAYER met2 ;
        RECT 1217.720 1600.000 1218.000 1604.000 ;
      LAYER met2 ;
        RECT 1218.280 1602.195 1222.500 1604.280 ;
      LAYER met2 ;
        RECT 1222.780 1600.000 1223.060 1604.000 ;
      LAYER met2 ;
        RECT 1223.340 1602.195 1227.100 1604.280 ;
      LAYER met2 ;
        RECT 1227.380 1600.000 1227.660 1604.000 ;
      LAYER met2 ;
        RECT 1227.940 1602.195 1232.160 1604.280 ;
      LAYER met2 ;
        RECT 1232.440 1600.000 1232.720 1604.000 ;
      LAYER met2 ;
        RECT 1233.000 1602.195 1236.760 1604.280 ;
      LAYER met2 ;
        RECT 1237.040 1600.000 1237.320 1604.000 ;
      LAYER met2 ;
        RECT 1237.600 1602.195 1241.820 1604.280 ;
      LAYER met2 ;
        RECT 1242.100 1600.000 1242.380 1604.000 ;
      LAYER met2 ;
        RECT 1242.660 1602.195 1246.420 1604.280 ;
      LAYER met2 ;
        RECT 1246.700 1600.000 1246.980 1604.000 ;
      LAYER met2 ;
        RECT 1247.260 1602.195 1251.480 1604.280 ;
      LAYER met2 ;
        RECT 1251.760 1600.000 1252.040 1604.000 ;
      LAYER met2 ;
        RECT 1252.320 1602.195 1256.540 1604.280 ;
      LAYER met2 ;
        RECT 1256.820 1600.000 1257.100 1604.000 ;
      LAYER met2 ;
        RECT 1257.380 1602.195 1261.140 1604.280 ;
      LAYER met2 ;
        RECT 1261.420 1600.000 1261.700 1604.000 ;
      LAYER met2 ;
        RECT 1261.980 1602.195 1266.200 1604.280 ;
      LAYER met2 ;
        RECT 1266.480 1600.000 1266.760 1604.000 ;
      LAYER met2 ;
        RECT 1267.040 1602.195 1270.800 1604.280 ;
      LAYER met2 ;
        RECT 1271.080 1600.000 1271.360 1604.000 ;
      LAYER met2 ;
        RECT 1271.640 1602.195 1275.860 1604.280 ;
      LAYER met2 ;
        RECT 1276.140 1600.000 1276.420 1604.000 ;
      LAYER met2 ;
        RECT 1276.700 1602.195 1280.460 1604.280 ;
      LAYER met2 ;
        RECT 1280.740 1600.000 1281.020 1604.000 ;
      LAYER met2 ;
        RECT 1281.300 1602.195 1285.520 1604.280 ;
      LAYER met2 ;
        RECT 1285.800 1600.000 1286.080 1604.000 ;
      LAYER met2 ;
        RECT 1286.360 1602.195 1290.120 1604.280 ;
      LAYER met2 ;
        RECT 1290.400 1600.000 1290.680 1604.000 ;
      LAYER met2 ;
        RECT 1290.960 1602.195 1295.180 1604.280 ;
      LAYER met2 ;
        RECT 1295.460 1600.000 1295.740 1604.000 ;
      LAYER met2 ;
        RECT 1296.020 1602.195 1299.780 1604.280 ;
      LAYER met2 ;
        RECT 1300.060 1600.000 1300.340 1604.000 ;
      LAYER met2 ;
        RECT 1300.620 1602.195 1304.840 1604.280 ;
      LAYER met2 ;
        RECT 1305.120 1600.000 1305.400 1604.000 ;
      LAYER met2 ;
        RECT 1305.680 1602.195 1309.440 1604.280 ;
      LAYER met2 ;
        RECT 1309.720 1600.000 1310.000 1604.000 ;
      LAYER met2 ;
        RECT 1310.280 1602.195 1314.500 1604.280 ;
      LAYER met2 ;
        RECT 1314.780 1600.000 1315.060 1604.000 ;
      LAYER met2 ;
        RECT 1315.340 1602.195 1319.100 1604.280 ;
      LAYER met2 ;
        RECT 1319.380 1600.000 1319.660 1604.000 ;
      LAYER met2 ;
        RECT 1319.940 1602.195 1324.160 1604.280 ;
      LAYER met2 ;
        RECT 1324.440 1600.000 1324.720 1604.000 ;
      LAYER met2 ;
        RECT 1325.000 1602.195 1329.220 1604.280 ;
      LAYER met2 ;
        RECT 1329.500 1600.000 1329.780 1604.000 ;
      LAYER met2 ;
        RECT 1330.060 1602.195 1333.820 1604.280 ;
      LAYER met2 ;
        RECT 1334.100 1600.000 1334.380 1604.000 ;
      LAYER met2 ;
        RECT 1334.660 1602.195 1338.880 1604.280 ;
      LAYER met2 ;
        RECT 1339.160 1600.000 1339.440 1604.000 ;
      LAYER met2 ;
        RECT 1339.720 1602.195 1343.480 1604.280 ;
      LAYER met2 ;
        RECT 1343.760 1600.000 1344.040 1604.000 ;
      LAYER met2 ;
        RECT 1344.320 1602.195 1348.540 1604.280 ;
      LAYER met2 ;
        RECT 1348.820 1600.000 1349.100 1604.000 ;
      LAYER met2 ;
        RECT 1349.380 1602.195 1353.140 1604.280 ;
      LAYER met2 ;
        RECT 1353.420 1600.000 1353.700 1604.000 ;
      LAYER met2 ;
        RECT 1353.980 1602.195 1358.200 1604.280 ;
      LAYER met2 ;
        RECT 1358.480 1600.000 1358.760 1604.000 ;
      LAYER met2 ;
        RECT 1359.040 1602.195 1362.800 1604.280 ;
      LAYER met2 ;
        RECT 1363.080 1600.000 1363.360 1604.000 ;
      LAYER met2 ;
        RECT 1363.640 1602.195 1367.860 1604.280 ;
      LAYER met2 ;
        RECT 1368.140 1600.000 1368.420 1604.000 ;
      LAYER met2 ;
        RECT 1368.700 1602.195 1372.460 1604.280 ;
      LAYER met2 ;
        RECT 1372.740 1600.000 1373.020 1604.000 ;
      LAYER met2 ;
        RECT 1373.300 1602.195 1377.520 1604.280 ;
      LAYER met2 ;
        RECT 1377.800 1600.000 1378.080 1604.000 ;
      LAYER met2 ;
        RECT 1378.360 1602.195 1382.120 1604.280 ;
      LAYER met2 ;
        RECT 1382.400 1600.000 1382.680 1604.000 ;
      LAYER met2 ;
        RECT 1382.960 1602.195 1387.180 1604.280 ;
      LAYER met2 ;
        RECT 1387.460 1600.000 1387.740 1604.000 ;
      LAYER met2 ;
        RECT 1388.020 1602.195 1391.780 1604.280 ;
      LAYER met2 ;
        RECT 1392.060 1600.000 1392.340 1604.000 ;
      LAYER met2 ;
        RECT 1392.620 1602.195 1396.840 1604.280 ;
      LAYER met2 ;
        RECT 1397.120 1600.000 1397.400 1604.000 ;
        RECT 1397.640 1603.965 1397.780 2901.230 ;
        RECT 1407.760 1607.365 1407.900 3250.750 ;
        RECT 1536.950 3230.155 1537.230 3230.525 ;
        RECT 1537.020 3229.650 1537.160 3230.155 ;
        RECT 1473.020 3229.330 1473.280 3229.650 ;
        RECT 1536.960 3229.330 1537.220 3229.650 ;
        RECT 1459.220 3222.190 1459.480 3222.510 ;
        RECT 1452.320 3215.390 1452.580 3215.710 ;
        RECT 1438.520 3208.590 1438.780 3208.910 ;
        RECT 1431.620 3201.450 1431.880 3201.770 ;
        RECT 1424.720 3194.650 1424.980 3194.970 ;
        RECT 1408.150 2894.915 1408.430 2895.285 ;
        RECT 1408.220 1612.125 1408.360 2894.915 ;
        RECT 1418.740 2794.130 1419.000 2794.450 ;
        RECT 1411.380 2791.070 1411.640 2791.390 ;
        RECT 1410.920 2789.030 1411.180 2789.350 ;
        RECT 1410.460 2152.550 1410.720 2152.870 ;
        RECT 1410.520 2147.285 1410.660 2152.550 ;
        RECT 1410.450 2146.915 1410.730 2147.285 ;
        RECT 1410.460 2131.810 1410.720 2132.130 ;
        RECT 1410.520 2126.885 1410.660 2131.810 ;
        RECT 1410.450 2126.515 1410.730 2126.885 ;
        RECT 1410.460 2117.530 1410.720 2117.850 ;
        RECT 1410.520 2111.925 1410.660 2117.530 ;
        RECT 1410.450 2111.555 1410.730 2111.925 ;
        RECT 1410.460 2096.790 1410.720 2097.110 ;
        RECT 1410.520 2091.525 1410.660 2096.790 ;
        RECT 1410.450 2091.155 1410.730 2091.525 ;
        RECT 1409.540 2090.330 1409.800 2090.650 ;
        RECT 1409.600 2086.765 1409.740 2090.330 ;
        RECT 1409.530 2086.395 1409.810 2086.765 ;
        RECT 1409.540 2080.810 1409.800 2081.130 ;
        RECT 1408.620 2080.470 1408.880 2080.790 ;
        RECT 1408.680 2051.405 1408.820 2080.470 ;
        RECT 1409.080 2080.130 1409.340 2080.450 ;
        RECT 1409.140 2056.165 1409.280 2080.130 ;
        RECT 1409.070 2055.795 1409.350 2056.165 ;
        RECT 1409.600 2053.330 1409.740 2080.810 ;
        RECT 1410.000 2060.070 1410.260 2060.390 ;
        RECT 1410.060 2056.650 1410.200 2060.070 ;
        RECT 1410.000 2056.330 1410.260 2056.650 ;
        RECT 1410.000 2054.290 1410.260 2054.610 ;
        RECT 1409.140 2053.190 1409.740 2053.330 ;
        RECT 1408.610 2051.035 1408.890 2051.405 ;
        RECT 1409.140 2046.645 1409.280 2053.190 ;
        RECT 1409.540 2052.590 1409.800 2052.910 ;
        RECT 1409.070 2046.275 1409.350 2046.645 ;
        RECT 1409.080 2045.790 1409.340 2046.110 ;
        RECT 1409.140 2027.750 1409.280 2045.790 ;
        RECT 1409.600 2036.445 1409.740 2052.590 ;
        RECT 1409.530 2036.075 1409.810 2036.445 ;
        RECT 1409.540 2034.230 1409.800 2034.550 ;
        RECT 1409.080 2027.430 1409.340 2027.750 ;
        RECT 1409.080 2021.485 1409.340 2021.630 ;
        RECT 1409.070 2021.115 1409.350 2021.485 ;
        RECT 1409.600 2015.250 1409.740 2034.230 ;
        RECT 1410.060 2025.710 1410.200 2054.290 ;
        RECT 1410.460 2053.270 1410.720 2053.590 ;
        RECT 1410.000 2025.390 1410.260 2025.710 ;
        RECT 1410.520 2016.045 1410.660 2053.270 ;
        RECT 1410.450 2015.675 1410.730 2016.045 ;
        RECT 1409.600 2015.110 1410.660 2015.250 ;
        RECT 1410.520 2011.285 1410.660 2015.110 ;
        RECT 1410.450 2010.915 1410.730 2011.285 ;
        RECT 1409.530 1965.355 1409.810 1965.725 ;
        RECT 1409.600 1962.470 1409.740 1965.355 ;
        RECT 1409.540 1962.150 1409.800 1962.470 ;
        RECT 1410.460 1956.370 1410.720 1956.690 ;
        RECT 1410.520 1955.525 1410.660 1956.370 ;
        RECT 1410.450 1955.155 1410.730 1955.525 ;
        RECT 1408.620 1895.170 1408.880 1895.490 ;
        RECT 1408.680 1895.005 1408.820 1895.170 ;
        RECT 1408.610 1894.635 1408.890 1895.005 ;
        RECT 1410.460 1869.670 1410.720 1869.990 ;
        RECT 1408.620 1826.830 1408.880 1827.150 ;
        RECT 1408.680 1824.285 1408.820 1826.830 ;
        RECT 1408.610 1823.915 1408.890 1824.285 ;
        RECT 1410.520 1822.050 1410.660 1869.670 ;
        RECT 1410.460 1821.730 1410.720 1822.050 ;
        RECT 1408.620 1819.525 1408.880 1819.670 ;
        RECT 1408.610 1819.155 1408.890 1819.525 ;
        RECT 1408.620 1814.085 1408.880 1814.230 ;
        RECT 1408.610 1813.715 1408.890 1814.085 ;
        RECT 1408.620 1809.325 1408.880 1809.470 ;
        RECT 1408.610 1808.955 1408.890 1809.325 ;
        RECT 1409.080 1799.630 1409.340 1799.950 ;
        RECT 1408.620 1799.125 1408.880 1799.270 ;
        RECT 1408.610 1798.755 1408.890 1799.125 ;
        RECT 1409.140 1794.365 1409.280 1799.630 ;
        RECT 1409.070 1793.995 1409.350 1794.365 ;
        RECT 1408.620 1778.725 1408.880 1778.870 ;
        RECT 1408.610 1778.355 1408.890 1778.725 ;
        RECT 1408.620 1777.870 1408.880 1778.190 ;
        RECT 1408.680 1773.965 1408.820 1777.870 ;
        RECT 1408.610 1773.595 1408.890 1773.965 ;
        RECT 1408.620 1769.370 1408.880 1769.690 ;
        RECT 1408.680 1768.525 1408.820 1769.370 ;
        RECT 1408.610 1768.155 1408.890 1768.525 ;
        RECT 1408.620 1764.950 1408.880 1765.270 ;
        RECT 1408.680 1763.765 1408.820 1764.950 ;
        RECT 1408.610 1763.395 1408.890 1763.765 ;
        RECT 1408.620 1756.450 1408.880 1756.770 ;
        RECT 1408.680 1753.565 1408.820 1756.450 ;
        RECT 1408.610 1753.195 1408.890 1753.565 ;
        RECT 1410.000 1738.090 1410.260 1738.410 ;
        RECT 1410.060 1733.165 1410.200 1738.090 ;
        RECT 1409.990 1732.795 1410.270 1733.165 ;
        RECT 1410.000 1717.690 1410.260 1718.010 ;
        RECT 1410.450 1717.835 1410.730 1718.205 ;
        RECT 1410.060 1713.445 1410.200 1717.690 ;
        RECT 1410.520 1717.670 1410.660 1717.835 ;
        RECT 1410.460 1717.350 1410.720 1717.670 ;
        RECT 1409.990 1713.075 1410.270 1713.445 ;
        RECT 1409.540 1703.245 1409.800 1703.390 ;
        RECT 1409.530 1702.875 1409.810 1703.245 ;
        RECT 1409.080 1699.330 1409.340 1699.650 ;
        RECT 1409.140 1698.485 1409.280 1699.330 ;
        RECT 1409.070 1698.115 1409.350 1698.485 ;
        RECT 1409.540 1694.570 1409.800 1694.890 ;
        RECT 1409.600 1693.045 1409.740 1694.570 ;
        RECT 1409.530 1692.675 1409.810 1693.045 ;
        RECT 1409.540 1688.285 1409.800 1688.430 ;
        RECT 1409.530 1687.915 1409.810 1688.285 ;
        RECT 1410.460 1672.810 1410.720 1673.130 ;
        RECT 1410.520 1672.645 1410.660 1672.810 ;
        RECT 1410.450 1672.275 1410.730 1672.645 ;
        RECT 1409.540 1668.390 1409.800 1668.710 ;
        RECT 1409.600 1667.885 1409.740 1668.390 ;
        RECT 1409.530 1667.515 1409.810 1667.885 ;
        RECT 1410.460 1647.990 1410.720 1648.310 ;
        RECT 1409.540 1647.485 1409.800 1647.630 ;
        RECT 1409.530 1647.115 1409.810 1647.485 ;
        RECT 1410.520 1642.725 1410.660 1647.990 ;
        RECT 1410.450 1642.355 1410.730 1642.725 ;
        RECT 1410.460 1635.070 1410.720 1635.390 ;
        RECT 1410.520 1632.525 1410.660 1635.070 ;
        RECT 1410.450 1632.155 1410.730 1632.525 ;
        RECT 1410.980 1617.565 1411.120 2789.030 ;
        RECT 1411.440 1637.285 1411.580 2791.070 ;
        RECT 1411.840 2790.390 1412.100 2790.710 ;
        RECT 1411.900 1788.925 1412.040 2790.390 ;
        RECT 1417.820 2788.690 1418.080 2789.010 ;
        RECT 1414.140 2145.410 1414.400 2145.730 ;
        RECT 1414.200 2142.525 1414.340 2145.410 ;
        RECT 1414.130 2142.155 1414.410 2142.525 ;
        RECT 1414.140 2138.610 1414.400 2138.930 ;
        RECT 1413.680 2138.270 1413.940 2138.590 ;
        RECT 1413.740 2132.325 1413.880 2138.270 ;
        RECT 1414.200 2137.085 1414.340 2138.610 ;
        RECT 1414.130 2136.715 1414.410 2137.085 ;
        RECT 1413.670 2131.955 1413.950 2132.325 ;
        RECT 1414.140 2125.010 1414.400 2125.330 ;
        RECT 1414.200 2122.125 1414.340 2125.010 ;
        RECT 1414.130 2121.755 1414.410 2122.125 ;
        RECT 1414.140 2117.870 1414.400 2118.190 ;
        RECT 1414.200 2117.365 1414.340 2117.870 ;
        RECT 1414.130 2116.995 1414.410 2117.365 ;
        RECT 1414.140 2111.070 1414.400 2111.390 ;
        RECT 1414.200 2107.165 1414.340 2111.070 ;
        RECT 1414.130 2106.795 1414.410 2107.165 ;
        RECT 1414.140 2104.270 1414.400 2104.590 ;
        RECT 1414.200 2101.725 1414.340 2104.270 ;
        RECT 1414.130 2101.355 1414.410 2101.725 ;
        RECT 1414.140 2097.130 1414.400 2097.450 ;
        RECT 1414.200 2096.965 1414.340 2097.130 ;
        RECT 1414.130 2096.595 1414.410 2096.965 ;
        RECT 1416.900 2086.930 1417.160 2087.250 ;
        RECT 1414.140 2083.530 1414.400 2083.850 ;
        RECT 1412.760 2082.510 1413.020 2082.830 ;
        RECT 1412.300 2082.170 1412.560 2082.490 ;
        RECT 1412.360 2063.450 1412.500 2082.170 ;
        RECT 1412.300 2063.130 1412.560 2063.450 ;
        RECT 1412.300 2053.950 1412.560 2054.270 ;
        RECT 1412.360 2028.430 1412.500 2053.950 ;
        RECT 1412.300 2028.110 1412.560 2028.430 ;
        RECT 1412.300 2027.430 1412.560 2027.750 ;
        RECT 1411.830 1788.555 1412.110 1788.925 ;
        RECT 1411.840 1682.845 1412.100 1682.990 ;
        RECT 1411.830 1682.475 1412.110 1682.845 ;
        RECT 1411.840 1678.085 1412.100 1678.230 ;
        RECT 1411.830 1677.715 1412.110 1678.085 ;
        RECT 1411.840 1669.410 1412.100 1669.730 ;
        RECT 1411.900 1663.125 1412.040 1669.410 ;
        RECT 1411.830 1662.755 1412.110 1663.125 ;
        RECT 1411.370 1636.915 1411.650 1637.285 ;
        RECT 1412.360 1622.325 1412.500 2027.430 ;
        RECT 1412.820 1748.805 1412.960 2082.510 ;
        RECT 1414.200 2082.005 1414.340 2083.530 ;
        RECT 1414.130 2081.635 1414.410 2082.005 ;
        RECT 1414.600 2081.150 1414.860 2081.470 ;
        RECT 1414.140 2076.730 1414.400 2077.050 ;
        RECT 1413.680 2076.390 1413.940 2076.710 ;
        RECT 1414.200 2076.565 1414.340 2076.730 ;
        RECT 1413.740 2071.805 1413.880 2076.390 ;
        RECT 1414.130 2076.195 1414.410 2076.565 ;
        RECT 1413.670 2071.435 1413.950 2071.805 ;
        RECT 1414.140 2069.590 1414.400 2069.910 ;
        RECT 1414.200 2066.365 1414.340 2069.590 ;
        RECT 1414.130 2065.995 1414.410 2066.365 ;
        RECT 1413.680 2063.130 1413.940 2063.450 ;
        RECT 1413.220 2052.930 1413.480 2053.250 ;
        RECT 1413.280 2026.245 1413.420 2052.930 ;
        RECT 1413.210 2025.875 1413.490 2026.245 ;
        RECT 1413.220 2025.390 1413.480 2025.710 ;
        RECT 1413.280 2014.830 1413.420 2025.390 ;
        RECT 1413.220 2014.510 1413.480 2014.830 ;
        RECT 1413.740 2001.085 1413.880 2063.130 ;
        RECT 1414.140 2062.790 1414.400 2063.110 ;
        RECT 1414.200 2061.605 1414.340 2062.790 ;
        RECT 1414.130 2061.235 1414.410 2061.605 ;
        RECT 1414.140 2053.610 1414.400 2053.930 ;
        RECT 1414.200 2034.550 1414.340 2053.610 ;
        RECT 1414.660 2041.205 1414.800 2081.150 ;
        RECT 1416.440 2068.570 1416.700 2068.890 ;
        RECT 1415.980 2068.230 1416.240 2068.550 ;
        RECT 1415.520 2067.210 1415.780 2067.530 ;
        RECT 1415.060 2066.190 1415.320 2066.510 ;
        RECT 1414.590 2040.835 1414.870 2041.205 ;
        RECT 1414.140 2034.230 1414.400 2034.550 ;
        RECT 1414.130 2030.635 1414.410 2031.005 ;
        RECT 1414.200 2029.110 1414.340 2030.635 ;
        RECT 1414.140 2028.790 1414.400 2029.110 ;
        RECT 1414.140 2028.110 1414.400 2028.430 ;
        RECT 1414.200 2005.845 1414.340 2028.110 ;
        RECT 1414.600 2014.510 1414.860 2014.830 ;
        RECT 1414.130 2005.475 1414.410 2005.845 ;
        RECT 1414.660 2005.050 1414.800 2014.510 ;
        RECT 1414.200 2004.910 1414.800 2005.050 ;
        RECT 1413.670 2000.715 1413.950 2001.085 ;
        RECT 1414.200 2000.290 1414.340 2004.910 ;
        RECT 1413.740 2000.150 1414.340 2000.290 ;
        RECT 1413.740 1952.010 1413.880 2000.150 ;
        RECT 1414.140 1995.810 1414.400 1996.130 ;
        RECT 1414.200 1995.645 1414.340 1995.810 ;
        RECT 1414.130 1995.275 1414.410 1995.645 ;
        RECT 1414.130 1990.515 1414.410 1990.885 ;
        RECT 1414.200 1989.670 1414.340 1990.515 ;
        RECT 1414.140 1989.350 1414.400 1989.670 ;
        RECT 1414.130 1985.755 1414.410 1986.125 ;
        RECT 1414.200 1984.570 1414.340 1985.755 ;
        RECT 1414.140 1984.250 1414.400 1984.570 ;
        RECT 1414.140 1981.190 1414.400 1981.510 ;
        RECT 1414.200 1980.685 1414.340 1981.190 ;
        RECT 1414.130 1980.315 1414.410 1980.685 ;
        RECT 1414.130 1975.555 1414.410 1975.925 ;
        RECT 1414.200 1974.030 1414.340 1975.555 ;
        RECT 1414.140 1973.710 1414.400 1974.030 ;
        RECT 1414.130 1970.115 1414.410 1970.485 ;
        RECT 1414.200 1969.610 1414.340 1970.115 ;
        RECT 1414.140 1969.290 1414.400 1969.610 ;
        RECT 1414.140 1961.470 1414.400 1961.790 ;
        RECT 1414.200 1960.285 1414.340 1961.470 ;
        RECT 1414.130 1959.915 1414.410 1960.285 ;
        RECT 1413.740 1951.870 1414.340 1952.010 ;
        RECT 1413.680 1951.270 1413.940 1951.590 ;
        RECT 1413.740 1950.765 1413.880 1951.270 ;
        RECT 1413.670 1950.395 1413.950 1950.765 ;
        RECT 1413.680 1945.325 1413.940 1945.470 ;
        RECT 1413.670 1944.955 1413.950 1945.325 ;
        RECT 1413.680 1942.770 1413.940 1943.090 ;
        RECT 1413.740 1940.565 1413.880 1942.770 ;
        RECT 1413.670 1940.195 1413.950 1940.565 ;
        RECT 1413.680 1936.310 1413.940 1936.630 ;
        RECT 1413.740 1935.125 1413.880 1936.310 ;
        RECT 1413.670 1934.755 1413.950 1935.125 ;
        RECT 1413.680 1930.365 1413.940 1930.510 ;
        RECT 1413.670 1929.995 1413.950 1930.365 ;
        RECT 1413.680 1926.450 1413.940 1926.770 ;
        RECT 1413.740 1925.605 1413.880 1926.450 ;
        RECT 1413.670 1925.235 1413.950 1925.605 ;
        RECT 1414.200 1923.450 1414.340 1951.870 ;
        RECT 1413.740 1923.310 1414.340 1923.450 ;
        RECT 1413.740 1894.210 1413.880 1923.310 ;
        RECT 1414.130 1922.770 1414.410 1922.885 ;
        RECT 1415.120 1922.770 1415.260 2066.190 ;
        RECT 1414.130 1922.630 1415.260 1922.770 ;
        RECT 1414.130 1922.515 1414.410 1922.630 ;
        RECT 1414.140 1915.405 1414.400 1915.550 ;
        RECT 1414.130 1915.035 1414.410 1915.405 ;
        RECT 1414.130 1910.530 1414.410 1910.645 ;
        RECT 1415.580 1910.530 1415.720 2067.210 ;
        RECT 1414.130 1910.390 1415.720 1910.530 ;
        RECT 1414.130 1910.275 1414.410 1910.390 ;
        RECT 1414.140 1906.390 1414.400 1906.710 ;
        RECT 1414.200 1905.205 1414.340 1906.390 ;
        RECT 1414.130 1904.835 1414.410 1905.205 ;
        RECT 1414.130 1901.010 1414.410 1901.125 ;
        RECT 1416.040 1901.010 1416.180 2068.230 ;
        RECT 1414.130 1900.870 1416.180 1901.010 ;
        RECT 1414.130 1900.755 1414.410 1900.870 ;
        RECT 1416.500 1895.490 1416.640 2068.570 ;
        RECT 1416.440 1895.170 1416.700 1895.490 ;
        RECT 1413.280 1894.070 1413.880 1894.210 ;
        RECT 1413.280 1869.990 1413.420 1894.070 ;
        RECT 1414.140 1890.245 1414.400 1890.390 ;
        RECT 1414.130 1889.875 1414.410 1890.245 ;
        RECT 1414.140 1885.650 1414.400 1885.970 ;
        RECT 1414.200 1884.805 1414.340 1885.650 ;
        RECT 1414.130 1884.435 1414.410 1884.805 ;
        RECT 1414.140 1881.570 1414.400 1881.890 ;
        RECT 1414.200 1880.045 1414.340 1881.570 ;
        RECT 1414.130 1879.675 1414.410 1880.045 ;
        RECT 1414.130 1874.235 1414.410 1874.605 ;
        RECT 1414.200 1872.710 1414.340 1874.235 ;
        RECT 1414.140 1872.390 1414.400 1872.710 ;
        RECT 1413.220 1869.670 1413.480 1869.990 ;
        RECT 1413.680 1869.670 1413.940 1869.990 ;
        RECT 1413.740 1864.405 1413.880 1869.670 ;
        RECT 1414.130 1869.475 1414.410 1869.845 ;
        RECT 1414.200 1865.910 1414.340 1869.475 ;
        RECT 1414.140 1865.590 1414.400 1865.910 ;
        RECT 1413.670 1864.035 1413.950 1864.405 ;
        RECT 1414.130 1859.275 1414.410 1859.645 ;
        RECT 1414.200 1858.430 1414.340 1859.275 ;
        RECT 1414.140 1858.110 1414.400 1858.430 ;
        RECT 1414.140 1855.730 1414.400 1856.050 ;
        RECT 1413.680 1855.390 1413.940 1855.710 ;
        RECT 1413.740 1849.445 1413.880 1855.390 ;
        RECT 1414.200 1854.885 1414.340 1855.730 ;
        RECT 1414.130 1854.515 1414.410 1854.885 ;
        RECT 1413.670 1849.075 1413.950 1849.445 ;
        RECT 1414.140 1848.930 1414.400 1849.250 ;
        RECT 1414.200 1844.685 1414.340 1848.930 ;
        RECT 1414.130 1844.315 1414.410 1844.685 ;
        RECT 1414.140 1840.770 1414.400 1841.090 ;
        RECT 1414.200 1839.245 1414.340 1840.770 ;
        RECT 1414.130 1838.875 1414.410 1839.245 ;
        RECT 1414.140 1834.990 1414.400 1835.310 ;
        RECT 1414.200 1834.485 1414.340 1834.990 ;
        RECT 1414.130 1834.115 1414.410 1834.485 ;
        RECT 1414.140 1830.910 1414.400 1831.230 ;
        RECT 1414.200 1829.045 1414.340 1830.910 ;
        RECT 1414.130 1828.675 1414.410 1829.045 ;
        RECT 1413.220 1821.730 1413.480 1822.050 ;
        RECT 1413.280 1759.005 1413.420 1821.730 ;
        RECT 1416.960 1819.670 1417.100 2086.930 ;
        RECT 1417.360 2079.110 1417.620 2079.430 ;
        RECT 1416.900 1819.350 1417.160 1819.670 ;
        RECT 1414.140 1807.450 1414.400 1807.770 ;
        RECT 1414.200 1803.885 1414.340 1807.450 ;
        RECT 1414.130 1803.515 1414.410 1803.885 ;
        RECT 1417.420 1799.270 1417.560 2079.110 ;
        RECT 1417.360 1798.950 1417.620 1799.270 ;
        RECT 1414.130 1783.795 1414.410 1784.165 ;
        RECT 1414.200 1783.290 1414.340 1783.795 ;
        RECT 1414.140 1782.970 1414.400 1783.290 ;
        RECT 1413.210 1758.635 1413.490 1759.005 ;
        RECT 1417.880 1756.770 1418.020 2788.690 ;
        RECT 1418.280 2788.350 1418.540 2788.670 ;
        RECT 1418.340 1765.270 1418.480 2788.350 ;
        RECT 1418.800 1769.690 1418.940 2794.130 ;
        RECT 1419.200 2793.790 1419.460 2794.110 ;
        RECT 1419.260 1778.870 1419.400 2793.790 ;
        RECT 1420.580 2792.090 1420.840 2792.410 ;
        RECT 1420.120 2790.050 1420.380 2790.370 ;
        RECT 1419.660 2789.710 1419.920 2790.030 ;
        RECT 1419.720 1814.230 1419.860 2789.710 ;
        RECT 1419.660 1813.910 1419.920 1814.230 ;
        RECT 1420.180 1809.470 1420.320 2790.050 ;
        RECT 1420.640 1827.150 1420.780 2792.090 ;
        RECT 1422.420 2087.270 1422.680 2087.590 ;
        RECT 1421.960 2081.490 1422.220 2081.810 ;
        RECT 1421.040 2059.390 1421.300 2059.710 ;
        RECT 1420.580 1826.830 1420.840 1827.150 ;
        RECT 1420.120 1809.150 1420.380 1809.470 ;
        RECT 1419.200 1778.550 1419.460 1778.870 ;
        RECT 1421.100 1778.190 1421.240 2059.390 ;
        RECT 1422.020 2021.630 1422.160 2081.490 ;
        RECT 1421.960 2021.310 1422.220 2021.630 ;
        RECT 1422.480 1799.950 1422.620 2087.270 ;
        RECT 1423.340 2062.110 1423.600 2062.430 ;
        RECT 1422.880 2061.090 1423.140 2061.410 ;
        RECT 1422.420 1799.630 1422.680 1799.950 ;
        RECT 1421.040 1777.870 1421.300 1778.190 ;
        RECT 1418.740 1769.370 1419.000 1769.690 ;
        RECT 1418.280 1764.950 1418.540 1765.270 ;
        RECT 1417.820 1756.450 1418.080 1756.770 ;
        RECT 1412.750 1748.435 1413.030 1748.805 ;
        RECT 1414.140 1745.230 1414.400 1745.550 ;
        RECT 1414.200 1743.365 1414.340 1745.230 ;
        RECT 1414.130 1742.995 1414.410 1743.365 ;
        RECT 1414.140 1738.605 1414.400 1738.750 ;
        RECT 1414.130 1738.235 1414.410 1738.605 ;
        RECT 1414.140 1728.910 1414.400 1729.230 ;
        RECT 1414.200 1728.405 1414.340 1728.910 ;
        RECT 1414.130 1728.035 1414.410 1728.405 ;
        RECT 1413.680 1723.645 1413.940 1723.790 ;
        RECT 1413.670 1723.275 1413.950 1723.645 ;
        RECT 1414.140 1710.890 1414.400 1711.210 ;
        RECT 1414.200 1708.005 1414.340 1710.890 ;
        RECT 1414.130 1707.635 1414.410 1708.005 ;
        RECT 1422.940 1699.650 1423.080 2061.090 ;
        RECT 1423.400 1703.390 1423.540 2062.110 ;
        RECT 1423.800 2061.770 1424.060 2062.090 ;
        RECT 1423.340 1703.070 1423.600 1703.390 ;
        RECT 1422.880 1699.330 1423.140 1699.650 ;
        RECT 1423.860 1694.890 1424.000 2061.770 ;
        RECT 1424.260 2061.430 1424.520 2061.750 ;
        RECT 1423.800 1694.570 1424.060 1694.890 ;
        RECT 1424.320 1688.430 1424.460 2061.430 ;
        RECT 1424.780 1717.670 1424.920 3194.650 ;
        RECT 1425.180 2790.730 1425.440 2791.050 ;
        RECT 1424.720 1717.350 1424.980 1717.670 ;
        RECT 1424.260 1688.110 1424.520 1688.430 ;
        RECT 1414.140 1655.810 1414.400 1656.130 ;
        RECT 1414.200 1652.925 1414.340 1655.810 ;
        RECT 1414.130 1652.555 1414.410 1652.925 ;
        RECT 1425.240 1647.630 1425.380 2790.730 ;
        RECT 1425.640 2087.610 1425.900 2087.930 ;
        RECT 1425.700 1648.310 1425.840 2087.610 ;
        RECT 1429.780 2076.050 1430.040 2076.370 ;
        RECT 1428.860 2075.370 1429.120 2075.690 ;
        RECT 1428.400 2074.350 1428.660 2074.670 ;
        RECT 1427.020 2062.450 1427.280 2062.770 ;
        RECT 1426.560 2060.750 1426.820 2061.070 ;
        RECT 1426.100 2060.410 1426.360 2060.730 ;
        RECT 1425.640 1647.990 1425.900 1648.310 ;
        RECT 1425.180 1647.310 1425.440 1647.630 ;
        RECT 1426.160 1635.390 1426.300 2060.410 ;
        RECT 1426.620 1668.710 1426.760 2060.750 ;
        RECT 1427.080 1673.130 1427.220 2062.450 ;
        RECT 1427.480 2059.050 1427.740 2059.370 ;
        RECT 1427.540 1682.990 1427.680 2059.050 ;
        RECT 1427.940 2058.710 1428.200 2059.030 ;
        RECT 1427.480 1682.670 1427.740 1682.990 ;
        RECT 1428.000 1678.230 1428.140 2058.710 ;
        RECT 1428.460 1956.690 1428.600 2074.350 ;
        RECT 1428.400 1956.370 1428.660 1956.690 ;
        RECT 1428.920 1951.590 1429.060 2075.370 ;
        RECT 1429.320 2066.530 1429.580 2066.850 ;
        RECT 1428.860 1951.270 1429.120 1951.590 ;
        RECT 1429.380 1936.630 1429.520 2066.530 ;
        RECT 1429.840 1945.470 1429.980 2076.050 ;
        RECT 1430.240 2072.990 1430.500 2073.310 ;
        RECT 1429.780 1945.150 1430.040 1945.470 ;
        RECT 1430.300 1943.090 1430.440 2072.990 ;
        RECT 1430.700 2067.550 1430.960 2067.870 ;
        RECT 1430.240 1942.770 1430.500 1943.090 ;
        RECT 1429.320 1936.310 1429.580 1936.630 ;
        RECT 1430.760 1926.770 1430.900 2067.550 ;
        RECT 1431.160 2066.870 1431.420 2067.190 ;
        RECT 1431.220 1930.510 1431.360 2066.870 ;
        RECT 1431.160 1930.190 1431.420 1930.510 ;
        RECT 1430.700 1926.450 1430.960 1926.770 ;
        RECT 1431.680 1723.790 1431.820 3201.450 ;
        RECT 1436.680 2083.190 1436.940 2083.510 ;
        RECT 1436.220 2082.850 1436.480 2083.170 ;
        RECT 1435.760 2081.830 1436.020 2082.150 ;
        RECT 1432.540 2072.310 1432.800 2072.630 ;
        RECT 1432.080 2065.170 1432.340 2065.490 ;
        RECT 1432.140 1831.230 1432.280 2065.170 ;
        RECT 1432.600 1841.090 1432.740 2072.310 ;
        RECT 1433.460 2069.250 1433.720 2069.570 ;
        RECT 1433.000 2065.510 1433.260 2065.830 ;
        RECT 1433.060 1881.890 1433.200 2065.510 ;
        RECT 1433.520 1890.390 1433.660 2069.250 ;
        RECT 1434.380 2068.910 1434.640 2069.230 ;
        RECT 1433.920 2065.850 1434.180 2066.170 ;
        RECT 1433.460 1890.070 1433.720 1890.390 ;
        RECT 1433.980 1885.970 1434.120 2065.850 ;
        RECT 1434.440 1906.710 1434.580 2068.910 ;
        RECT 1434.840 2067.890 1435.100 2068.210 ;
        RECT 1434.900 1915.550 1435.040 2067.890 ;
        RECT 1435.820 2029.110 1435.960 2081.830 ;
        RECT 1435.760 2028.790 1436.020 2029.110 ;
        RECT 1436.280 1996.130 1436.420 2082.850 ;
        RECT 1436.220 1995.810 1436.480 1996.130 ;
        RECT 1436.740 1989.670 1436.880 2083.190 ;
        RECT 1438.060 2074.010 1438.320 2074.330 ;
        RECT 1437.600 2073.670 1437.860 2073.990 ;
        RECT 1437.140 2073.330 1437.400 2073.650 ;
        RECT 1436.680 1989.350 1436.940 1989.670 ;
        RECT 1437.200 1984.570 1437.340 2073.330 ;
        RECT 1437.140 1984.250 1437.400 1984.570 ;
        RECT 1437.660 1981.510 1437.800 2073.670 ;
        RECT 1437.600 1981.190 1437.860 1981.510 ;
        RECT 1438.120 1974.030 1438.260 2074.010 ;
        RECT 1438.060 1973.710 1438.320 1974.030 ;
        RECT 1434.840 1915.230 1435.100 1915.550 ;
        RECT 1434.380 1906.390 1434.640 1906.710 ;
        RECT 1433.920 1885.650 1434.180 1885.970 ;
        RECT 1433.000 1881.570 1433.260 1881.890 ;
        RECT 1432.540 1840.770 1432.800 1841.090 ;
        RECT 1432.080 1830.910 1432.340 1831.230 ;
        RECT 1438.580 1729.230 1438.720 3208.590 ;
        RECT 1440.360 2079.790 1440.620 2080.110 ;
        RECT 1439.440 2079.450 1439.700 2079.770 ;
        RECT 1438.980 2059.730 1439.240 2060.050 ;
        RECT 1439.040 1783.290 1439.180 2059.730 ;
        RECT 1439.500 1865.910 1439.640 2079.450 ;
        RECT 1439.900 2072.650 1440.160 2072.970 ;
        RECT 1439.440 1865.590 1439.700 1865.910 ;
        RECT 1439.960 1858.430 1440.100 2072.650 ;
        RECT 1440.420 1872.710 1440.560 2079.790 ;
        RECT 1440.820 2075.710 1441.080 2076.030 ;
        RECT 1440.880 1961.790 1441.020 2075.710 ;
        RECT 1441.280 2075.030 1441.540 2075.350 ;
        RECT 1441.340 1962.470 1441.480 2075.030 ;
        RECT 1441.740 2074.690 1442.000 2075.010 ;
        RECT 1441.800 1969.610 1441.940 2074.690 ;
        RECT 1441.740 1969.290 1442.000 1969.610 ;
        RECT 1441.280 1962.150 1441.540 1962.470 ;
        RECT 1440.820 1961.470 1441.080 1961.790 ;
        RECT 1440.360 1872.390 1440.620 1872.710 ;
        RECT 1439.900 1858.110 1440.160 1858.430 ;
        RECT 1438.980 1782.970 1439.240 1783.290 ;
        RECT 1452.380 1738.410 1452.520 3215.390 ;
        RECT 1459.280 1738.750 1459.420 3222.190 ;
        RECT 1459.680 2898.170 1459.940 2898.490 ;
        RECT 1459.220 1738.430 1459.480 1738.750 ;
        RECT 1452.320 1738.090 1452.580 1738.410 ;
        RECT 1438.520 1728.910 1438.780 1729.230 ;
        RECT 1431.620 1723.470 1431.880 1723.790 ;
        RECT 1427.940 1677.910 1428.200 1678.230 ;
        RECT 1427.020 1672.810 1427.280 1673.130 ;
        RECT 1459.740 1669.730 1459.880 2898.170 ;
        RECT 1466.120 2064.830 1466.380 2065.150 ;
        RECT 1460.140 2058.370 1460.400 2058.690 ;
        RECT 1459.680 1669.410 1459.940 1669.730 ;
        RECT 1426.560 1668.390 1426.820 1668.710 ;
        RECT 1460.200 1656.130 1460.340 2058.370 ;
        RECT 1466.180 1835.310 1466.320 2064.830 ;
        RECT 1466.120 1834.990 1466.380 1835.310 ;
        RECT 1473.080 1745.550 1473.220 3229.330 ;
        RECT 1535.570 3224.715 1535.850 3225.085 ;
        RECT 1535.640 3222.510 1535.780 3224.715 ;
        RECT 1535.580 3222.190 1535.840 3222.510 ;
        RECT 1535.570 3217.235 1535.850 3217.605 ;
        RECT 1535.640 3215.710 1535.780 3217.235 ;
        RECT 1535.580 3215.390 1535.840 3215.710 ;
        RECT 1538.330 3210.435 1538.610 3210.805 ;
        RECT 1538.400 3208.910 1538.540 3210.435 ;
        RECT 1538.340 3208.590 1538.600 3208.910 ;
        RECT 1538.330 3202.275 1538.610 3202.645 ;
        RECT 1538.400 3201.770 1538.540 3202.275 ;
        RECT 1538.340 3201.450 1538.600 3201.770 ;
        RECT 1533.270 3196.835 1533.550 3197.205 ;
        RECT 1533.340 3194.970 1533.480 3196.835 ;
        RECT 1533.280 3194.650 1533.540 3194.970 ;
        RECT 1534.190 3189.355 1534.470 3189.725 ;
        RECT 1534.260 3188.170 1534.400 3189.355 ;
        RECT 1473.480 3187.850 1473.740 3188.170 ;
        RECT 1534.200 3187.850 1534.460 3188.170 ;
        RECT 1473.020 1745.230 1473.280 1745.550 ;
        RECT 1473.540 1718.010 1473.680 3187.850 ;
        RECT 1538.330 2898.995 1538.610 2899.365 ;
        RECT 1538.400 2898.490 1538.540 2898.995 ;
        RECT 1538.340 2898.170 1538.600 2898.490 ;
      LAYER met2 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met2 ;
        RECT 1935.780 3251.090 1936.040 3251.410 ;
        RECT 1935.840 3249.565 1935.980 3251.090 ;
        RECT 1935.770 3249.195 1936.050 3249.565 ;
        RECT 2190.610 3230.155 2190.890 3230.525 ;
        RECT 1732.910 2795.635 1733.190 2796.005 ;
        RECT 1732.980 2795.130 1733.120 2795.635 ;
        RECT 1732.920 2794.810 1733.180 2795.130 ;
        RECT 1613.310 2794.275 1613.590 2794.645 ;
        RECT 1642.750 2794.275 1643.030 2794.645 ;
        RECT 1652.870 2794.275 1653.150 2794.645 ;
        RECT 1659.310 2794.275 1659.590 2794.645 ;
        RECT 1669.430 2794.275 1669.710 2794.645 ;
        RECT 1670.350 2794.275 1670.630 2794.645 ;
        RECT 1677.250 2794.275 1677.530 2794.645 ;
        RECT 1695.190 2794.275 1695.470 2794.645 ;
        RECT 1699.330 2794.275 1699.610 2794.645 ;
        RECT 1706.230 2794.275 1706.510 2794.645 ;
        RECT 1712.670 2794.275 1712.950 2794.645 ;
        RECT 1718.190 2794.275 1718.470 2794.645 ;
        RECT 1723.710 2794.275 1723.990 2794.645 ;
        RECT 1728.770 2794.275 1729.050 2794.645 ;
        RECT 1741.190 2794.275 1741.470 2794.645 ;
        RECT 1747.630 2794.275 1747.910 2794.645 ;
        RECT 1760.050 2794.275 1760.330 2794.645 ;
        RECT 1596.290 2792.235 1596.570 2792.605 ;
        RECT 1596.360 2792.070 1596.500 2792.235 ;
        RECT 1549.380 2791.750 1549.640 2792.070 ;
        RECT 1548.920 2787.670 1549.180 2787.990 ;
        RECT 1494.180 2078.770 1494.440 2079.090 ;
        RECT 1493.720 2058.030 1493.980 2058.350 ;
        RECT 1473.480 1717.690 1473.740 1718.010 ;
        RECT 1493.780 1711.210 1493.920 2058.030 ;
        RECT 1494.240 1807.770 1494.380 2078.770 ;
        RECT 1494.640 2071.970 1494.900 2072.290 ;
        RECT 1494.700 1869.990 1494.840 2071.970 ;
        RECT 1494.640 1869.670 1494.900 1869.990 ;
        RECT 1548.980 1849.250 1549.120 2787.670 ;
        RECT 1549.440 1855.710 1549.580 2791.750 ;
        RECT 1587.090 2791.555 1587.370 2791.925 ;
        RECT 1596.300 2791.750 1596.560 2792.070 ;
        RECT 1600.890 2791.555 1601.170 2791.925 ;
        RECT 1587.160 2791.390 1587.300 2791.555 ;
        RECT 1587.100 2791.070 1587.360 2791.390 ;
        RECT 1600.960 2791.050 1601.100 2791.555 ;
        RECT 1600.900 2790.730 1601.160 2791.050 ;
        RECT 1613.380 2790.710 1613.520 2794.275 ;
        RECT 1642.820 2793.770 1642.960 2794.275 ;
        RECT 1642.760 2793.450 1643.020 2793.770 ;
        RECT 1636.770 2792.915 1637.050 2793.285 ;
        RECT 1613.320 2790.390 1613.580 2790.710 ;
        RECT 1624.820 2790.390 1625.080 2790.710 ;
        RECT 1549.840 2789.370 1550.100 2789.690 ;
        RECT 1549.900 1856.050 1550.040 2789.370 ;
        RECT 1624.880 2788.525 1625.020 2790.390 ;
        RECT 1636.840 2790.370 1636.980 2792.915 ;
        RECT 1636.780 2790.050 1637.040 2790.370 ;
        RECT 1642.290 2790.195 1642.570 2790.565 ;
        RECT 1642.360 2789.690 1642.500 2790.195 ;
        RECT 1642.820 2790.030 1642.960 2793.450 ;
        RECT 1652.940 2792.750 1653.080 2794.275 ;
        RECT 1652.880 2792.430 1653.140 2792.750 ;
        RECT 1659.380 2791.050 1659.520 2794.275 ;
        RECT 1662.540 2792.090 1662.800 2792.410 ;
        RECT 1662.600 2791.050 1662.740 2792.090 ;
        RECT 1669.500 2791.050 1669.640 2794.275 ;
        RECT 1670.420 2791.390 1670.560 2794.275 ;
        RECT 1677.320 2793.090 1677.460 2794.275 ;
        RECT 1688.750 2793.850 1689.030 2793.965 ;
        RECT 1687.900 2793.770 1689.420 2793.850 ;
        RECT 1687.840 2793.710 1689.480 2793.770 ;
        RECT 1687.840 2793.450 1688.100 2793.710 ;
        RECT 1688.750 2793.595 1689.030 2793.710 ;
        RECT 1688.820 2793.295 1688.960 2793.595 ;
        RECT 1689.220 2793.450 1689.480 2793.710 ;
        RECT 1677.260 2792.770 1677.520 2793.090 ;
        RECT 1682.310 2792.915 1682.590 2793.285 ;
        RECT 1670.360 2791.070 1670.620 2791.390 ;
        RECT 1659.320 2790.730 1659.580 2791.050 ;
        RECT 1662.540 2790.730 1662.800 2791.050 ;
        RECT 1669.440 2790.730 1669.700 2791.050 ;
        RECT 1642.760 2789.710 1643.020 2790.030 ;
        RECT 1642.300 2789.370 1642.560 2789.690 ;
        RECT 1645.520 2789.370 1645.780 2789.690 ;
        RECT 1648.270 2789.515 1648.550 2789.885 ;
        RECT 1648.280 2789.370 1648.540 2789.515 ;
        RECT 1617.910 2788.155 1618.190 2788.525 ;
        RECT 1624.810 2788.155 1625.090 2788.525 ;
        RECT 1628.490 2788.155 1628.770 2788.525 ;
        RECT 1617.920 2788.010 1618.180 2788.155 ;
        RECT 1580.190 2787.475 1580.470 2787.845 ;
        RECT 1593.990 2787.475 1594.270 2787.845 ;
        RECT 1601.350 2787.475 1601.630 2787.845 ;
        RECT 1607.790 2787.475 1608.070 2787.845 ;
        RECT 1614.690 2787.475 1614.970 2787.845 ;
        RECT 1580.260 2058.350 1580.400 2787.475 ;
        RECT 1594.060 2087.930 1594.200 2787.475 ;
        RECT 1594.000 2087.610 1594.260 2087.930 ;
        RECT 1601.420 2058.690 1601.560 2787.475 ;
        RECT 1607.860 2065.490 1608.000 2787.475 ;
        RECT 1607.800 2065.170 1608.060 2065.490 ;
        RECT 1614.760 2065.150 1614.900 2787.475 ;
        RECT 1617.980 2087.590 1618.120 2788.010 ;
        RECT 1621.590 2787.475 1621.870 2787.845 ;
        RECT 1617.920 2087.270 1618.180 2087.590 ;
        RECT 1621.660 2072.630 1621.800 2787.475 ;
        RECT 1624.880 2079.430 1625.020 2788.155 ;
        RECT 1628.560 2787.990 1628.700 2788.155 ;
        RECT 1631.780 2787.990 1631.920 2788.145 ;
        RECT 1628.500 2787.670 1628.760 2787.990 ;
        RECT 1631.720 2787.845 1631.980 2787.990 ;
        RECT 1631.710 2787.475 1631.990 2787.845 ;
        RECT 1624.820 2079.110 1625.080 2079.430 ;
        RECT 1631.780 2079.090 1631.920 2787.475 ;
        RECT 1645.580 2087.250 1645.720 2789.370 ;
        RECT 1649.650 2788.155 1649.930 2788.525 ;
        RECT 1669.500 2788.330 1669.640 2790.730 ;
        RECT 1649.190 2787.475 1649.470 2787.845 ;
        RECT 1645.520 2086.930 1645.780 2087.250 ;
        RECT 1631.720 2078.770 1631.980 2079.090 ;
        RECT 1649.260 2072.970 1649.400 2787.475 ;
        RECT 1649.200 2072.650 1649.460 2072.970 ;
        RECT 1621.600 2072.310 1621.860 2072.630 ;
        RECT 1649.720 2072.290 1649.860 2788.155 ;
        RECT 1669.440 2788.010 1669.700 2788.330 ;
        RECT 1677.320 2787.990 1677.460 2792.770 ;
        RECT 1682.380 2791.730 1682.520 2792.915 ;
        RECT 1695.260 2792.750 1695.400 2794.275 ;
        RECT 1690.600 2792.430 1690.860 2792.750 ;
        RECT 1695.200 2792.430 1695.460 2792.750 ;
        RECT 1682.320 2791.410 1682.580 2791.730 ;
        RECT 1690.660 2789.690 1690.800 2792.430 ;
        RECT 1699.400 2792.070 1699.540 2794.275 ;
        RECT 1706.300 2792.410 1706.440 2794.275 ;
        RECT 1706.240 2792.090 1706.500 2792.410 ;
        RECT 1699.340 2791.750 1699.600 2792.070 ;
        RECT 1712.740 2791.050 1712.880 2794.275 ;
        RECT 1718.260 2791.390 1718.400 2794.275 ;
        RECT 1723.780 2793.770 1723.920 2794.275 ;
        RECT 1723.720 2793.450 1723.980 2793.770 ;
        RECT 1723.780 2793.090 1723.920 2793.450 ;
        RECT 1723.720 2792.770 1723.980 2793.090 ;
        RECT 1728.840 2791.730 1728.980 2794.275 ;
        RECT 1741.260 2793.090 1741.400 2794.275 ;
        RECT 1741.200 2792.770 1741.460 2793.090 ;
        RECT 1728.780 2791.410 1729.040 2791.730 ;
        RECT 1718.200 2791.070 1718.460 2791.390 ;
        RECT 1724.640 2791.070 1724.900 2791.390 ;
        RECT 1712.680 2790.730 1712.940 2791.050 ;
        RECT 1724.700 2790.710 1724.840 2791.070 ;
        RECT 1724.640 2790.390 1724.900 2790.710 ;
        RECT 1741.260 2790.370 1741.400 2792.770 ;
        RECT 1747.700 2791.730 1747.840 2794.275 ;
        RECT 1752.690 2792.235 1752.970 2792.605 ;
        RECT 1752.700 2792.090 1752.960 2792.235 ;
        RECT 1747.640 2791.410 1747.900 2791.730 ;
        RECT 1759.590 2791.555 1759.870 2791.925 ;
        RECT 1759.660 2791.050 1759.800 2791.555 ;
        RECT 1759.600 2790.730 1759.860 2791.050 ;
        RECT 1760.120 2790.710 1760.260 2794.275 ;
        RECT 1766.490 2793.595 1766.770 2793.965 ;
        RECT 1780.290 2793.595 1780.570 2793.965 ;
        RECT 1766.500 2793.450 1766.760 2793.595 ;
        RECT 1780.360 2793.430 1780.500 2793.595 ;
        RECT 1780.300 2793.110 1780.560 2793.430 ;
        RECT 1787.190 2792.915 1787.470 2793.285 ;
        RECT 1787.200 2792.770 1787.460 2792.915 ;
        RECT 1773.390 2791.555 1773.670 2791.925 ;
        RECT 1794.090 2791.555 1794.370 2791.925 ;
        RECT 1773.460 2791.390 1773.600 2791.555 ;
        RECT 1794.100 2791.410 1794.360 2791.555 ;
        RECT 2090.800 2791.410 2091.060 2791.730 ;
        RECT 1773.400 2791.070 1773.660 2791.390 ;
        RECT 1797.320 2790.730 1797.580 2791.050 ;
        RECT 1760.060 2790.390 1760.320 2790.710 ;
        RECT 1783.520 2790.390 1783.780 2790.710 ;
        RECT 1741.200 2790.050 1741.460 2790.370 ;
        RECT 1690.600 2789.370 1690.860 2789.690 ;
        RECT 1762.820 2789.370 1763.080 2789.690 ;
        RECT 1683.690 2788.155 1683.970 2788.525 ;
        RECT 1718.190 2788.155 1718.470 2788.525 ;
        RECT 1760.510 2788.155 1760.790 2788.525 ;
        RECT 1656.090 2787.475 1656.370 2787.845 ;
        RECT 1662.990 2787.475 1663.270 2787.845 ;
        RECT 1669.890 2787.475 1670.170 2787.845 ;
        RECT 1676.790 2787.475 1677.070 2787.845 ;
        RECT 1677.260 2787.670 1677.520 2787.990 ;
        RECT 1656.160 2079.770 1656.300 2787.475 ;
        RECT 1663.060 2080.110 1663.200 2787.475 ;
        RECT 1663.000 2079.790 1663.260 2080.110 ;
        RECT 1656.100 2079.450 1656.360 2079.770 ;
        RECT 1649.660 2071.970 1649.920 2072.290 ;
        RECT 1669.960 2065.830 1670.100 2787.475 ;
        RECT 1676.860 2066.170 1677.000 2787.475 ;
        RECT 1683.760 2068.890 1683.900 2788.155 ;
        RECT 1684.150 2787.475 1684.430 2787.845 ;
        RECT 1690.590 2787.475 1690.870 2787.845 ;
        RECT 1697.490 2787.475 1697.770 2787.845 ;
        RECT 1704.390 2787.475 1704.670 2787.845 ;
        RECT 1711.290 2787.475 1711.570 2787.845 ;
        RECT 1684.220 2069.570 1684.360 2787.475 ;
        RECT 1684.160 2069.250 1684.420 2069.570 ;
        RECT 1683.700 2068.570 1683.960 2068.890 ;
        RECT 1690.660 2068.550 1690.800 2787.475 ;
        RECT 1697.560 2069.230 1697.700 2787.475 ;
        RECT 1697.500 2068.910 1697.760 2069.230 ;
        RECT 1690.600 2068.230 1690.860 2068.550 ;
        RECT 1704.460 2067.530 1704.600 2787.475 ;
        RECT 1711.360 2068.210 1711.500 2787.475 ;
        RECT 1711.300 2067.890 1711.560 2068.210 ;
        RECT 1718.260 2067.870 1718.400 2788.155 ;
        RECT 1718.650 2787.475 1718.930 2787.845 ;
        RECT 1725.090 2787.475 1725.370 2787.845 ;
        RECT 1731.990 2787.475 1732.270 2787.845 ;
        RECT 1738.890 2787.475 1739.170 2787.845 ;
        RECT 1745.790 2787.475 1746.070 2787.845 ;
        RECT 1752.690 2787.475 1752.970 2787.845 ;
        RECT 1760.050 2787.475 1760.330 2787.845 ;
        RECT 1718.200 2067.550 1718.460 2067.870 ;
        RECT 1704.400 2067.210 1704.660 2067.530 ;
        RECT 1718.720 2066.510 1718.860 2787.475 ;
        RECT 1725.160 2067.190 1725.300 2787.475 ;
        RECT 1725.100 2066.870 1725.360 2067.190 ;
        RECT 1732.060 2066.850 1732.200 2787.475 ;
        RECT 1738.960 2073.310 1739.100 2787.475 ;
        RECT 1745.860 2076.370 1746.000 2787.475 ;
        RECT 1745.800 2076.050 1746.060 2076.370 ;
        RECT 1752.760 2075.690 1752.900 2787.475 ;
        RECT 1752.700 2075.370 1752.960 2075.690 ;
        RECT 1760.120 2074.670 1760.260 2787.475 ;
        RECT 1760.580 2076.030 1760.720 2788.155 ;
        RECT 1762.880 2097.110 1763.020 2789.370 ;
        RECT 1766.490 2787.475 1766.770 2787.845 ;
        RECT 1773.850 2787.475 1774.130 2787.845 ;
        RECT 1780.290 2787.475 1780.570 2787.845 ;
        RECT 1762.820 2096.790 1763.080 2097.110 ;
        RECT 1760.520 2075.710 1760.780 2076.030 ;
        RECT 1766.560 2075.350 1766.700 2787.475 ;
        RECT 1766.500 2075.030 1766.760 2075.350 ;
        RECT 1773.920 2075.010 1774.060 2787.475 ;
        RECT 1773.860 2074.690 1774.120 2075.010 ;
        RECT 1760.060 2074.350 1760.320 2074.670 ;
        RECT 1780.360 2074.330 1780.500 2787.475 ;
        RECT 1783.580 2090.650 1783.720 2790.390 ;
        RECT 1790.420 2790.050 1790.680 2790.370 ;
        RECT 1787.190 2787.475 1787.470 2787.845 ;
        RECT 1783.520 2090.330 1783.780 2090.650 ;
        RECT 1780.300 2074.010 1780.560 2074.330 ;
        RECT 1787.260 2073.990 1787.400 2787.475 ;
        RECT 1790.480 2097.450 1790.620 2790.050 ;
        RECT 1794.550 2787.475 1794.830 2787.845 ;
        RECT 1790.420 2097.130 1790.680 2097.450 ;
        RECT 1787.200 2073.670 1787.460 2073.990 ;
        RECT 1794.620 2073.650 1794.760 2787.475 ;
        RECT 1797.380 2104.590 1797.520 2790.730 ;
        RECT 1797.780 2789.710 1798.040 2790.030 ;
        RECT 1797.840 2111.390 1797.980 2789.710 ;
        RECT 2090.860 2788.330 2091.000 2791.410 ;
        RECT 1828.140 2788.010 1828.400 2788.330 ;
        RECT 1869.540 2788.010 1869.800 2788.330 ;
        RECT 2090.800 2788.010 2091.060 2788.330 ;
        RECT 1828.200 2787.845 1828.340 2788.010 ;
        RECT 1869.600 2787.845 1869.740 2788.010 ;
        RECT 1828.130 2787.475 1828.410 2787.845 ;
        RECT 1869.530 2787.475 1869.810 2787.845 ;
        RECT 1797.780 2111.070 1798.040 2111.390 ;
        RECT 1797.320 2104.270 1797.580 2104.590 ;
        RECT 1794.560 2073.330 1794.820 2073.650 ;
        RECT 1738.900 2072.990 1739.160 2073.310 ;
        RECT 1732.000 2066.530 1732.260 2066.850 ;
        RECT 1718.660 2066.190 1718.920 2066.510 ;
        RECT 1676.800 2065.850 1677.060 2066.170 ;
        RECT 1669.900 2065.510 1670.160 2065.830 ;
        RECT 1614.700 2064.830 1614.960 2065.150 ;
        RECT 2190.680 2062.430 2190.820 3230.155 ;
        RECT 2191.070 3224.715 2191.350 3225.085 ;
        RECT 2190.620 2062.110 2190.880 2062.430 ;
        RECT 2191.140 2061.410 2191.280 3224.715 ;
        RECT 2191.530 3215.875 2191.810 3216.245 ;
        RECT 2191.600 2062.090 2191.740 3215.875 ;
        RECT 2191.990 3209.755 2192.270 3210.125 ;
        RECT 2191.540 2061.770 2191.800 2062.090 ;
        RECT 2192.060 2061.750 2192.200 3209.755 ;
        RECT 2192.450 3201.595 2192.730 3201.965 ;
        RECT 2192.000 2061.430 2192.260 2061.750 ;
        RECT 2191.080 2061.090 2191.340 2061.410 ;
        RECT 2192.520 2059.370 2192.660 3201.595 ;
        RECT 2192.910 3196.155 2193.190 3196.525 ;
        RECT 2192.460 2059.050 2192.720 2059.370 ;
        RECT 2192.980 2059.030 2193.120 3196.155 ;
        RECT 2193.370 3187.995 2193.650 3188.365 ;
        RECT 2193.440 2062.770 2193.580 3187.995 ;
        RECT 2193.830 2898.315 2194.110 2898.685 ;
        RECT 2193.900 2087.445 2194.040 2898.315 ;
      LAYER met2 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met2 ;
        RECT 2582.140 3249.565 2582.280 3252.110 ;
        RECT 2582.070 3249.195 2582.350 3249.565 ;
        RECT 2594.560 2946.965 2594.700 3263.670 ;
        RECT 2594.490 2946.595 2594.770 2946.965 ;
        RECT 2594.560 2938.805 2594.700 2946.595 ;
        RECT 2594.490 2938.435 2594.770 2938.805 ;
        RECT 2242.590 2794.275 2242.870 2794.645 ;
        RECT 2256.390 2794.275 2256.670 2794.645 ;
        RECT 2263.290 2794.275 2263.570 2794.645 ;
        RECT 2268.350 2794.275 2268.630 2794.645 ;
        RECT 2270.190 2794.275 2270.470 2794.645 ;
        RECT 2277.090 2794.275 2277.370 2794.645 ;
        RECT 2283.990 2794.275 2284.270 2794.645 ;
        RECT 2290.890 2794.275 2291.170 2794.645 ;
        RECT 2297.790 2794.275 2298.070 2794.645 ;
        RECT 2304.690 2794.275 2304.970 2794.645 ;
        RECT 2308.830 2794.275 2309.110 2794.645 ;
        RECT 2311.590 2794.275 2311.870 2794.645 ;
        RECT 2318.490 2794.275 2318.770 2794.645 ;
        RECT 2325.390 2794.275 2325.670 2794.645 ;
        RECT 2332.290 2794.275 2332.570 2794.645 ;
        RECT 2339.650 2794.275 2339.930 2794.645 ;
        RECT 2343.790 2794.275 2344.070 2794.645 ;
        RECT 2346.090 2794.275 2346.370 2794.645 ;
        RECT 2352.990 2794.275 2353.270 2794.645 ;
        RECT 2359.890 2794.275 2360.170 2794.645 ;
        RECT 2366.790 2794.275 2367.070 2794.645 ;
        RECT 2374.150 2794.275 2374.430 2794.645 ;
        RECT 2385.650 2794.275 2385.930 2794.645 ;
        RECT 2391.630 2794.275 2391.910 2794.645 ;
        RECT 2394.850 2794.275 2395.130 2794.645 ;
        RECT 2415.090 2794.275 2415.370 2794.645 ;
        RECT 2428.890 2794.275 2429.170 2794.645 ;
        RECT 2218.220 2789.030 2218.480 2789.350 ;
        RECT 2218.280 2117.850 2218.420 2789.030 ;
        RECT 2235.690 2788.835 2235.970 2789.205 ;
        RECT 2235.700 2788.690 2235.960 2788.835 ;
        RECT 2238.920 2788.690 2239.180 2789.010 ;
        RECT 2232.020 2788.010 2232.280 2788.330 ;
        RECT 2228.790 2787.475 2229.070 2787.845 ;
        RECT 2218.220 2117.530 2218.480 2117.850 ;
        RECT 2193.830 2087.075 2194.110 2087.445 ;
        RECT 2193.380 2062.450 2193.640 2062.770 ;
        RECT 2228.860 2061.070 2229.000 2787.475 ;
        RECT 2232.080 2118.190 2232.220 2788.010 ;
        RECT 2238.980 2125.330 2239.120 2788.690 ;
        RECT 2238.920 2125.010 2239.180 2125.330 ;
        RECT 2232.020 2117.870 2232.280 2118.190 ;
        RECT 2228.800 2060.750 2229.060 2061.070 ;
        RECT 2242.660 2060.390 2242.800 2794.275 ;
        RECT 2245.820 2793.450 2246.080 2793.770 ;
        RECT 2245.880 2132.130 2246.020 2793.450 ;
        RECT 2252.720 2787.670 2252.980 2787.990 ;
        RECT 2252.780 2138.590 2252.920 2787.670 ;
        RECT 2252.720 2138.270 2252.980 2138.590 ;
        RECT 2245.820 2131.810 2246.080 2132.130 ;
        RECT 2256.460 2060.730 2256.600 2794.275 ;
        RECT 2263.360 2083.510 2263.500 2794.275 ;
        RECT 2263.750 2793.595 2264.030 2793.965 ;
        RECT 2263.300 2083.190 2263.560 2083.510 ;
        RECT 2263.820 2083.170 2263.960 2793.595 ;
        RECT 2266.510 2792.915 2266.790 2793.285 ;
        RECT 2266.580 2792.410 2266.720 2792.915 ;
        RECT 2268.420 2792.750 2268.560 2794.275 ;
        RECT 2268.360 2792.430 2268.620 2792.750 ;
        RECT 2266.520 2792.090 2266.780 2792.410 ;
        RECT 2263.760 2082.850 2264.020 2083.170 ;
        RECT 2266.580 2082.830 2266.720 2792.090 ;
        RECT 2266.980 2791.070 2267.240 2791.390 ;
        RECT 2267.040 2138.930 2267.180 2791.070 ;
        RECT 2266.980 2138.610 2267.240 2138.930 ;
        RECT 2266.520 2082.510 2266.780 2082.830 ;
        RECT 2270.260 2082.490 2270.400 2794.275 ;
        RECT 2273.410 2793.595 2273.690 2793.965 ;
        RECT 2273.480 2793.090 2273.620 2793.595 ;
        RECT 2273.420 2792.770 2273.680 2793.090 ;
        RECT 2270.200 2082.170 2270.460 2082.490 ;
        RECT 2256.400 2060.410 2256.660 2060.730 ;
        RECT 2242.600 2060.070 2242.860 2060.390 ;
        RECT 2192.920 2058.710 2193.180 2059.030 ;
        RECT 1601.360 2058.370 1601.620 2058.690 ;
        RECT 1580.200 2058.030 1580.460 2058.350 ;
        RECT 2273.480 2054.610 2273.620 2792.770 ;
        RECT 2273.420 2054.290 2273.680 2054.610 ;
        RECT 2277.160 2054.270 2277.300 2794.275 ;
        RECT 2279.850 2793.595 2280.130 2793.965 ;
        RECT 2279.920 2791.730 2280.060 2793.595 ;
        RECT 2279.860 2791.410 2280.120 2791.730 ;
        RECT 2277.100 2053.950 2277.360 2054.270 ;
        RECT 2284.060 2053.930 2284.200 2794.275 ;
        RECT 2284.460 2793.965 2284.720 2794.110 ;
        RECT 2284.450 2793.595 2284.730 2793.965 ;
        RECT 2284.520 2792.410 2284.660 2793.595 ;
        RECT 2284.460 2792.090 2284.720 2792.410 ;
        RECT 2284.000 2053.610 2284.260 2053.930 ;
        RECT 2290.960 2053.590 2291.100 2794.275 ;
        RECT 2294.110 2792.915 2294.390 2793.285 ;
        RECT 2294.180 2788.330 2294.320 2792.915 ;
        RECT 2294.120 2788.010 2294.380 2788.330 ;
        RECT 2294.180 2059.710 2294.320 2788.010 ;
        RECT 2297.860 2081.810 2298.000 2794.275 ;
        RECT 2298.250 2793.595 2298.530 2793.965 ;
        RECT 2301.020 2793.790 2301.280 2794.110 ;
        RECT 2304.240 2793.965 2304.500 2794.110 ;
        RECT 2298.320 2793.430 2298.460 2793.595 ;
        RECT 2298.260 2793.110 2298.520 2793.430 ;
        RECT 2297.800 2081.490 2298.060 2081.810 ;
        RECT 2301.080 2060.050 2301.220 2793.790 ;
        RECT 2304.230 2793.595 2304.510 2793.965 ;
        RECT 2301.480 2791.410 2301.740 2791.730 ;
        RECT 2301.540 2145.730 2301.680 2791.410 ;
        RECT 2301.480 2145.410 2301.740 2145.730 ;
        RECT 2301.020 2059.730 2301.280 2060.050 ;
        RECT 2294.120 2059.390 2294.380 2059.710 ;
        RECT 2290.900 2053.270 2291.160 2053.590 ;
        RECT 2304.760 2053.250 2304.900 2794.275 ;
        RECT 2305.150 2793.595 2305.430 2793.965 ;
        RECT 2308.900 2793.770 2309.040 2794.275 ;
        RECT 2305.220 2082.150 2305.360 2793.595 ;
        RECT 2308.840 2793.450 2309.100 2793.770 ;
        RECT 2307.910 2790.875 2308.190 2791.245 ;
        RECT 2307.980 2152.870 2308.120 2790.875 ;
        RECT 2307.920 2152.550 2308.180 2152.870 ;
        RECT 2305.160 2081.830 2305.420 2082.150 ;
        RECT 2304.700 2052.930 2304.960 2053.250 ;
        RECT 2311.660 2052.910 2311.800 2794.275 ;
        RECT 2315.270 2793.595 2315.550 2793.965 ;
        RECT 2315.340 2792.750 2315.480 2793.595 ;
        RECT 2315.280 2792.430 2315.540 2792.750 ;
        RECT 2318.560 2081.470 2318.700 2794.275 ;
        RECT 2321.710 2793.595 2321.990 2793.965 ;
        RECT 2321.780 2793.090 2321.920 2793.595 ;
        RECT 2321.720 2792.770 2321.980 2793.090 ;
        RECT 2318.500 2081.150 2318.760 2081.470 ;
        RECT 2325.460 2081.130 2325.600 2794.275 ;
        RECT 2326.770 2793.595 2327.050 2793.965 ;
        RECT 2326.840 2792.070 2326.980 2793.595 ;
        RECT 2326.780 2791.750 2327.040 2792.070 ;
        RECT 2325.400 2080.810 2325.660 2081.130 ;
        RECT 2332.360 2080.790 2332.500 2794.275 ;
        RECT 2333.670 2793.595 2333.950 2793.965 ;
        RECT 2339.190 2793.595 2339.470 2793.965 ;
        RECT 2333.740 2792.410 2333.880 2793.595 ;
        RECT 2333.680 2792.090 2333.940 2792.410 ;
        RECT 2333.740 2788.330 2333.880 2792.090 ;
        RECT 2333.680 2788.010 2333.940 2788.330 ;
        RECT 2332.300 2080.470 2332.560 2080.790 ;
        RECT 2339.260 2063.110 2339.400 2793.595 ;
        RECT 2339.720 2080.450 2339.860 2794.275 ;
        RECT 2343.860 2793.430 2344.000 2794.275 ;
        RECT 2340.110 2792.915 2340.390 2793.285 ;
        RECT 2343.800 2793.110 2344.060 2793.430 ;
        RECT 2340.180 2792.410 2340.320 2792.915 ;
        RECT 2340.120 2792.090 2340.380 2792.410 ;
        RECT 2339.660 2080.130 2339.920 2080.450 ;
        RECT 2346.160 2069.910 2346.300 2794.275 ;
        RECT 2347.480 2793.965 2347.740 2794.110 ;
        RECT 2347.470 2793.595 2347.750 2793.965 ;
        RECT 2347.540 2792.410 2347.680 2793.595 ;
        RECT 2347.480 2792.090 2347.740 2792.410 ;
        RECT 2353.060 2076.710 2353.200 2794.275 ;
        RECT 2356.670 2793.595 2356.950 2793.965 ;
        RECT 2356.680 2793.450 2356.940 2793.595 ;
        RECT 2359.960 2077.050 2360.100 2794.275 ;
        RECT 2361.270 2793.595 2361.550 2793.965 ;
        RECT 2361.340 2792.750 2361.480 2793.595 ;
        RECT 2361.280 2792.430 2361.540 2792.750 ;
        RECT 2366.860 2083.850 2367.000 2794.275 ;
        RECT 2367.250 2793.595 2367.530 2793.965 ;
        RECT 2367.320 2793.090 2367.460 2793.595 ;
        RECT 2367.260 2792.770 2367.520 2793.090 ;
        RECT 2373.690 2792.915 2373.970 2793.285 ;
        RECT 2373.760 2790.710 2373.900 2792.915 ;
        RECT 2374.220 2792.070 2374.360 2794.275 ;
        RECT 2385.720 2794.110 2385.860 2794.275 ;
        RECT 2377.370 2793.595 2377.650 2793.965 ;
        RECT 2385.660 2793.790 2385.920 2794.110 ;
        RECT 2374.160 2791.750 2374.420 2792.070 ;
        RECT 2377.440 2790.710 2377.580 2793.595 ;
        RECT 2391.700 2793.430 2391.840 2794.275 ;
        RECT 2391.640 2793.110 2391.900 2793.430 ;
        RECT 2394.920 2792.410 2395.060 2794.275 ;
        RECT 2415.100 2794.130 2415.360 2794.275 ;
        RECT 2428.960 2794.110 2429.100 2794.275 ;
        RECT 2402.670 2793.595 2402.950 2793.965 ;
        RECT 2421.990 2793.595 2422.270 2793.965 ;
        RECT 2428.900 2793.790 2429.160 2794.110 ;
        RECT 2435.790 2793.595 2436.070 2793.965 ;
        RECT 2402.680 2793.450 2402.940 2793.595 ;
        RECT 2402.670 2792.915 2402.950 2793.285 ;
        RECT 2408.190 2792.915 2408.470 2793.285 ;
        RECT 2415.090 2792.915 2415.370 2793.285 ;
        RECT 2394.860 2792.090 2395.120 2792.410 ;
        RECT 2387.490 2791.555 2387.770 2791.925 ;
        RECT 2387.560 2791.050 2387.700 2791.555 ;
        RECT 2394.920 2791.050 2395.060 2792.090 ;
        RECT 2387.500 2790.730 2387.760 2791.050 ;
        RECT 2394.860 2790.730 2395.120 2791.050 ;
        RECT 2373.700 2790.390 2373.960 2790.710 ;
        RECT 2377.380 2790.390 2377.640 2790.710 ;
        RECT 2377.440 2788.330 2377.580 2790.390 ;
        RECT 2380.590 2790.195 2380.870 2790.565 ;
        RECT 2394.390 2790.195 2394.670 2790.565 ;
        RECT 2380.600 2790.050 2380.860 2790.195 ;
        RECT 2394.460 2790.030 2394.600 2790.195 ;
        RECT 2380.590 2789.515 2380.870 2789.885 ;
        RECT 2394.400 2789.710 2394.660 2790.030 ;
        RECT 2380.600 2789.370 2380.860 2789.515 ;
        RECT 2402.740 2789.350 2402.880 2792.915 ;
        RECT 2408.260 2792.750 2408.400 2792.915 ;
        RECT 2415.100 2792.770 2415.360 2792.915 ;
        RECT 2408.200 2792.430 2408.460 2792.750 ;
        RECT 2415.090 2792.235 2415.370 2792.605 ;
        RECT 2415.160 2792.070 2415.300 2792.235 ;
        RECT 2415.100 2791.750 2415.360 2792.070 ;
        RECT 2408.190 2790.875 2408.470 2791.245 ;
        RECT 2402.680 2789.030 2402.940 2789.350 ;
        RECT 2408.260 2789.010 2408.400 2790.875 ;
        RECT 2422.060 2790.710 2422.200 2793.595 ;
        RECT 2435.860 2793.430 2436.000 2793.595 ;
        RECT 2435.800 2793.110 2436.060 2793.430 ;
        RECT 2442.690 2792.915 2442.970 2793.285 ;
        RECT 2428.890 2791.555 2429.170 2791.925 ;
        RECT 2435.790 2791.555 2436.070 2791.925 ;
        RECT 2428.960 2791.390 2429.100 2791.555 ;
        RECT 2435.800 2791.410 2436.060 2791.555 ;
        RECT 2428.900 2791.070 2429.160 2791.390 ;
        RECT 2442.760 2791.050 2442.900 2792.915 ;
        RECT 2442.700 2790.730 2442.960 2791.050 ;
        RECT 2422.000 2790.390 2422.260 2790.710 ;
        RECT 2408.200 2788.690 2408.460 2789.010 ;
        RECT 2415.090 2788.835 2415.370 2789.205 ;
        RECT 2415.160 2788.670 2415.300 2788.835 ;
        RECT 2415.100 2788.350 2415.360 2788.670 ;
        RECT 2377.380 2788.010 2377.640 2788.330 ;
        RECT 2421.990 2788.155 2422.270 2788.525 ;
        RECT 2422.060 2787.990 2422.200 2788.155 ;
        RECT 2422.000 2787.670 2422.260 2787.990 ;
        RECT 2366.800 2083.530 2367.060 2083.850 ;
        RECT 2359.900 2076.730 2360.160 2077.050 ;
        RECT 2353.000 2076.390 2353.260 2076.710 ;
        RECT 2346.100 2069.590 2346.360 2069.910 ;
        RECT 2339.200 2062.790 2339.460 2063.110 ;
        RECT 2311.600 2052.590 2311.860 2052.910 ;
        RECT 1549.840 1855.730 1550.100 1856.050 ;
        RECT 1549.380 1855.390 1549.640 1855.710 ;
        RECT 1548.920 1848.930 1549.180 1849.250 ;
        RECT 1494.180 1807.450 1494.440 1807.770 ;
        RECT 1493.720 1710.890 1493.980 1711.210 ;
        RECT 1460.140 1655.810 1460.400 1656.130 ;
        RECT 1426.100 1635.070 1426.360 1635.390 ;
        RECT 1412.290 1621.955 1412.570 1622.325 ;
        RECT 1410.910 1617.195 1411.190 1617.565 ;
        RECT 1408.150 1611.755 1408.430 1612.125 ;
        RECT 1407.690 1606.995 1407.970 1607.365 ;
      LAYER met2 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
      LAYER met2 ;
        RECT 1397.570 1603.595 1397.850 1603.965 ;
      LAYER met2 ;
        RECT 1550.030 1495.720 1554.800 1497.365 ;
      LAYER met2 ;
        RECT 1555.080 1496.000 1555.360 1500.000 ;
      LAYER met2 ;
        RECT 1555.640 1495.720 1564.920 1497.365 ;
      LAYER met2 ;
        RECT 1565.200 1496.000 1565.480 1500.000 ;
      LAYER met2 ;
        RECT 1565.760 1495.720 1575.500 1497.365 ;
      LAYER met2 ;
        RECT 1575.780 1496.000 1576.060 1500.000 ;
      LAYER met2 ;
        RECT 1576.340 1495.720 1585.620 1497.365 ;
      LAYER met2 ;
        RECT 1585.900 1496.000 1586.180 1500.000 ;
      LAYER met2 ;
        RECT 1586.460 1495.720 1596.200 1497.365 ;
      LAYER met2 ;
        RECT 1596.480 1496.000 1596.760 1500.000 ;
      LAYER met2 ;
        RECT 1597.040 1495.720 1606.320 1497.365 ;
      LAYER met2 ;
        RECT 1606.600 1496.000 1606.880 1500.000 ;
      LAYER met2 ;
        RECT 1607.160 1495.720 1616.900 1497.365 ;
      LAYER met2 ;
        RECT 1617.180 1496.000 1617.460 1500.000 ;
      LAYER met2 ;
        RECT 1617.740 1495.720 1627.020 1497.365 ;
      LAYER met2 ;
        RECT 1627.300 1496.000 1627.580 1500.000 ;
      LAYER met2 ;
        RECT 1627.860 1495.720 1637.600 1497.365 ;
      LAYER met2 ;
        RECT 1637.880 1496.000 1638.160 1500.000 ;
      LAYER met2 ;
        RECT 1638.440 1495.720 1648.180 1497.365 ;
      LAYER met2 ;
        RECT 1648.460 1496.000 1648.740 1500.000 ;
      LAYER met2 ;
        RECT 1649.020 1495.720 1658.300 1497.365 ;
      LAYER met2 ;
        RECT 1658.580 1496.000 1658.860 1500.000 ;
      LAYER met2 ;
        RECT 1659.140 1495.720 1668.880 1497.365 ;
      LAYER met2 ;
        RECT 1669.160 1496.000 1669.440 1500.000 ;
      LAYER met2 ;
        RECT 1669.720 1495.720 1679.000 1497.365 ;
      LAYER met2 ;
        RECT 1679.280 1496.000 1679.560 1500.000 ;
      LAYER met2 ;
        RECT 1679.840 1495.720 1689.580 1497.365 ;
      LAYER met2 ;
        RECT 1689.860 1496.000 1690.140 1500.000 ;
      LAYER met2 ;
        RECT 1690.420 1495.720 1699.700 1497.365 ;
      LAYER met2 ;
        RECT 1699.980 1496.000 1700.260 1500.000 ;
      LAYER met2 ;
        RECT 1700.540 1495.720 1710.280 1497.365 ;
      LAYER met2 ;
        RECT 1710.560 1496.000 1710.840 1500.000 ;
      LAYER met2 ;
        RECT 1711.120 1495.720 1720.400 1497.365 ;
      LAYER met2 ;
        RECT 1720.680 1496.000 1720.960 1500.000 ;
      LAYER met2 ;
        RECT 1721.240 1495.720 1730.980 1497.365 ;
      LAYER met2 ;
        RECT 1731.260 1496.000 1731.540 1500.000 ;
      LAYER met2 ;
        RECT 1731.820 1495.720 1741.560 1497.365 ;
      LAYER met2 ;
        RECT 1741.840 1496.000 1742.120 1500.000 ;
      LAYER met2 ;
        RECT 1742.400 1495.720 1751.680 1497.365 ;
      LAYER met2 ;
        RECT 1751.960 1496.000 1752.240 1500.000 ;
      LAYER met2 ;
        RECT 1752.520 1495.720 1762.260 1497.365 ;
      LAYER met2 ;
        RECT 1762.540 1496.000 1762.820 1500.000 ;
      LAYER met2 ;
        RECT 1763.100 1495.720 1772.380 1497.365 ;
      LAYER met2 ;
        RECT 1772.660 1496.000 1772.940 1500.000 ;
      LAYER met2 ;
        RECT 1773.220 1495.720 1782.960 1497.365 ;
      LAYER met2 ;
        RECT 1783.240 1496.000 1783.520 1500.000 ;
      LAYER met2 ;
        RECT 1783.800 1495.720 1793.080 1497.365 ;
      LAYER met2 ;
        RECT 1793.360 1496.000 1793.640 1500.000 ;
      LAYER met2 ;
        RECT 1793.920 1495.720 1803.660 1497.365 ;
      LAYER met2 ;
        RECT 1803.940 1496.000 1804.220 1500.000 ;
      LAYER met2 ;
        RECT 1804.500 1495.720 1813.780 1497.365 ;
      LAYER met2 ;
        RECT 1814.060 1496.000 1814.340 1500.000 ;
      LAYER met2 ;
        RECT 1814.620 1495.720 1824.360 1497.365 ;
      LAYER met2 ;
        RECT 1824.640 1496.000 1824.920 1500.000 ;
      LAYER met2 ;
        RECT 1825.200 1495.720 1834.940 1497.365 ;
      LAYER met2 ;
        RECT 1835.220 1496.000 1835.500 1500.000 ;
      LAYER met2 ;
        RECT 1835.780 1495.720 1845.060 1497.365 ;
      LAYER met2 ;
        RECT 1845.340 1496.000 1845.620 1500.000 ;
      LAYER met2 ;
        RECT 1845.900 1495.720 1855.640 1497.365 ;
      LAYER met2 ;
        RECT 1855.920 1496.000 1856.200 1500.000 ;
      LAYER met2 ;
        RECT 1856.480 1495.720 1865.760 1497.365 ;
      LAYER met2 ;
        RECT 1866.040 1496.000 1866.320 1500.000 ;
      LAYER met2 ;
        RECT 1866.600 1495.720 1876.340 1497.365 ;
      LAYER met2 ;
        RECT 1876.620 1496.000 1876.900 1500.000 ;
      LAYER met2 ;
        RECT 1877.180 1495.720 1886.460 1497.365 ;
      LAYER met2 ;
        RECT 1886.740 1496.000 1887.020 1500.000 ;
      LAYER met2 ;
        RECT 1887.300 1495.720 1897.040 1497.365 ;
      LAYER met2 ;
        RECT 1897.320 1496.000 1897.600 1500.000 ;
      LAYER met2 ;
        RECT 1897.880 1495.720 1907.160 1497.365 ;
      LAYER met2 ;
        RECT 1907.440 1496.000 1907.720 1500.000 ;
      LAYER met2 ;
        RECT 1908.000 1495.720 1917.740 1497.365 ;
      LAYER met2 ;
        RECT 1918.020 1496.000 1918.300 1500.000 ;
      LAYER met2 ;
        RECT 1918.580 1495.720 1928.320 1497.365 ;
      LAYER met2 ;
        RECT 1928.600 1496.000 1928.880 1500.000 ;
      LAYER met2 ;
        RECT 1929.160 1495.720 1938.440 1497.365 ;
      LAYER met2 ;
        RECT 1938.720 1496.000 1939.000 1500.000 ;
      LAYER met2 ;
        RECT 1939.280 1495.720 1949.020 1497.365 ;
      LAYER met2 ;
        RECT 1949.300 1496.000 1949.580 1500.000 ;
      LAYER met2 ;
        RECT 1949.860 1495.720 1959.140 1497.365 ;
      LAYER met2 ;
        RECT 1959.420 1496.000 1959.700 1500.000 ;
      LAYER met2 ;
        RECT 1959.980 1495.720 1969.720 1497.365 ;
      LAYER met2 ;
        RECT 1970.000 1496.000 1970.280 1500.000 ;
      LAYER met2 ;
        RECT 1970.560 1495.720 1979.840 1497.365 ;
      LAYER met2 ;
        RECT 1980.120 1496.000 1980.400 1500.000 ;
      LAYER met2 ;
        RECT 1980.680 1495.720 1990.420 1497.365 ;
      LAYER met2 ;
        RECT 1990.700 1496.000 1990.980 1500.000 ;
      LAYER met2 ;
        RECT 1991.260 1495.720 2000.540 1497.365 ;
      LAYER met2 ;
        RECT 2000.820 1496.000 2001.100 1500.000 ;
      LAYER met2 ;
        RECT 2001.380 1495.720 2011.120 1497.365 ;
      LAYER met2 ;
        RECT 2011.400 1496.000 2011.680 1500.000 ;
      LAYER met2 ;
        RECT 2011.960 1495.720 2021.700 1497.365 ;
      LAYER met2 ;
        RECT 2021.980 1496.000 2022.260 1500.000 ;
      LAYER met2 ;
        RECT 2022.540 1495.720 2031.820 1497.365 ;
      LAYER met2 ;
        RECT 2032.100 1496.000 2032.380 1500.000 ;
      LAYER met2 ;
        RECT 2032.660 1495.720 2042.400 1497.365 ;
      LAYER met2 ;
        RECT 2042.680 1496.000 2042.960 1500.000 ;
      LAYER met2 ;
        RECT 2043.240 1495.720 2052.520 1497.365 ;
      LAYER met2 ;
        RECT 2052.800 1496.000 2053.080 1500.000 ;
      LAYER met2 ;
        RECT 2053.360 1495.720 2063.100 1497.365 ;
      LAYER met2 ;
        RECT 2063.380 1496.000 2063.660 1500.000 ;
      LAYER met2 ;
        RECT 2063.940 1495.720 2073.220 1497.365 ;
      LAYER met2 ;
        RECT 2073.500 1496.000 2073.780 1500.000 ;
      LAYER met2 ;
        RECT 2074.060 1495.720 2083.800 1497.365 ;
      LAYER met2 ;
        RECT 2084.080 1496.000 2084.360 1500.000 ;
      LAYER met2 ;
        RECT 2084.640 1495.720 2093.920 1497.365 ;
      LAYER met2 ;
        RECT 2094.200 1496.000 2094.480 1500.000 ;
      LAYER met2 ;
        RECT 2094.760 1495.720 2104.500 1497.365 ;
      LAYER met2 ;
        RECT 2104.780 1496.000 2105.060 1500.000 ;
      LAYER met2 ;
        RECT 2105.340 1495.720 2115.080 1497.365 ;
      LAYER met2 ;
        RECT 2115.360 1496.000 2115.640 1500.000 ;
      LAYER met2 ;
        RECT 2115.920 1495.720 2125.200 1497.365 ;
      LAYER met2 ;
        RECT 2125.480 1496.000 2125.760 1500.000 ;
      LAYER met2 ;
        RECT 2126.040 1495.720 2135.780 1497.365 ;
      LAYER met2 ;
        RECT 2136.060 1496.000 2136.340 1500.000 ;
      LAYER met2 ;
        RECT 2136.620 1495.720 2145.900 1497.365 ;
      LAYER met2 ;
        RECT 2146.180 1496.000 2146.460 1500.000 ;
      LAYER met2 ;
        RECT 2146.740 1495.720 2156.480 1497.365 ;
      LAYER met2 ;
        RECT 2156.760 1496.000 2157.040 1500.000 ;
      LAYER met2 ;
        RECT 2157.320 1495.720 2166.600 1497.365 ;
      LAYER met2 ;
        RECT 2166.880 1496.000 2167.160 1500.000 ;
      LAYER met2 ;
        RECT 2167.440 1495.720 2177.180 1497.365 ;
      LAYER met2 ;
        RECT 2177.460 1496.000 2177.740 1500.000 ;
      LAYER met2 ;
        RECT 2178.020 1495.720 2187.300 1497.365 ;
      LAYER met2 ;
        RECT 2187.580 1496.000 2187.860 1500.000 ;
      LAYER met2 ;
        RECT 2188.140 1495.720 2197.880 1497.365 ;
      LAYER met2 ;
        RECT 2198.160 1496.000 2198.440 1500.000 ;
      LAYER met2 ;
        RECT 2198.720 1495.720 2208.460 1497.365 ;
      LAYER met2 ;
        RECT 2208.740 1496.000 2209.020 1500.000 ;
      LAYER met2 ;
        RECT 2209.300 1495.720 2218.580 1497.365 ;
      LAYER met2 ;
        RECT 2218.860 1496.000 2219.140 1500.000 ;
      LAYER met2 ;
        RECT 2219.420 1495.720 2229.160 1497.365 ;
      LAYER met2 ;
        RECT 2229.440 1496.000 2229.720 1500.000 ;
      LAYER met2 ;
        RECT 2230.000 1495.720 2239.280 1497.365 ;
      LAYER met2 ;
        RECT 2239.560 1496.000 2239.840 1500.000 ;
      LAYER met2 ;
        RECT 2240.120 1495.720 2249.860 1497.365 ;
      LAYER met2 ;
        RECT 2250.140 1496.000 2250.420 1500.000 ;
      LAYER met2 ;
        RECT 2250.700 1495.720 2259.980 1497.365 ;
      LAYER met2 ;
        RECT 2260.260 1496.000 2260.540 1500.000 ;
      LAYER met2 ;
        RECT 2260.820 1495.720 2270.560 1497.365 ;
      LAYER met2 ;
        RECT 2270.840 1496.000 2271.120 1500.000 ;
      LAYER met2 ;
        RECT 2271.400 1495.720 2280.680 1497.365 ;
      LAYER met2 ;
        RECT 2280.960 1496.000 2281.240 1500.000 ;
      LAYER met2 ;
        RECT 2281.520 1495.720 2291.260 1497.365 ;
      LAYER met2 ;
        RECT 2291.540 1496.000 2291.820 1500.000 ;
      LAYER met2 ;
        RECT 2292.100 1495.720 2301.840 1497.365 ;
      LAYER met2 ;
        RECT 2302.120 1496.000 2302.400 1500.000 ;
      LAYER met2 ;
        RECT 2302.680 1495.720 2311.960 1497.365 ;
      LAYER met2 ;
        RECT 2312.240 1496.000 2312.520 1500.000 ;
      LAYER met2 ;
        RECT 2312.800 1495.720 2322.540 1497.365 ;
      LAYER met2 ;
        RECT 2322.820 1496.000 2323.100 1500.000 ;
      LAYER met2 ;
        RECT 2323.380 1495.720 2332.660 1497.365 ;
      LAYER met2 ;
        RECT 2332.940 1496.000 2333.220 1500.000 ;
      LAYER met2 ;
        RECT 2333.500 1495.720 2343.240 1497.365 ;
      LAYER met2 ;
        RECT 2343.520 1496.000 2343.800 1500.000 ;
      LAYER met2 ;
        RECT 2344.080 1495.720 2353.360 1497.365 ;
      LAYER met2 ;
        RECT 2353.640 1496.000 2353.920 1500.000 ;
      LAYER met2 ;
        RECT 2354.200 1495.720 2363.940 1497.365 ;
      LAYER met2 ;
        RECT 2364.220 1496.000 2364.500 1500.000 ;
      LAYER met2 ;
        RECT 2364.780 1495.720 2374.060 1497.365 ;
      LAYER met2 ;
        RECT 2374.340 1496.000 2374.620 1500.000 ;
      LAYER met2 ;
        RECT 2374.900 1495.720 2384.640 1497.365 ;
      LAYER met2 ;
        RECT 2384.920 1496.000 2385.200 1500.000 ;
      LAYER met2 ;
        RECT 2385.480 1495.720 2395.220 1497.365 ;
      LAYER met2 ;
        RECT 2395.500 1496.000 2395.780 1500.000 ;
      LAYER met2 ;
        RECT 2396.060 1495.720 2405.340 1497.365 ;
      LAYER met2 ;
        RECT 2405.620 1496.000 2405.900 1500.000 ;
      LAYER met2 ;
        RECT 2406.180 1495.720 2415.920 1497.365 ;
      LAYER met2 ;
        RECT 2416.200 1496.000 2416.480 1500.000 ;
      LAYER met2 ;
        RECT 2416.760 1495.720 2426.040 1497.365 ;
      LAYER met2 ;
        RECT 2426.320 1496.000 2426.600 1500.000 ;
      LAYER met2 ;
        RECT 2426.880 1495.720 2436.620 1497.365 ;
      LAYER met2 ;
        RECT 2436.900 1496.000 2437.180 1500.000 ;
      LAYER met2 ;
        RECT 2437.460 1495.720 2446.740 1497.365 ;
      LAYER met2 ;
        RECT 2447.020 1496.000 2447.300 1500.000 ;
      LAYER met2 ;
        RECT 2447.580 1495.720 2457.320 1497.365 ;
      LAYER met2 ;
        RECT 2457.600 1496.000 2457.880 1500.000 ;
      LAYER met2 ;
        RECT 2458.160 1495.720 2467.440 1497.365 ;
      LAYER met2 ;
        RECT 2467.720 1496.000 2468.000 1500.000 ;
      LAYER met2 ;
        RECT 2468.280 1495.720 2478.020 1497.365 ;
      LAYER met2 ;
        RECT 2478.300 1496.000 2478.580 1500.000 ;
      LAYER met2 ;
        RECT 2478.860 1495.720 2488.600 1497.365 ;
      LAYER met2 ;
        RECT 2488.880 1496.000 2489.160 1500.000 ;
      LAYER met2 ;
        RECT 2489.440 1495.720 2498.720 1497.365 ;
      LAYER met2 ;
        RECT 2499.000 1496.000 2499.280 1500.000 ;
      LAYER met2 ;
        RECT 2499.560 1495.720 2509.300 1497.365 ;
      LAYER met2 ;
        RECT 2509.580 1496.000 2509.860 1500.000 ;
      LAYER met2 ;
        RECT 2510.140 1495.720 2519.420 1497.365 ;
      LAYER met2 ;
        RECT 2519.700 1496.000 2519.980 1500.000 ;
      LAYER met2 ;
        RECT 2520.260 1495.720 2530.000 1497.365 ;
      LAYER met2 ;
        RECT 2530.280 1496.000 2530.560 1500.000 ;
      LAYER met2 ;
        RECT 2530.840 1495.720 2540.120 1497.365 ;
      LAYER met2 ;
        RECT 2540.400 1496.000 2540.680 1500.000 ;
      LAYER met2 ;
        RECT 2540.960 1495.720 2550.700 1497.365 ;
      LAYER met2 ;
        RECT 2550.980 1496.000 2551.260 1500.000 ;
      LAYER met2 ;
        RECT 2551.540 1495.720 2560.820 1497.365 ;
      LAYER met2 ;
        RECT 2561.100 1496.000 2561.380 1500.000 ;
      LAYER met2 ;
        RECT 2561.660 1495.720 2571.400 1497.365 ;
      LAYER met2 ;
        RECT 2571.680 1496.000 2571.960 1500.000 ;
      LAYER met2 ;
        RECT 2572.240 1495.720 2581.980 1497.365 ;
      LAYER met2 ;
        RECT 2582.260 1496.000 2582.540 1500.000 ;
      LAYER met2 ;
        RECT 2582.820 1495.720 2592.100 1497.365 ;
      LAYER met2 ;
        RECT 2592.380 1496.000 2592.660 1500.000 ;
      LAYER met2 ;
        RECT 2592.940 1495.720 2602.680 1497.365 ;
      LAYER met2 ;
        RECT 2602.960 1496.000 2603.240 1500.000 ;
      LAYER met2 ;
        RECT 2603.520 1495.720 2612.800 1497.365 ;
      LAYER met2 ;
        RECT 2613.080 1496.000 2613.360 1500.000 ;
      LAYER met2 ;
        RECT 2613.640 1495.720 2623.380 1497.365 ;
      LAYER met2 ;
        RECT 2623.660 1496.000 2623.940 1500.000 ;
      LAYER met2 ;
        RECT 2624.220 1495.720 2633.500 1497.365 ;
      LAYER met2 ;
        RECT 2633.780 1496.000 2634.060 1500.000 ;
      LAYER met2 ;
        RECT 2634.340 1495.720 2644.080 1497.365 ;
      LAYER met2 ;
        RECT 2644.360 1496.000 2644.640 1500.000 ;
      LAYER met2 ;
        RECT 2644.920 1495.720 2647.390 1497.365 ;
        RECT 1550.030 404.280 2647.390 1495.720 ;
        RECT 1550.030 402.195 1552.040 404.280 ;
      LAYER met2 ;
        RECT 1552.320 400.000 1552.600 404.000 ;
      LAYER met2 ;
        RECT 1552.880 402.195 1556.640 404.280 ;
      LAYER met2 ;
        RECT 1556.920 400.000 1557.200 404.000 ;
      LAYER met2 ;
        RECT 1557.480 402.195 1561.700 404.280 ;
      LAYER met2 ;
        RECT 1561.980 400.000 1562.260 404.000 ;
      LAYER met2 ;
        RECT 1562.540 402.195 1566.300 404.280 ;
      LAYER met2 ;
        RECT 1566.580 400.000 1566.860 404.000 ;
      LAYER met2 ;
        RECT 1567.140 402.195 1571.360 404.280 ;
      LAYER met2 ;
        RECT 1571.640 400.000 1571.920 404.000 ;
      LAYER met2 ;
        RECT 1572.200 402.195 1575.960 404.280 ;
      LAYER met2 ;
        RECT 1576.240 400.000 1576.520 404.000 ;
      LAYER met2 ;
        RECT 1576.800 402.195 1581.020 404.280 ;
      LAYER met2 ;
        RECT 1581.300 400.000 1581.580 404.000 ;
      LAYER met2 ;
        RECT 1581.860 402.195 1585.620 404.280 ;
      LAYER met2 ;
        RECT 1585.900 400.000 1586.180 404.000 ;
      LAYER met2 ;
        RECT 1586.460 402.195 1590.680 404.280 ;
      LAYER met2 ;
        RECT 1590.960 400.000 1591.240 404.000 ;
      LAYER met2 ;
        RECT 1591.520 402.195 1595.280 404.280 ;
      LAYER met2 ;
        RECT 1595.560 400.000 1595.840 404.000 ;
      LAYER met2 ;
        RECT 1596.120 402.195 1600.340 404.280 ;
      LAYER met2 ;
        RECT 1600.620 400.000 1600.900 404.000 ;
      LAYER met2 ;
        RECT 1601.180 402.195 1604.940 404.280 ;
      LAYER met2 ;
        RECT 1605.220 400.000 1605.500 404.000 ;
      LAYER met2 ;
        RECT 1605.780 402.195 1610.000 404.280 ;
      LAYER met2 ;
        RECT 1610.280 400.000 1610.560 404.000 ;
      LAYER met2 ;
        RECT 1610.840 402.195 1614.600 404.280 ;
      LAYER met2 ;
        RECT 1614.880 400.000 1615.160 404.000 ;
      LAYER met2 ;
        RECT 1615.440 402.195 1619.660 404.280 ;
      LAYER met2 ;
        RECT 1619.940 400.000 1620.220 404.000 ;
      LAYER met2 ;
        RECT 1620.500 402.195 1624.260 404.280 ;
      LAYER met2 ;
        RECT 1624.540 400.000 1624.820 404.000 ;
      LAYER met2 ;
        RECT 1625.100 402.195 1629.320 404.280 ;
      LAYER met2 ;
        RECT 1629.600 400.000 1629.880 404.000 ;
      LAYER met2 ;
        RECT 1630.160 402.195 1634.380 404.280 ;
      LAYER met2 ;
        RECT 1634.660 400.000 1634.940 404.000 ;
      LAYER met2 ;
        RECT 1635.220 402.195 1638.980 404.280 ;
      LAYER met2 ;
        RECT 1639.260 400.000 1639.540 404.000 ;
      LAYER met2 ;
        RECT 1639.820 402.195 1644.040 404.280 ;
      LAYER met2 ;
        RECT 1644.320 400.000 1644.600 404.000 ;
      LAYER met2 ;
        RECT 1644.880 402.195 1648.640 404.280 ;
      LAYER met2 ;
        RECT 1648.920 400.000 1649.200 404.000 ;
      LAYER met2 ;
        RECT 1649.480 402.195 1653.700 404.280 ;
      LAYER met2 ;
        RECT 1653.980 400.000 1654.260 404.000 ;
      LAYER met2 ;
        RECT 1654.540 402.195 1658.300 404.280 ;
      LAYER met2 ;
        RECT 1658.580 400.000 1658.860 404.000 ;
      LAYER met2 ;
        RECT 1659.140 402.195 1663.360 404.280 ;
      LAYER met2 ;
        RECT 1663.640 400.000 1663.920 404.000 ;
      LAYER met2 ;
        RECT 1664.200 402.195 1667.960 404.280 ;
      LAYER met2 ;
        RECT 1668.240 400.000 1668.520 404.000 ;
      LAYER met2 ;
        RECT 1668.800 402.195 1673.020 404.280 ;
      LAYER met2 ;
        RECT 1673.300 400.000 1673.580 404.000 ;
      LAYER met2 ;
        RECT 1673.860 402.195 1677.620 404.280 ;
      LAYER met2 ;
        RECT 1677.900 400.000 1678.180 404.000 ;
      LAYER met2 ;
        RECT 1678.460 402.195 1682.680 404.280 ;
      LAYER met2 ;
        RECT 1682.960 400.000 1683.240 404.000 ;
      LAYER met2 ;
        RECT 1683.520 402.195 1687.280 404.280 ;
      LAYER met2 ;
        RECT 1687.560 400.000 1687.840 404.000 ;
      LAYER met2 ;
        RECT 1688.120 402.195 1692.340 404.280 ;
      LAYER met2 ;
        RECT 1692.620 400.000 1692.900 404.000 ;
      LAYER met2 ;
        RECT 1693.180 402.195 1696.940 404.280 ;
      LAYER met2 ;
        RECT 1697.220 400.000 1697.500 404.000 ;
      LAYER met2 ;
        RECT 1697.780 402.195 1702.000 404.280 ;
      LAYER met2 ;
        RECT 1702.280 400.000 1702.560 404.000 ;
      LAYER met2 ;
        RECT 1702.840 402.195 1707.060 404.280 ;
      LAYER met2 ;
        RECT 1707.340 400.000 1707.620 404.000 ;
      LAYER met2 ;
        RECT 1707.900 402.195 1711.660 404.280 ;
      LAYER met2 ;
        RECT 1711.940 400.000 1712.220 404.000 ;
      LAYER met2 ;
        RECT 1712.500 402.195 1716.720 404.280 ;
      LAYER met2 ;
        RECT 1717.000 400.000 1717.280 404.000 ;
      LAYER met2 ;
        RECT 1717.560 402.195 1721.320 404.280 ;
      LAYER met2 ;
        RECT 1721.600 400.000 1721.880 404.000 ;
      LAYER met2 ;
        RECT 1722.160 402.195 1726.380 404.280 ;
      LAYER met2 ;
        RECT 1726.660 400.000 1726.940 404.000 ;
      LAYER met2 ;
        RECT 1727.220 402.195 1730.980 404.280 ;
      LAYER met2 ;
        RECT 1731.260 400.000 1731.540 404.000 ;
      LAYER met2 ;
        RECT 1731.820 402.195 1736.040 404.280 ;
      LAYER met2 ;
        RECT 1736.320 400.000 1736.600 404.000 ;
      LAYER met2 ;
        RECT 1736.880 402.195 1740.640 404.280 ;
      LAYER met2 ;
        RECT 1740.920 400.000 1741.200 404.000 ;
      LAYER met2 ;
        RECT 1741.480 402.195 1745.700 404.280 ;
      LAYER met2 ;
        RECT 1745.980 400.000 1746.260 404.000 ;
      LAYER met2 ;
        RECT 1746.540 402.195 1750.300 404.280 ;
      LAYER met2 ;
        RECT 1750.580 400.000 1750.860 404.000 ;
      LAYER met2 ;
        RECT 1751.140 402.195 1755.360 404.280 ;
      LAYER met2 ;
        RECT 1755.640 400.000 1755.920 404.000 ;
      LAYER met2 ;
        RECT 1756.200 402.195 1759.960 404.280 ;
      LAYER met2 ;
        RECT 1760.240 400.000 1760.520 404.000 ;
      LAYER met2 ;
        RECT 1760.800 402.195 1765.020 404.280 ;
      LAYER met2 ;
        RECT 1765.300 400.000 1765.580 404.000 ;
      LAYER met2 ;
        RECT 1765.860 402.195 1769.620 404.280 ;
      LAYER met2 ;
        RECT 1769.900 400.000 1770.180 404.000 ;
      LAYER met2 ;
        RECT 1770.460 402.195 1774.680 404.280 ;
      LAYER met2 ;
        RECT 1774.960 400.000 1775.240 404.000 ;
      LAYER met2 ;
        RECT 1775.520 402.195 1779.740 404.280 ;
      LAYER met2 ;
        RECT 1780.020 400.000 1780.300 404.000 ;
      LAYER met2 ;
        RECT 1780.580 402.195 1784.340 404.280 ;
      LAYER met2 ;
        RECT 1784.620 400.000 1784.900 404.000 ;
      LAYER met2 ;
        RECT 1785.180 402.195 1789.400 404.280 ;
      LAYER met2 ;
        RECT 1789.680 400.000 1789.960 404.000 ;
      LAYER met2 ;
        RECT 1790.240 402.195 1794.000 404.280 ;
      LAYER met2 ;
        RECT 1794.280 400.000 1794.560 404.000 ;
      LAYER met2 ;
        RECT 1794.840 402.195 1799.060 404.280 ;
      LAYER met2 ;
        RECT 1799.340 400.000 1799.620 404.000 ;
      LAYER met2 ;
        RECT 1799.900 402.195 1803.660 404.280 ;
      LAYER met2 ;
        RECT 1803.940 400.000 1804.220 404.000 ;
      LAYER met2 ;
        RECT 1804.500 402.195 1808.720 404.280 ;
      LAYER met2 ;
        RECT 1809.000 400.000 1809.280 404.000 ;
      LAYER met2 ;
        RECT 1809.560 402.195 1813.320 404.280 ;
      LAYER met2 ;
        RECT 1813.600 400.000 1813.880 404.000 ;
      LAYER met2 ;
        RECT 1814.160 402.195 1818.380 404.280 ;
      LAYER met2 ;
        RECT 1818.660 400.000 1818.940 404.000 ;
      LAYER met2 ;
        RECT 1819.220 402.195 1822.980 404.280 ;
      LAYER met2 ;
        RECT 1823.260 400.000 1823.540 404.000 ;
      LAYER met2 ;
        RECT 1823.820 402.195 1828.040 404.280 ;
      LAYER met2 ;
        RECT 1828.320 400.000 1828.600 404.000 ;
      LAYER met2 ;
        RECT 1828.880 402.195 1832.640 404.280 ;
      LAYER met2 ;
        RECT 1832.920 400.000 1833.200 404.000 ;
      LAYER met2 ;
        RECT 1833.480 402.195 1837.700 404.280 ;
      LAYER met2 ;
        RECT 1837.980 400.000 1838.260 404.000 ;
      LAYER met2 ;
        RECT 1838.540 402.195 1842.300 404.280 ;
      LAYER met2 ;
        RECT 1842.580 400.000 1842.860 404.000 ;
      LAYER met2 ;
        RECT 1843.140 402.195 1847.360 404.280 ;
      LAYER met2 ;
        RECT 1847.640 400.000 1847.920 404.000 ;
      LAYER met2 ;
        RECT 1848.200 402.195 1852.420 404.280 ;
      LAYER met2 ;
        RECT 1852.700 400.000 1852.980 404.000 ;
      LAYER met2 ;
        RECT 1853.260 402.195 1857.020 404.280 ;
      LAYER met2 ;
        RECT 1857.300 400.000 1857.580 404.000 ;
      LAYER met2 ;
        RECT 1857.860 402.195 1862.080 404.280 ;
      LAYER met2 ;
        RECT 1862.360 400.000 1862.640 404.000 ;
      LAYER met2 ;
        RECT 1862.920 402.195 1866.680 404.280 ;
      LAYER met2 ;
        RECT 1866.960 400.000 1867.240 404.000 ;
      LAYER met2 ;
        RECT 1867.520 402.195 1871.740 404.280 ;
      LAYER met2 ;
        RECT 1872.020 400.000 1872.300 404.000 ;
      LAYER met2 ;
        RECT 1872.580 402.195 1876.340 404.280 ;
      LAYER met2 ;
        RECT 1876.620 400.000 1876.900 404.000 ;
      LAYER met2 ;
        RECT 1877.180 402.195 1881.400 404.280 ;
      LAYER met2 ;
        RECT 1881.680 400.000 1881.960 404.000 ;
      LAYER met2 ;
        RECT 1882.240 402.195 1886.000 404.280 ;
      LAYER met2 ;
        RECT 1886.280 400.000 1886.560 404.000 ;
      LAYER met2 ;
        RECT 1886.840 402.195 1891.060 404.280 ;
      LAYER met2 ;
        RECT 1891.340 400.000 1891.620 404.000 ;
      LAYER met2 ;
        RECT 1891.900 402.195 1895.660 404.280 ;
      LAYER met2 ;
        RECT 1895.940 400.000 1896.220 404.000 ;
      LAYER met2 ;
        RECT 1896.500 402.195 1900.720 404.280 ;
      LAYER met2 ;
        RECT 1901.000 400.000 1901.280 404.000 ;
      LAYER met2 ;
        RECT 1901.560 402.195 1905.320 404.280 ;
      LAYER met2 ;
        RECT 1905.600 400.000 1905.880 404.000 ;
      LAYER met2 ;
        RECT 1906.160 402.195 1910.380 404.280 ;
      LAYER met2 ;
        RECT 1910.660 400.000 1910.940 404.000 ;
      LAYER met2 ;
        RECT 1911.220 402.195 1914.980 404.280 ;
      LAYER met2 ;
        RECT 1915.260 400.000 1915.540 404.000 ;
      LAYER met2 ;
        RECT 1915.820 402.195 1920.040 404.280 ;
      LAYER met2 ;
        RECT 1920.320 400.000 1920.600 404.000 ;
      LAYER met2 ;
        RECT 1920.880 402.195 1925.100 404.280 ;
      LAYER met2 ;
        RECT 1925.380 400.000 1925.660 404.000 ;
      LAYER met2 ;
        RECT 1925.940 402.195 1929.700 404.280 ;
      LAYER met2 ;
        RECT 1929.980 400.000 1930.260 404.000 ;
      LAYER met2 ;
        RECT 1930.540 402.195 1934.760 404.280 ;
      LAYER met2 ;
        RECT 1935.040 400.000 1935.320 404.000 ;
      LAYER met2 ;
        RECT 1935.600 402.195 1939.360 404.280 ;
      LAYER met2 ;
        RECT 1939.640 400.000 1939.920 404.000 ;
      LAYER met2 ;
        RECT 1940.200 402.195 1944.420 404.280 ;
      LAYER met2 ;
        RECT 1944.700 400.000 1944.980 404.000 ;
      LAYER met2 ;
        RECT 1945.260 402.195 1949.020 404.280 ;
      LAYER met2 ;
        RECT 1949.300 400.000 1949.580 404.000 ;
      LAYER met2 ;
        RECT 1949.860 402.195 1954.080 404.280 ;
      LAYER met2 ;
        RECT 1954.360 400.000 1954.640 404.000 ;
      LAYER met2 ;
        RECT 1954.920 402.195 1958.680 404.280 ;
      LAYER met2 ;
        RECT 1958.960 400.000 1959.240 404.000 ;
      LAYER met2 ;
        RECT 1959.520 402.195 1963.740 404.280 ;
      LAYER met2 ;
        RECT 1964.020 400.000 1964.300 404.000 ;
      LAYER met2 ;
        RECT 1964.580 402.195 1968.340 404.280 ;
      LAYER met2 ;
        RECT 1968.620 400.000 1968.900 404.000 ;
      LAYER met2 ;
        RECT 1969.180 402.195 1973.400 404.280 ;
      LAYER met2 ;
        RECT 1973.680 400.000 1973.960 404.000 ;
      LAYER met2 ;
        RECT 1974.240 402.195 1978.000 404.280 ;
      LAYER met2 ;
        RECT 1978.280 400.000 1978.560 404.000 ;
      LAYER met2 ;
        RECT 1978.840 402.195 1983.060 404.280 ;
      LAYER met2 ;
        RECT 1983.340 400.000 1983.620 404.000 ;
      LAYER met2 ;
        RECT 1983.900 402.195 1987.660 404.280 ;
      LAYER met2 ;
        RECT 1987.940 400.000 1988.220 404.000 ;
      LAYER met2 ;
        RECT 1988.500 402.195 1992.720 404.280 ;
      LAYER met2 ;
        RECT 1993.000 400.000 1993.280 404.000 ;
      LAYER met2 ;
        RECT 1993.560 402.195 1997.780 404.280 ;
      LAYER met2 ;
        RECT 1998.060 400.000 1998.340 404.000 ;
      LAYER met2 ;
        RECT 1998.620 402.195 2002.380 404.280 ;
      LAYER met2 ;
        RECT 2002.660 400.000 2002.940 404.000 ;
      LAYER met2 ;
        RECT 2003.220 402.195 2007.440 404.280 ;
      LAYER met2 ;
        RECT 2007.720 400.000 2008.000 404.000 ;
      LAYER met2 ;
        RECT 2008.280 402.195 2012.040 404.280 ;
      LAYER met2 ;
        RECT 2012.320 400.000 2012.600 404.000 ;
      LAYER met2 ;
        RECT 2012.880 402.195 2017.100 404.280 ;
      LAYER met2 ;
        RECT 2017.380 400.000 2017.660 404.000 ;
      LAYER met2 ;
        RECT 2017.940 402.195 2021.700 404.280 ;
      LAYER met2 ;
        RECT 2021.980 400.000 2022.260 404.000 ;
      LAYER met2 ;
        RECT 2022.540 402.195 2026.760 404.280 ;
      LAYER met2 ;
        RECT 2027.040 400.000 2027.320 404.000 ;
      LAYER met2 ;
        RECT 2027.600 402.195 2031.360 404.280 ;
      LAYER met2 ;
        RECT 2031.640 400.000 2031.920 404.000 ;
      LAYER met2 ;
        RECT 2032.200 402.195 2036.420 404.280 ;
      LAYER met2 ;
        RECT 2036.700 400.000 2036.980 404.000 ;
      LAYER met2 ;
        RECT 2037.260 402.195 2041.020 404.280 ;
      LAYER met2 ;
        RECT 2041.300 400.000 2041.580 404.000 ;
      LAYER met2 ;
        RECT 2041.860 402.195 2046.080 404.280 ;
      LAYER met2 ;
        RECT 2046.360 400.000 2046.640 404.000 ;
      LAYER met2 ;
        RECT 2046.920 402.195 2050.680 404.280 ;
      LAYER met2 ;
        RECT 2050.960 400.000 2051.240 404.000 ;
      LAYER met2 ;
        RECT 2051.520 402.195 2055.740 404.280 ;
      LAYER met2 ;
        RECT 2056.020 400.000 2056.300 404.000 ;
      LAYER met2 ;
        RECT 2056.580 402.195 2060.340 404.280 ;
      LAYER met2 ;
        RECT 2060.620 400.000 2060.900 404.000 ;
      LAYER met2 ;
        RECT 2061.180 402.195 2065.400 404.280 ;
      LAYER met2 ;
        RECT 2065.680 400.000 2065.960 404.000 ;
      LAYER met2 ;
        RECT 2066.240 402.195 2070.460 404.280 ;
      LAYER met2 ;
        RECT 2070.740 400.000 2071.020 404.000 ;
      LAYER met2 ;
        RECT 2071.300 402.195 2075.060 404.280 ;
      LAYER met2 ;
        RECT 2075.340 400.000 2075.620 404.000 ;
      LAYER met2 ;
        RECT 2075.900 402.195 2080.120 404.280 ;
      LAYER met2 ;
        RECT 2080.400 400.000 2080.680 404.000 ;
      LAYER met2 ;
        RECT 2080.960 402.195 2084.720 404.280 ;
      LAYER met2 ;
        RECT 2085.000 400.000 2085.280 404.000 ;
      LAYER met2 ;
        RECT 2085.560 402.195 2089.780 404.280 ;
      LAYER met2 ;
        RECT 2090.060 400.000 2090.340 404.000 ;
      LAYER met2 ;
        RECT 2090.620 402.195 2094.380 404.280 ;
      LAYER met2 ;
        RECT 2094.660 400.000 2094.940 404.000 ;
      LAYER met2 ;
        RECT 2095.220 402.195 2099.440 404.280 ;
      LAYER met2 ;
        RECT 2099.720 400.000 2100.000 404.000 ;
      LAYER met2 ;
        RECT 2100.280 402.195 2104.040 404.280 ;
      LAYER met2 ;
        RECT 2104.320 400.000 2104.600 404.000 ;
      LAYER met2 ;
        RECT 2104.880 402.195 2109.100 404.280 ;
      LAYER met2 ;
        RECT 2109.380 400.000 2109.660 404.000 ;
      LAYER met2 ;
        RECT 2109.940 402.195 2113.700 404.280 ;
      LAYER met2 ;
        RECT 2113.980 400.000 2114.260 404.000 ;
      LAYER met2 ;
        RECT 2114.540 402.195 2118.760 404.280 ;
      LAYER met2 ;
        RECT 2119.040 400.000 2119.320 404.000 ;
      LAYER met2 ;
        RECT 2119.600 402.195 2123.360 404.280 ;
      LAYER met2 ;
        RECT 2123.640 400.000 2123.920 404.000 ;
      LAYER met2 ;
        RECT 2124.200 402.195 2128.420 404.280 ;
      LAYER met2 ;
        RECT 2128.700 400.000 2128.980 404.000 ;
      LAYER met2 ;
        RECT 2129.260 402.195 2133.020 404.280 ;
      LAYER met2 ;
        RECT 2133.300 400.000 2133.580 404.000 ;
      LAYER met2 ;
        RECT 2133.860 402.195 2138.080 404.280 ;
      LAYER met2 ;
        RECT 2138.360 400.000 2138.640 404.000 ;
      LAYER met2 ;
        RECT 2138.920 402.195 2143.140 404.280 ;
      LAYER met2 ;
        RECT 2143.420 400.000 2143.700 404.000 ;
      LAYER met2 ;
        RECT 2143.980 402.195 2147.740 404.280 ;
      LAYER met2 ;
        RECT 2148.020 400.000 2148.300 404.000 ;
      LAYER met2 ;
        RECT 2148.580 402.195 2152.800 404.280 ;
      LAYER met2 ;
        RECT 2153.080 400.000 2153.360 404.000 ;
      LAYER met2 ;
        RECT 2153.640 402.195 2157.400 404.280 ;
      LAYER met2 ;
        RECT 2157.680 400.000 2157.960 404.000 ;
      LAYER met2 ;
        RECT 2158.240 402.195 2162.460 404.280 ;
      LAYER met2 ;
        RECT 2162.740 400.000 2163.020 404.000 ;
      LAYER met2 ;
        RECT 2163.300 402.195 2167.060 404.280 ;
      LAYER met2 ;
        RECT 2167.340 400.000 2167.620 404.000 ;
      LAYER met2 ;
        RECT 2167.900 402.195 2172.120 404.280 ;
      LAYER met2 ;
        RECT 2172.400 400.000 2172.680 404.000 ;
      LAYER met2 ;
        RECT 2172.960 402.195 2176.720 404.280 ;
      LAYER met2 ;
        RECT 2177.000 400.000 2177.280 404.000 ;
      LAYER met2 ;
        RECT 2177.560 402.195 2181.780 404.280 ;
      LAYER met2 ;
        RECT 2182.060 400.000 2182.340 404.000 ;
      LAYER met2 ;
        RECT 2182.620 402.195 2186.380 404.280 ;
      LAYER met2 ;
        RECT 2186.660 400.000 2186.940 404.000 ;
      LAYER met2 ;
        RECT 2187.220 402.195 2191.440 404.280 ;
      LAYER met2 ;
        RECT 2191.720 400.000 2192.000 404.000 ;
      LAYER met2 ;
        RECT 2192.280 402.195 2196.040 404.280 ;
      LAYER met2 ;
        RECT 2196.320 400.000 2196.600 404.000 ;
      LAYER met2 ;
        RECT 2196.880 402.195 2201.100 404.280 ;
      LAYER met2 ;
        RECT 2201.380 400.000 2201.660 404.000 ;
      LAYER met2 ;
        RECT 2201.940 402.195 2205.700 404.280 ;
      LAYER met2 ;
        RECT 2205.980 400.000 2206.260 404.000 ;
      LAYER met2 ;
        RECT 2206.540 402.195 2210.760 404.280 ;
      LAYER met2 ;
        RECT 2211.040 400.000 2211.320 404.000 ;
      LAYER met2 ;
        RECT 2211.600 402.195 2215.820 404.280 ;
      LAYER met2 ;
        RECT 2216.100 400.000 2216.380 404.000 ;
      LAYER met2 ;
        RECT 2216.660 402.195 2220.420 404.280 ;
      LAYER met2 ;
        RECT 2220.700 400.000 2220.980 404.000 ;
      LAYER met2 ;
        RECT 2221.260 402.195 2225.480 404.280 ;
      LAYER met2 ;
        RECT 2225.760 400.000 2226.040 404.000 ;
      LAYER met2 ;
        RECT 2226.320 402.195 2230.080 404.280 ;
      LAYER met2 ;
        RECT 2230.360 400.000 2230.640 404.000 ;
      LAYER met2 ;
        RECT 2230.920 402.195 2235.140 404.280 ;
      LAYER met2 ;
        RECT 2235.420 400.000 2235.700 404.000 ;
      LAYER met2 ;
        RECT 2235.980 402.195 2239.740 404.280 ;
      LAYER met2 ;
        RECT 2240.020 400.000 2240.300 404.000 ;
      LAYER met2 ;
        RECT 2240.580 402.195 2244.800 404.280 ;
      LAYER met2 ;
        RECT 2245.080 400.000 2245.360 404.000 ;
      LAYER met2 ;
        RECT 2245.640 402.195 2249.400 404.280 ;
      LAYER met2 ;
        RECT 2249.680 400.000 2249.960 404.000 ;
      LAYER met2 ;
        RECT 2250.240 402.195 2254.460 404.280 ;
      LAYER met2 ;
        RECT 2254.740 400.000 2255.020 404.000 ;
      LAYER met2 ;
        RECT 2255.300 402.195 2259.060 404.280 ;
      LAYER met2 ;
        RECT 2259.340 400.000 2259.620 404.000 ;
      LAYER met2 ;
        RECT 2259.900 402.195 2264.120 404.280 ;
      LAYER met2 ;
        RECT 2264.400 400.000 2264.680 404.000 ;
      LAYER met2 ;
        RECT 2264.960 402.195 2268.720 404.280 ;
      LAYER met2 ;
        RECT 2269.000 400.000 2269.280 404.000 ;
      LAYER met2 ;
        RECT 2269.560 402.195 2273.780 404.280 ;
      LAYER met2 ;
        RECT 2274.060 400.000 2274.340 404.000 ;
      LAYER met2 ;
        RECT 2274.620 402.195 2278.380 404.280 ;
      LAYER met2 ;
        RECT 2278.660 400.000 2278.940 404.000 ;
      LAYER met2 ;
        RECT 2279.220 402.195 2283.440 404.280 ;
      LAYER met2 ;
        RECT 2283.720 400.000 2284.000 404.000 ;
      LAYER met2 ;
        RECT 2284.280 402.195 2288.500 404.280 ;
      LAYER met2 ;
        RECT 2288.780 400.000 2289.060 404.000 ;
      LAYER met2 ;
        RECT 2289.340 402.195 2293.100 404.280 ;
      LAYER met2 ;
        RECT 2293.380 400.000 2293.660 404.000 ;
      LAYER met2 ;
        RECT 2293.940 402.195 2298.160 404.280 ;
      LAYER met2 ;
        RECT 2298.440 400.000 2298.720 404.000 ;
      LAYER met2 ;
        RECT 2299.000 402.195 2302.760 404.280 ;
      LAYER met2 ;
        RECT 2303.040 400.000 2303.320 404.000 ;
      LAYER met2 ;
        RECT 2303.600 402.195 2307.820 404.280 ;
      LAYER met2 ;
        RECT 2308.100 400.000 2308.380 404.000 ;
      LAYER met2 ;
        RECT 2308.660 402.195 2312.420 404.280 ;
      LAYER met2 ;
        RECT 2312.700 400.000 2312.980 404.000 ;
      LAYER met2 ;
        RECT 2313.260 402.195 2317.480 404.280 ;
      LAYER met2 ;
        RECT 2317.760 400.000 2318.040 404.000 ;
      LAYER met2 ;
        RECT 2318.320 402.195 2322.080 404.280 ;
      LAYER met2 ;
        RECT 2322.360 400.000 2322.640 404.000 ;
      LAYER met2 ;
        RECT 2322.920 402.195 2327.140 404.280 ;
      LAYER met2 ;
        RECT 2327.420 400.000 2327.700 404.000 ;
      LAYER met2 ;
        RECT 2327.980 402.195 2331.740 404.280 ;
      LAYER met2 ;
        RECT 2332.020 400.000 2332.300 404.000 ;
      LAYER met2 ;
        RECT 2332.580 402.195 2336.800 404.280 ;
      LAYER met2 ;
        RECT 2337.080 400.000 2337.360 404.000 ;
      LAYER met2 ;
        RECT 2337.640 402.195 2341.400 404.280 ;
      LAYER met2 ;
        RECT 2341.680 400.000 2341.960 404.000 ;
      LAYER met2 ;
        RECT 2342.240 402.195 2346.460 404.280 ;
      LAYER met2 ;
        RECT 2346.740 400.000 2347.020 404.000 ;
      LAYER met2 ;
        RECT 2347.300 402.195 2351.060 404.280 ;
      LAYER met2 ;
        RECT 2351.340 400.000 2351.620 404.000 ;
      LAYER met2 ;
        RECT 2351.900 402.195 2356.120 404.280 ;
      LAYER met2 ;
        RECT 2356.400 400.000 2356.680 404.000 ;
      LAYER met2 ;
        RECT 2356.960 402.195 2361.180 404.280 ;
      LAYER met2 ;
        RECT 2361.460 400.000 2361.740 404.000 ;
      LAYER met2 ;
        RECT 2362.020 402.195 2365.780 404.280 ;
      LAYER met2 ;
        RECT 2366.060 400.000 2366.340 404.000 ;
      LAYER met2 ;
        RECT 2366.620 402.195 2370.840 404.280 ;
      LAYER met2 ;
        RECT 2371.120 400.000 2371.400 404.000 ;
      LAYER met2 ;
        RECT 2371.680 402.195 2375.440 404.280 ;
      LAYER met2 ;
        RECT 2375.720 400.000 2376.000 404.000 ;
      LAYER met2 ;
        RECT 2376.280 402.195 2380.500 404.280 ;
      LAYER met2 ;
        RECT 2380.780 400.000 2381.060 404.000 ;
      LAYER met2 ;
        RECT 2381.340 402.195 2385.100 404.280 ;
      LAYER met2 ;
        RECT 2385.380 400.000 2385.660 404.000 ;
      LAYER met2 ;
        RECT 2385.940 402.195 2390.160 404.280 ;
      LAYER met2 ;
        RECT 2390.440 400.000 2390.720 404.000 ;
      LAYER met2 ;
        RECT 2391.000 402.195 2394.760 404.280 ;
      LAYER met2 ;
        RECT 2395.040 400.000 2395.320 404.000 ;
      LAYER met2 ;
        RECT 2395.600 402.195 2399.820 404.280 ;
      LAYER met2 ;
        RECT 2400.100 400.000 2400.380 404.000 ;
      LAYER met2 ;
        RECT 2400.660 402.195 2404.420 404.280 ;
      LAYER met2 ;
        RECT 2404.700 400.000 2404.980 404.000 ;
      LAYER met2 ;
        RECT 2405.260 402.195 2409.480 404.280 ;
      LAYER met2 ;
        RECT 2409.760 400.000 2410.040 404.000 ;
      LAYER met2 ;
        RECT 2410.320 402.195 2414.080 404.280 ;
      LAYER met2 ;
        RECT 2414.360 400.000 2414.640 404.000 ;
      LAYER met2 ;
        RECT 2414.920 402.195 2419.140 404.280 ;
      LAYER met2 ;
        RECT 2419.420 400.000 2419.700 404.000 ;
      LAYER met2 ;
        RECT 2419.980 402.195 2423.740 404.280 ;
      LAYER met2 ;
        RECT 2424.020 400.000 2424.300 404.000 ;
      LAYER met2 ;
        RECT 2424.580 402.195 2428.800 404.280 ;
      LAYER met2 ;
        RECT 2429.080 400.000 2429.360 404.000 ;
      LAYER met2 ;
        RECT 2429.640 402.195 2433.860 404.280 ;
      LAYER met2 ;
        RECT 2434.140 400.000 2434.420 404.000 ;
      LAYER met2 ;
        RECT 2434.700 402.195 2438.460 404.280 ;
      LAYER met2 ;
        RECT 2438.740 400.000 2439.020 404.000 ;
      LAYER met2 ;
        RECT 2439.300 402.195 2443.520 404.280 ;
      LAYER met2 ;
        RECT 2443.800 400.000 2444.080 404.000 ;
      LAYER met2 ;
        RECT 2444.360 402.195 2448.120 404.280 ;
      LAYER met2 ;
        RECT 2448.400 400.000 2448.680 404.000 ;
      LAYER met2 ;
        RECT 2448.960 402.195 2453.180 404.280 ;
      LAYER met2 ;
        RECT 2453.460 400.000 2453.740 404.000 ;
      LAYER met2 ;
        RECT 2454.020 402.195 2457.780 404.280 ;
      LAYER met2 ;
        RECT 2458.060 400.000 2458.340 404.000 ;
      LAYER met2 ;
        RECT 2458.620 402.195 2462.840 404.280 ;
      LAYER met2 ;
        RECT 2463.120 400.000 2463.400 404.000 ;
      LAYER met2 ;
        RECT 2463.680 402.195 2467.440 404.280 ;
      LAYER met2 ;
        RECT 2467.720 400.000 2468.000 404.000 ;
      LAYER met2 ;
        RECT 2468.280 402.195 2472.500 404.280 ;
      LAYER met2 ;
        RECT 2472.780 400.000 2473.060 404.000 ;
      LAYER met2 ;
        RECT 2473.340 402.195 2477.100 404.280 ;
      LAYER met2 ;
        RECT 2477.380 400.000 2477.660 404.000 ;
      LAYER met2 ;
        RECT 2477.940 402.195 2482.160 404.280 ;
      LAYER met2 ;
        RECT 2482.440 400.000 2482.720 404.000 ;
      LAYER met2 ;
        RECT 2483.000 402.195 2486.760 404.280 ;
      LAYER met2 ;
        RECT 2487.040 400.000 2487.320 404.000 ;
      LAYER met2 ;
        RECT 2487.600 402.195 2491.820 404.280 ;
      LAYER met2 ;
        RECT 2492.100 400.000 2492.380 404.000 ;
      LAYER met2 ;
        RECT 2492.660 402.195 2496.420 404.280 ;
      LAYER met2 ;
        RECT 2496.700 400.000 2496.980 404.000 ;
      LAYER met2 ;
        RECT 2497.260 402.195 2501.480 404.280 ;
      LAYER met2 ;
        RECT 2501.760 400.000 2502.040 404.000 ;
      LAYER met2 ;
        RECT 2502.320 402.195 2506.540 404.280 ;
      LAYER met2 ;
        RECT 2506.820 400.000 2507.100 404.000 ;
      LAYER met2 ;
        RECT 2507.380 402.195 2511.140 404.280 ;
      LAYER met2 ;
        RECT 2511.420 400.000 2511.700 404.000 ;
      LAYER met2 ;
        RECT 2511.980 402.195 2516.200 404.280 ;
      LAYER met2 ;
        RECT 2516.480 400.000 2516.760 404.000 ;
      LAYER met2 ;
        RECT 2517.040 402.195 2520.800 404.280 ;
      LAYER met2 ;
        RECT 2521.080 400.000 2521.360 404.000 ;
      LAYER met2 ;
        RECT 2521.640 402.195 2525.860 404.280 ;
      LAYER met2 ;
        RECT 2526.140 400.000 2526.420 404.000 ;
      LAYER met2 ;
        RECT 2526.700 402.195 2530.460 404.280 ;
      LAYER met2 ;
        RECT 2530.740 400.000 2531.020 404.000 ;
      LAYER met2 ;
        RECT 2531.300 402.195 2535.520 404.280 ;
      LAYER met2 ;
        RECT 2535.800 400.000 2536.080 404.000 ;
      LAYER met2 ;
        RECT 2536.360 402.195 2540.120 404.280 ;
      LAYER met2 ;
        RECT 2540.400 400.000 2540.680 404.000 ;
      LAYER met2 ;
        RECT 2540.960 402.195 2545.180 404.280 ;
      LAYER met2 ;
        RECT 2545.460 400.000 2545.740 404.000 ;
      LAYER met2 ;
        RECT 2546.020 402.195 2549.780 404.280 ;
      LAYER met2 ;
        RECT 2550.060 400.000 2550.340 404.000 ;
      LAYER met2 ;
        RECT 2550.620 402.195 2554.840 404.280 ;
      LAYER met2 ;
        RECT 2555.120 400.000 2555.400 404.000 ;
      LAYER met2 ;
        RECT 2555.680 402.195 2559.440 404.280 ;
      LAYER met2 ;
        RECT 2559.720 400.000 2560.000 404.000 ;
      LAYER met2 ;
        RECT 2560.280 402.195 2564.500 404.280 ;
      LAYER met2 ;
        RECT 2564.780 400.000 2565.060 404.000 ;
      LAYER met2 ;
        RECT 2565.340 402.195 2569.100 404.280 ;
      LAYER met2 ;
        RECT 2569.380 400.000 2569.660 404.000 ;
      LAYER met2 ;
        RECT 2569.940 402.195 2574.160 404.280 ;
      LAYER met2 ;
        RECT 2574.440 400.000 2574.720 404.000 ;
      LAYER met2 ;
        RECT 2575.000 402.195 2579.220 404.280 ;
      LAYER met2 ;
        RECT 2579.500 400.000 2579.780 404.000 ;
      LAYER met2 ;
        RECT 2580.060 402.195 2583.820 404.280 ;
      LAYER met2 ;
        RECT 2584.100 400.000 2584.380 404.000 ;
      LAYER met2 ;
        RECT 2584.660 402.195 2588.880 404.280 ;
      LAYER met2 ;
        RECT 2589.160 400.000 2589.440 404.000 ;
      LAYER met2 ;
        RECT 2589.720 402.195 2593.480 404.280 ;
      LAYER met2 ;
        RECT 2593.760 400.000 2594.040 404.000 ;
      LAYER met2 ;
        RECT 2594.320 402.195 2598.540 404.280 ;
      LAYER met2 ;
        RECT 2598.820 400.000 2599.100 404.000 ;
      LAYER met2 ;
        RECT 2599.380 402.195 2603.140 404.280 ;
      LAYER met2 ;
        RECT 2603.420 400.000 2603.700 404.000 ;
      LAYER met2 ;
        RECT 2603.980 402.195 2608.200 404.280 ;
      LAYER met2 ;
        RECT 2608.480 400.000 2608.760 404.000 ;
      LAYER met2 ;
        RECT 2609.040 402.195 2612.800 404.280 ;
      LAYER met2 ;
        RECT 2613.080 400.000 2613.360 404.000 ;
      LAYER met2 ;
        RECT 2613.640 402.195 2617.860 404.280 ;
      LAYER met2 ;
        RECT 2618.140 400.000 2618.420 404.000 ;
      LAYER met2 ;
        RECT 2618.700 402.195 2622.460 404.280 ;
      LAYER met2 ;
        RECT 2622.740 400.000 2623.020 404.000 ;
      LAYER met2 ;
        RECT 2623.300 402.195 2627.520 404.280 ;
      LAYER met2 ;
        RECT 2627.800 400.000 2628.080 404.000 ;
      LAYER met2 ;
        RECT 2628.360 402.195 2632.120 404.280 ;
      LAYER met2 ;
        RECT 2632.400 400.000 2632.680 404.000 ;
      LAYER met2 ;
        RECT 2632.960 402.195 2637.180 404.280 ;
      LAYER met2 ;
        RECT 2637.460 400.000 2637.740 404.000 ;
      LAYER met2 ;
        RECT 2638.020 402.195 2641.780 404.280 ;
      LAYER met2 ;
        RECT 2642.060 400.000 2642.340 404.000 ;
      LAYER met2 ;
        RECT 2642.620 402.195 2646.840 404.280 ;
      LAYER met2 ;
        RECT 2647.120 400.000 2647.400 404.000 ;
      LAYER via2 ;
        RECT 646.390 3264.200 646.670 3264.480 ;
        RECT 668.010 3264.200 668.290 3264.480 ;
        RECT 1293.150 3264.200 1293.430 3264.480 ;
        RECT 1890.690 3264.200 1890.970 3264.480 ;
        RECT 1917.830 3264.200 1918.110 3264.480 ;
        RECT 2542.050 3264.200 2542.330 3264.480 ;
        RECT 2566.890 3264.200 2567.170 3264.480 ;
        RECT 289.430 3230.200 289.710 3230.480 ;
        RECT 288.970 3224.760 289.250 3225.040 ;
        RECT 288.510 3215.920 288.790 3216.200 ;
        RECT 288.050 3209.800 288.330 3210.080 ;
        RECT 287.590 3201.640 287.870 3201.920 ;
        RECT 287.130 3196.200 287.410 3196.480 ;
        RECT 286.670 3188.040 286.950 3188.320 ;
        RECT 286.210 2898.360 286.490 2898.640 ;
        RECT 688.250 3248.275 688.530 3248.555 ;
        RECT 1317.530 3258.080 1317.810 3258.360 ;
        RECT 821.190 3251.280 821.470 3251.560 ;
        RECT 869.030 3251.280 869.310 3251.560 ;
        RECT 941.710 3230.200 941.990 3230.480 ;
        RECT 696.990 2948.000 697.270 2948.280 ;
        RECT 939.410 2898.360 939.690 2898.640 ;
        RECT 337.730 2794.320 338.010 2794.600 ;
        RECT 344.630 2794.320 344.910 2794.600 ;
        RECT 351.530 2794.320 351.810 2794.600 ;
        RECT 358.430 2794.320 358.710 2794.600 ;
        RECT 362.110 2794.320 362.390 2794.600 ;
        RECT 365.330 2794.320 365.610 2794.600 ;
        RECT 368.550 2794.320 368.830 2794.600 ;
        RECT 371.310 2794.320 371.590 2794.600 ;
        RECT 374.990 2794.320 375.270 2794.600 ;
        RECT 378.670 2794.320 378.950 2794.600 ;
        RECT 380.050 2794.320 380.330 2794.600 ;
        RECT 384.650 2794.320 384.930 2794.600 ;
        RECT 386.950 2794.320 387.230 2794.600 ;
        RECT 390.630 2794.320 390.910 2794.600 ;
        RECT 392.470 2794.320 392.750 2794.600 ;
        RECT 396.610 2794.320 396.890 2794.600 ;
        RECT 399.830 2794.320 400.110 2794.600 ;
        RECT 403.970 2794.320 404.250 2794.600 ;
        RECT 406.270 2794.320 406.550 2794.600 ;
        RECT 409.950 2794.320 410.230 2794.600 ;
        RECT 413.630 2794.320 413.910 2794.600 ;
        RECT 414.550 2794.320 414.830 2794.600 ;
        RECT 418.690 2794.320 418.970 2794.600 ;
        RECT 420.990 2794.320 421.270 2794.600 ;
        RECT 427.430 2794.320 427.710 2794.600 ;
        RECT 432.030 2794.320 432.310 2794.600 ;
        RECT 305.070 2714.760 305.350 2715.040 ;
        RECT 351.070 2792.280 351.350 2792.560 ;
        RECT 397.070 2793.640 397.350 2793.920 ;
        RECT 410.410 2790.920 410.690 2791.200 ;
        RECT 426.970 2793.640 427.250 2793.920 ;
        RECT 434.330 2794.320 434.610 2794.600 ;
        RECT 439.390 2794.320 439.670 2794.600 ;
        RECT 441.230 2794.320 441.510 2794.600 ;
        RECT 444.450 2794.320 444.730 2794.600 ;
        RECT 448.130 2794.320 448.410 2794.600 ;
        RECT 450.430 2794.320 450.710 2794.600 ;
        RECT 455.030 2794.320 455.310 2794.600 ;
        RECT 461.930 2794.320 462.210 2794.600 ;
        RECT 466.530 2794.320 466.810 2794.600 ;
        RECT 468.370 2794.320 468.650 2794.600 ;
        RECT 475.730 2794.320 476.010 2794.600 ;
        RECT 478.490 2794.320 478.770 2794.600 ;
        RECT 482.630 2794.320 482.910 2794.600 ;
        RECT 484.930 2794.320 485.210 2794.600 ;
        RECT 489.070 2794.320 489.350 2794.600 ;
        RECT 492.750 2794.320 493.030 2794.600 ;
        RECT 496.430 2794.320 496.710 2794.600 ;
        RECT 433.870 2793.640 434.150 2793.920 ;
        RECT 455.490 2793.640 455.770 2793.920 ;
        RECT 462.390 2793.640 462.670 2793.920 ;
        RECT 468.830 2793.640 469.110 2793.920 ;
        RECT 475.270 2793.640 475.550 2793.920 ;
        RECT 501.950 2794.320 502.230 2794.600 ;
        RECT 509.770 2794.320 510.050 2794.600 ;
        RECT 513.910 2794.320 514.190 2794.600 ;
        RECT 517.130 2794.320 517.410 2794.600 ;
        RECT 524.030 2794.320 524.310 2794.600 ;
        RECT 526.790 2794.320 527.070 2794.600 ;
        RECT 530.930 2794.320 531.210 2794.600 ;
        RECT 537.370 2794.320 537.650 2794.600 ;
        RECT 539.210 2794.320 539.490 2794.600 ;
        RECT 544.270 2794.320 544.550 2794.600 ;
        RECT 551.630 2794.320 551.910 2794.600 ;
        RECT 500.110 2792.960 500.390 2793.240 ;
        RECT 501.030 2793.640 501.310 2793.920 ;
        RECT 508.850 2793.640 509.130 2793.920 ;
        RECT 510.230 2793.640 510.510 2793.920 ;
        RECT 520.810 2792.960 521.090 2793.240 ;
        RECT 534.610 2793.640 534.890 2793.920 ;
        RECT 541.510 2792.960 541.790 2793.240 ;
        RECT 686.410 2714.760 686.690 2715.040 ;
        RECT 942.170 3224.760 942.450 3225.040 ;
        RECT 942.630 3215.920 942.910 3216.200 ;
        RECT 943.090 3209.800 943.370 3210.080 ;
        RECT 943.550 3201.640 943.830 3201.920 ;
        RECT 944.010 3196.200 944.290 3196.480 ;
        RECT 944.470 3188.040 944.750 3188.320 ;
        RECT 1332.250 3249.240 1332.530 3249.520 ;
        RECT 1345.590 2946.640 1345.870 2946.920 ;
        RECT 1345.590 2935.760 1345.870 2936.040 ;
        RECT 1352.030 2901.760 1352.310 2902.040 ;
        RECT 1054.870 2799.760 1055.150 2800.040 ;
        RECT 1053.030 2795.680 1053.310 2795.960 ;
        RECT 979.890 2794.320 980.170 2794.600 ;
        RECT 1013.930 2794.320 1014.210 2794.600 ;
        RECT 1018.990 2794.320 1019.270 2794.600 ;
        RECT 1020.830 2794.320 1021.110 2794.600 ;
        RECT 1027.730 2794.320 1028.010 2794.600 ;
        RECT 1034.630 2794.320 1034.910 2794.600 ;
        RECT 1042.450 2794.320 1042.730 2794.600 ;
        RECT 986.790 2793.640 987.070 2793.920 ;
        RECT 1001.050 2793.640 1001.330 2793.920 ;
        RECT 1010.710 2792.960 1010.990 2793.240 ;
        RECT 1007.490 2788.200 1007.770 2788.480 ;
        RECT 1024.510 2792.960 1024.790 2793.240 ;
        RECT 1045.210 2792.960 1045.490 2793.240 ;
        RECT 1038.310 2788.200 1038.590 2788.480 ;
        RECT 1034.630 2787.520 1034.910 2787.800 ;
        RECT 1041.530 2787.520 1041.810 2787.800 ;
        RECT 1048.430 2787.520 1048.710 2787.800 ;
        RECT 1059.010 2794.320 1059.290 2794.600 ;
        RECT 1065.450 2794.320 1065.730 2794.600 ;
        RECT 1069.590 2794.320 1069.870 2794.600 ;
        RECT 1082.930 2794.320 1083.210 2794.600 ;
        RECT 1087.530 2794.320 1087.810 2794.600 ;
        RECT 1089.830 2794.320 1090.110 2794.600 ;
        RECT 1094.430 2794.320 1094.710 2794.600 ;
        RECT 1096.730 2794.320 1097.010 2794.600 ;
        RECT 1100.870 2794.320 1101.150 2794.600 ;
        RECT 1103.630 2794.320 1103.910 2794.600 ;
        RECT 1105.470 2794.320 1105.750 2794.600 ;
        RECT 1110.530 2794.320 1110.810 2794.600 ;
        RECT 1111.450 2794.320 1111.730 2794.600 ;
        RECT 1118.350 2794.320 1118.630 2794.600 ;
        RECT 1124.330 2794.320 1124.610 2794.600 ;
        RECT 1129.390 2794.320 1129.670 2794.600 ;
        RECT 1131.230 2794.320 1131.510 2794.600 ;
        RECT 1135.830 2794.320 1136.110 2794.600 ;
        RECT 1138.130 2794.320 1138.410 2794.600 ;
        RECT 1139.970 2794.320 1140.250 2794.600 ;
        RECT 1145.030 2794.320 1145.310 2794.600 ;
        RECT 1146.410 2794.320 1146.690 2794.600 ;
        RECT 1151.930 2794.320 1152.210 2794.600 ;
        RECT 1158.830 2794.320 1159.110 2794.600 ;
        RECT 1165.270 2794.320 1165.550 2794.600 ;
        RECT 1172.630 2794.320 1172.910 2794.600 ;
        RECT 1179.530 2794.320 1179.810 2794.600 ;
        RECT 1186.430 2794.320 1186.710 2794.600 ;
        RECT 1200.230 2794.320 1200.510 2794.600 ;
        RECT 1076.490 2793.640 1076.770 2793.920 ;
        RECT 1055.330 2788.200 1055.610 2788.480 ;
        RECT 1062.230 2787.520 1062.510 2787.800 ;
        RECT 1069.130 2787.520 1069.410 2787.800 ;
        RECT 1076.030 2787.520 1076.310 2787.800 ;
        RECT 1083.390 2793.640 1083.670 2793.920 ;
        RECT 1089.370 2793.640 1089.650 2793.920 ;
        RECT 1117.430 2792.280 1117.710 2792.560 ;
        RECT 1122.030 2793.640 1122.310 2793.920 ;
        RECT 1130.770 2793.640 1131.050 2793.920 ;
        RECT 1152.390 2792.280 1152.670 2792.560 ;
        RECT 1159.290 2791.600 1159.570 2791.880 ;
        RECT 1159.290 2790.920 1159.570 2791.200 ;
        RECT 1165.730 2793.640 1166.010 2793.920 ;
        RECT 1166.190 2792.960 1166.470 2793.240 ;
        RECT 1173.090 2793.640 1173.370 2793.920 ;
        RECT 1179.990 2793.640 1180.270 2793.920 ;
        RECT 1186.890 2793.640 1187.170 2793.920 ;
        RECT 1193.790 2791.600 1194.070 2791.880 ;
        RECT 1193.330 2790.240 1193.610 2790.520 ;
        RECT 1536.950 3230.200 1537.230 3230.480 ;
        RECT 1408.150 2894.960 1408.430 2895.240 ;
        RECT 1410.450 2146.960 1410.730 2147.240 ;
        RECT 1410.450 2126.560 1410.730 2126.840 ;
        RECT 1410.450 2111.600 1410.730 2111.880 ;
        RECT 1410.450 2091.200 1410.730 2091.480 ;
        RECT 1409.530 2086.440 1409.810 2086.720 ;
        RECT 1409.070 2055.840 1409.350 2056.120 ;
        RECT 1408.610 2051.080 1408.890 2051.360 ;
        RECT 1409.070 2046.320 1409.350 2046.600 ;
        RECT 1409.530 2036.120 1409.810 2036.400 ;
        RECT 1409.070 2021.160 1409.350 2021.440 ;
        RECT 1410.450 2015.720 1410.730 2016.000 ;
        RECT 1410.450 2010.960 1410.730 2011.240 ;
        RECT 1409.530 1965.400 1409.810 1965.680 ;
        RECT 1410.450 1955.200 1410.730 1955.480 ;
        RECT 1408.610 1894.680 1408.890 1894.960 ;
        RECT 1408.610 1823.960 1408.890 1824.240 ;
        RECT 1408.610 1819.200 1408.890 1819.480 ;
        RECT 1408.610 1813.760 1408.890 1814.040 ;
        RECT 1408.610 1809.000 1408.890 1809.280 ;
        RECT 1408.610 1798.800 1408.890 1799.080 ;
        RECT 1409.070 1794.040 1409.350 1794.320 ;
        RECT 1408.610 1778.400 1408.890 1778.680 ;
        RECT 1408.610 1773.640 1408.890 1773.920 ;
        RECT 1408.610 1768.200 1408.890 1768.480 ;
        RECT 1408.610 1763.440 1408.890 1763.720 ;
        RECT 1408.610 1753.240 1408.890 1753.520 ;
        RECT 1409.990 1732.840 1410.270 1733.120 ;
        RECT 1410.450 1717.880 1410.730 1718.160 ;
        RECT 1409.990 1713.120 1410.270 1713.400 ;
        RECT 1409.530 1702.920 1409.810 1703.200 ;
        RECT 1409.070 1698.160 1409.350 1698.440 ;
        RECT 1409.530 1692.720 1409.810 1693.000 ;
        RECT 1409.530 1687.960 1409.810 1688.240 ;
        RECT 1410.450 1672.320 1410.730 1672.600 ;
        RECT 1409.530 1667.560 1409.810 1667.840 ;
        RECT 1409.530 1647.160 1409.810 1647.440 ;
        RECT 1410.450 1642.400 1410.730 1642.680 ;
        RECT 1410.450 1632.200 1410.730 1632.480 ;
        RECT 1414.130 2142.200 1414.410 2142.480 ;
        RECT 1414.130 2136.760 1414.410 2137.040 ;
        RECT 1413.670 2132.000 1413.950 2132.280 ;
        RECT 1414.130 2121.800 1414.410 2122.080 ;
        RECT 1414.130 2117.040 1414.410 2117.320 ;
        RECT 1414.130 2106.840 1414.410 2107.120 ;
        RECT 1414.130 2101.400 1414.410 2101.680 ;
        RECT 1414.130 2096.640 1414.410 2096.920 ;
        RECT 1411.830 1788.600 1412.110 1788.880 ;
        RECT 1411.830 1682.520 1412.110 1682.800 ;
        RECT 1411.830 1677.760 1412.110 1678.040 ;
        RECT 1411.830 1662.800 1412.110 1663.080 ;
        RECT 1411.370 1636.960 1411.650 1637.240 ;
        RECT 1414.130 2081.680 1414.410 2081.960 ;
        RECT 1414.130 2076.240 1414.410 2076.520 ;
        RECT 1413.670 2071.480 1413.950 2071.760 ;
        RECT 1414.130 2066.040 1414.410 2066.320 ;
        RECT 1413.210 2025.920 1413.490 2026.200 ;
        RECT 1414.130 2061.280 1414.410 2061.560 ;
        RECT 1414.590 2040.880 1414.870 2041.160 ;
        RECT 1414.130 2030.680 1414.410 2030.960 ;
        RECT 1414.130 2005.520 1414.410 2005.800 ;
        RECT 1413.670 2000.760 1413.950 2001.040 ;
        RECT 1414.130 1995.320 1414.410 1995.600 ;
        RECT 1414.130 1990.560 1414.410 1990.840 ;
        RECT 1414.130 1985.800 1414.410 1986.080 ;
        RECT 1414.130 1980.360 1414.410 1980.640 ;
        RECT 1414.130 1975.600 1414.410 1975.880 ;
        RECT 1414.130 1970.160 1414.410 1970.440 ;
        RECT 1414.130 1959.960 1414.410 1960.240 ;
        RECT 1413.670 1950.440 1413.950 1950.720 ;
        RECT 1413.670 1945.000 1413.950 1945.280 ;
        RECT 1413.670 1940.240 1413.950 1940.520 ;
        RECT 1413.670 1934.800 1413.950 1935.080 ;
        RECT 1413.670 1930.040 1413.950 1930.320 ;
        RECT 1413.670 1925.280 1413.950 1925.560 ;
        RECT 1414.130 1922.560 1414.410 1922.840 ;
        RECT 1414.130 1915.080 1414.410 1915.360 ;
        RECT 1414.130 1910.320 1414.410 1910.600 ;
        RECT 1414.130 1904.880 1414.410 1905.160 ;
        RECT 1414.130 1900.800 1414.410 1901.080 ;
        RECT 1414.130 1889.920 1414.410 1890.200 ;
        RECT 1414.130 1884.480 1414.410 1884.760 ;
        RECT 1414.130 1879.720 1414.410 1880.000 ;
        RECT 1414.130 1874.280 1414.410 1874.560 ;
        RECT 1414.130 1869.520 1414.410 1869.800 ;
        RECT 1413.670 1864.080 1413.950 1864.360 ;
        RECT 1414.130 1859.320 1414.410 1859.600 ;
        RECT 1414.130 1854.560 1414.410 1854.840 ;
        RECT 1413.670 1849.120 1413.950 1849.400 ;
        RECT 1414.130 1844.360 1414.410 1844.640 ;
        RECT 1414.130 1838.920 1414.410 1839.200 ;
        RECT 1414.130 1834.160 1414.410 1834.440 ;
        RECT 1414.130 1828.720 1414.410 1829.000 ;
        RECT 1414.130 1803.560 1414.410 1803.840 ;
        RECT 1414.130 1783.840 1414.410 1784.120 ;
        RECT 1413.210 1758.680 1413.490 1758.960 ;
        RECT 1412.750 1748.480 1413.030 1748.760 ;
        RECT 1414.130 1743.040 1414.410 1743.320 ;
        RECT 1414.130 1738.280 1414.410 1738.560 ;
        RECT 1414.130 1728.080 1414.410 1728.360 ;
        RECT 1413.670 1723.320 1413.950 1723.600 ;
        RECT 1414.130 1707.680 1414.410 1707.960 ;
        RECT 1414.130 1652.600 1414.410 1652.880 ;
        RECT 1535.570 3224.760 1535.850 3225.040 ;
        RECT 1535.570 3217.280 1535.850 3217.560 ;
        RECT 1538.330 3210.480 1538.610 3210.760 ;
        RECT 1538.330 3202.320 1538.610 3202.600 ;
        RECT 1533.270 3196.880 1533.550 3197.160 ;
        RECT 1534.190 3189.400 1534.470 3189.680 ;
        RECT 1538.330 2899.040 1538.610 2899.320 ;
        RECT 1935.770 3249.240 1936.050 3249.520 ;
        RECT 2190.610 3230.200 2190.890 3230.480 ;
        RECT 1732.910 2795.680 1733.190 2795.960 ;
        RECT 1613.310 2794.320 1613.590 2794.600 ;
        RECT 1642.750 2794.320 1643.030 2794.600 ;
        RECT 1652.870 2794.320 1653.150 2794.600 ;
        RECT 1659.310 2794.320 1659.590 2794.600 ;
        RECT 1669.430 2794.320 1669.710 2794.600 ;
        RECT 1670.350 2794.320 1670.630 2794.600 ;
        RECT 1677.250 2794.320 1677.530 2794.600 ;
        RECT 1695.190 2794.320 1695.470 2794.600 ;
        RECT 1699.330 2794.320 1699.610 2794.600 ;
        RECT 1706.230 2794.320 1706.510 2794.600 ;
        RECT 1712.670 2794.320 1712.950 2794.600 ;
        RECT 1718.190 2794.320 1718.470 2794.600 ;
        RECT 1723.710 2794.320 1723.990 2794.600 ;
        RECT 1728.770 2794.320 1729.050 2794.600 ;
        RECT 1741.190 2794.320 1741.470 2794.600 ;
        RECT 1747.630 2794.320 1747.910 2794.600 ;
        RECT 1760.050 2794.320 1760.330 2794.600 ;
        RECT 1596.290 2792.280 1596.570 2792.560 ;
        RECT 1587.090 2791.600 1587.370 2791.880 ;
        RECT 1600.890 2791.600 1601.170 2791.880 ;
        RECT 1636.770 2792.960 1637.050 2793.240 ;
        RECT 1642.290 2790.240 1642.570 2790.520 ;
        RECT 1688.750 2793.640 1689.030 2793.920 ;
        RECT 1682.310 2792.960 1682.590 2793.240 ;
        RECT 1648.270 2789.560 1648.550 2789.840 ;
        RECT 1617.910 2788.200 1618.190 2788.480 ;
        RECT 1624.810 2788.200 1625.090 2788.480 ;
        RECT 1628.490 2788.200 1628.770 2788.480 ;
        RECT 1580.190 2787.520 1580.470 2787.800 ;
        RECT 1593.990 2787.520 1594.270 2787.800 ;
        RECT 1601.350 2787.520 1601.630 2787.800 ;
        RECT 1607.790 2787.520 1608.070 2787.800 ;
        RECT 1614.690 2787.520 1614.970 2787.800 ;
        RECT 1621.590 2787.520 1621.870 2787.800 ;
        RECT 1631.710 2787.520 1631.990 2787.800 ;
        RECT 1649.650 2788.200 1649.930 2788.480 ;
        RECT 1649.190 2787.520 1649.470 2787.800 ;
        RECT 1752.690 2792.280 1752.970 2792.560 ;
        RECT 1759.590 2791.600 1759.870 2791.880 ;
        RECT 1766.490 2793.640 1766.770 2793.920 ;
        RECT 1780.290 2793.640 1780.570 2793.920 ;
        RECT 1787.190 2792.960 1787.470 2793.240 ;
        RECT 1773.390 2791.600 1773.670 2791.880 ;
        RECT 1794.090 2791.600 1794.370 2791.880 ;
        RECT 1683.690 2788.200 1683.970 2788.480 ;
        RECT 1718.190 2788.200 1718.470 2788.480 ;
        RECT 1760.510 2788.200 1760.790 2788.480 ;
        RECT 1656.090 2787.520 1656.370 2787.800 ;
        RECT 1662.990 2787.520 1663.270 2787.800 ;
        RECT 1669.890 2787.520 1670.170 2787.800 ;
        RECT 1676.790 2787.520 1677.070 2787.800 ;
        RECT 1684.150 2787.520 1684.430 2787.800 ;
        RECT 1690.590 2787.520 1690.870 2787.800 ;
        RECT 1697.490 2787.520 1697.770 2787.800 ;
        RECT 1704.390 2787.520 1704.670 2787.800 ;
        RECT 1711.290 2787.520 1711.570 2787.800 ;
        RECT 1718.650 2787.520 1718.930 2787.800 ;
        RECT 1725.090 2787.520 1725.370 2787.800 ;
        RECT 1731.990 2787.520 1732.270 2787.800 ;
        RECT 1738.890 2787.520 1739.170 2787.800 ;
        RECT 1745.790 2787.520 1746.070 2787.800 ;
        RECT 1752.690 2787.520 1752.970 2787.800 ;
        RECT 1760.050 2787.520 1760.330 2787.800 ;
        RECT 1766.490 2787.520 1766.770 2787.800 ;
        RECT 1773.850 2787.520 1774.130 2787.800 ;
        RECT 1780.290 2787.520 1780.570 2787.800 ;
        RECT 1787.190 2787.520 1787.470 2787.800 ;
        RECT 1794.550 2787.520 1794.830 2787.800 ;
        RECT 1828.130 2787.520 1828.410 2787.800 ;
        RECT 1869.530 2787.520 1869.810 2787.800 ;
        RECT 2191.070 3224.760 2191.350 3225.040 ;
        RECT 2191.530 3215.920 2191.810 3216.200 ;
        RECT 2191.990 3209.800 2192.270 3210.080 ;
        RECT 2192.450 3201.640 2192.730 3201.920 ;
        RECT 2192.910 3196.200 2193.190 3196.480 ;
        RECT 2193.370 3188.040 2193.650 3188.320 ;
        RECT 2193.830 2898.360 2194.110 2898.640 ;
        RECT 2582.070 3249.240 2582.350 3249.520 ;
        RECT 2594.490 2946.640 2594.770 2946.920 ;
        RECT 2594.490 2938.480 2594.770 2938.760 ;
        RECT 2242.590 2794.320 2242.870 2794.600 ;
        RECT 2256.390 2794.320 2256.670 2794.600 ;
        RECT 2263.290 2794.320 2263.570 2794.600 ;
        RECT 2268.350 2794.320 2268.630 2794.600 ;
        RECT 2270.190 2794.320 2270.470 2794.600 ;
        RECT 2277.090 2794.320 2277.370 2794.600 ;
        RECT 2283.990 2794.320 2284.270 2794.600 ;
        RECT 2290.890 2794.320 2291.170 2794.600 ;
        RECT 2297.790 2794.320 2298.070 2794.600 ;
        RECT 2304.690 2794.320 2304.970 2794.600 ;
        RECT 2308.830 2794.320 2309.110 2794.600 ;
        RECT 2311.590 2794.320 2311.870 2794.600 ;
        RECT 2318.490 2794.320 2318.770 2794.600 ;
        RECT 2325.390 2794.320 2325.670 2794.600 ;
        RECT 2332.290 2794.320 2332.570 2794.600 ;
        RECT 2339.650 2794.320 2339.930 2794.600 ;
        RECT 2343.790 2794.320 2344.070 2794.600 ;
        RECT 2346.090 2794.320 2346.370 2794.600 ;
        RECT 2352.990 2794.320 2353.270 2794.600 ;
        RECT 2359.890 2794.320 2360.170 2794.600 ;
        RECT 2366.790 2794.320 2367.070 2794.600 ;
        RECT 2374.150 2794.320 2374.430 2794.600 ;
        RECT 2385.650 2794.320 2385.930 2794.600 ;
        RECT 2391.630 2794.320 2391.910 2794.600 ;
        RECT 2394.850 2794.320 2395.130 2794.600 ;
        RECT 2415.090 2794.320 2415.370 2794.600 ;
        RECT 2428.890 2794.320 2429.170 2794.600 ;
        RECT 2235.690 2788.880 2235.970 2789.160 ;
        RECT 2228.790 2787.520 2229.070 2787.800 ;
        RECT 2193.830 2087.120 2194.110 2087.400 ;
        RECT 2263.750 2793.640 2264.030 2793.920 ;
        RECT 2266.510 2792.960 2266.790 2793.240 ;
        RECT 2273.410 2793.640 2273.690 2793.920 ;
        RECT 2279.850 2793.640 2280.130 2793.920 ;
        RECT 2284.450 2793.640 2284.730 2793.920 ;
        RECT 2294.110 2792.960 2294.390 2793.240 ;
        RECT 2298.250 2793.640 2298.530 2793.920 ;
        RECT 2304.230 2793.640 2304.510 2793.920 ;
        RECT 2305.150 2793.640 2305.430 2793.920 ;
        RECT 2307.910 2790.920 2308.190 2791.200 ;
        RECT 2315.270 2793.640 2315.550 2793.920 ;
        RECT 2321.710 2793.640 2321.990 2793.920 ;
        RECT 2326.770 2793.640 2327.050 2793.920 ;
        RECT 2333.670 2793.640 2333.950 2793.920 ;
        RECT 2339.190 2793.640 2339.470 2793.920 ;
        RECT 2340.110 2792.960 2340.390 2793.240 ;
        RECT 2347.470 2793.640 2347.750 2793.920 ;
        RECT 2356.670 2793.640 2356.950 2793.920 ;
        RECT 2361.270 2793.640 2361.550 2793.920 ;
        RECT 2367.250 2793.640 2367.530 2793.920 ;
        RECT 2373.690 2792.960 2373.970 2793.240 ;
        RECT 2377.370 2793.640 2377.650 2793.920 ;
        RECT 2402.670 2793.640 2402.950 2793.920 ;
        RECT 2421.990 2793.640 2422.270 2793.920 ;
        RECT 2435.790 2793.640 2436.070 2793.920 ;
        RECT 2402.670 2792.960 2402.950 2793.240 ;
        RECT 2408.190 2792.960 2408.470 2793.240 ;
        RECT 2415.090 2792.960 2415.370 2793.240 ;
        RECT 2387.490 2791.600 2387.770 2791.880 ;
        RECT 2380.590 2790.240 2380.870 2790.520 ;
        RECT 2394.390 2790.240 2394.670 2790.520 ;
        RECT 2380.590 2789.560 2380.870 2789.840 ;
        RECT 2415.090 2792.280 2415.370 2792.560 ;
        RECT 2408.190 2790.920 2408.470 2791.200 ;
        RECT 2442.690 2792.960 2442.970 2793.240 ;
        RECT 2428.890 2791.600 2429.170 2791.880 ;
        RECT 2435.790 2791.600 2436.070 2791.880 ;
        RECT 2415.090 2788.880 2415.370 2789.160 ;
        RECT 2421.990 2788.200 2422.270 2788.480 ;
        RECT 1412.290 1622.000 1412.570 1622.280 ;
        RECT 1410.910 1617.240 1411.190 1617.520 ;
        RECT 1408.150 1611.800 1408.430 1612.080 ;
        RECT 1407.690 1607.040 1407.970 1607.320 ;
        RECT 1397.570 1603.640 1397.850 1603.920 ;
      LAYER met3 ;
        RECT 646.365 3264.500 646.695 3264.505 ;
        RECT 646.110 3264.490 646.695 3264.500 ;
        RECT 645.910 3264.190 646.695 3264.490 ;
        RECT 646.110 3264.180 646.695 3264.190 ;
        RECT 646.365 3264.175 646.695 3264.180 ;
        RECT 667.985 3264.500 668.315 3264.505 ;
        RECT 1293.125 3264.500 1293.455 3264.505 ;
        RECT 667.985 3264.490 668.570 3264.500 ;
        RECT 1292.870 3264.490 1293.455 3264.500 ;
        RECT 667.985 3264.190 668.770 3264.490 ;
        RECT 1292.670 3264.190 1293.455 3264.490 ;
        RECT 667.985 3264.180 668.570 3264.190 ;
        RECT 1292.870 3264.180 1293.455 3264.190 ;
        RECT 667.985 3264.175 668.315 3264.180 ;
        RECT 1293.125 3264.175 1293.455 3264.180 ;
        RECT 1890.665 3264.500 1890.995 3264.505 ;
        RECT 1917.805 3264.500 1918.135 3264.505 ;
        RECT 1890.665 3264.490 1891.250 3264.500 ;
        RECT 1917.550 3264.490 1918.135 3264.500 ;
        RECT 1890.665 3264.190 1891.450 3264.490 ;
        RECT 1917.350 3264.190 1918.135 3264.490 ;
        RECT 1890.665 3264.180 1891.250 3264.190 ;
        RECT 1917.550 3264.180 1918.135 3264.190 ;
        RECT 1890.665 3264.175 1890.995 3264.180 ;
        RECT 1917.805 3264.175 1918.135 3264.180 ;
        RECT 2542.025 3264.500 2542.355 3264.505 ;
        RECT 2566.865 3264.500 2567.195 3264.505 ;
        RECT 2542.025 3264.490 2542.610 3264.500 ;
        RECT 2566.865 3264.490 2567.450 3264.500 ;
        RECT 2542.025 3264.190 2542.810 3264.490 ;
        RECT 2566.865 3264.190 2567.650 3264.490 ;
        RECT 2542.025 3264.180 2542.610 3264.190 ;
        RECT 2566.865 3264.180 2567.450 3264.190 ;
        RECT 2542.025 3264.175 2542.355 3264.180 ;
        RECT 2566.865 3264.175 2567.195 3264.180 ;
        RECT 1317.505 3258.380 1317.835 3258.385 ;
        RECT 1317.505 3258.370 1318.205 3258.380 ;
        RECT 1317.505 3258.070 1318.290 3258.370 ;
        RECT 1317.505 3258.060 1318.205 3258.070 ;
        RECT 1317.505 3258.055 1317.835 3258.060 ;
        RECT 659.280 3251.235 661.020 3252.140 ;
        RECT 821.165 3251.570 821.495 3251.585 ;
        RECT 869.005 3251.570 869.335 3251.585 ;
        RECT 821.165 3251.270 869.335 3251.570 ;
        RECT 821.165 3251.255 821.495 3251.270 ;
        RECT 869.005 3251.255 869.335 3251.270 ;
        RECT 1309.280 3251.235 1311.020 3252.140 ;
        RECT 1909.280 3251.235 1911.020 3252.140 ;
        RECT 2559.280 3251.235 2561.020 3252.140 ;
        RECT 300.000 3232.785 304.600 3233.085 ;
        RECT 289.405 3230.490 289.735 3230.505 ;
        RECT 300.230 3230.490 300.530 3232.785 ;
        RECT 289.405 3230.190 300.530 3230.490 ;
        RECT 289.405 3230.175 289.735 3230.190 ;
        RECT 300.000 3227.145 304.600 3227.445 ;
        RECT 288.945 3225.050 289.275 3225.065 ;
        RECT 300.230 3225.050 300.530 3227.145 ;
        RECT 288.945 3224.750 300.530 3225.050 ;
        RECT 288.945 3224.735 289.275 3224.750 ;
        RECT 300.000 3218.645 304.600 3218.945 ;
        RECT 288.485 3216.210 288.815 3216.225 ;
        RECT 300.230 3216.210 300.530 3218.645 ;
        RECT 288.485 3215.910 300.530 3216.210 ;
        RECT 288.485 3215.895 288.815 3215.910 ;
        RECT 300.000 3213.005 304.600 3213.305 ;
        RECT 288.025 3210.090 288.355 3210.105 ;
        RECT 300.230 3210.090 300.530 3213.005 ;
        RECT 288.025 3209.790 300.530 3210.090 ;
        RECT 288.025 3209.775 288.355 3209.790 ;
        RECT 300.000 3204.505 304.600 3204.805 ;
        RECT 287.565 3201.930 287.895 3201.945 ;
        RECT 300.230 3201.930 300.530 3204.505 ;
        RECT 287.565 3201.630 300.530 3201.930 ;
        RECT 287.565 3201.615 287.895 3201.630 ;
        RECT 300.000 3198.865 304.600 3199.165 ;
        RECT 287.105 3196.490 287.435 3196.505 ;
        RECT 300.230 3196.490 300.530 3198.865 ;
        RECT 287.105 3196.190 300.530 3196.490 ;
        RECT 287.105 3196.175 287.435 3196.190 ;
        RECT 300.000 3190.365 304.600 3190.665 ;
        RECT 286.645 3188.330 286.975 3188.345 ;
        RECT 300.230 3188.330 300.530 3190.365 ;
        RECT 286.645 3188.030 300.530 3188.330 ;
        RECT 286.645 3188.015 286.975 3188.030 ;
        RECT 300.000 2901.125 304.600 2901.425 ;
        RECT 286.185 2898.650 286.515 2898.665 ;
        RECT 300.230 2898.650 300.530 2901.125 ;
        RECT 286.185 2898.350 300.530 2898.650 ;
        RECT 286.185 2898.335 286.515 2898.350 ;
        RECT 302.950 2894.940 303.330 2895.260 ;
        RECT 302.990 2892.925 303.290 2894.940 ;
        RECT 300.000 2892.625 304.600 2892.925 ;
      LAYER met3 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met3 ;
        RECT 688.225 3248.565 688.555 3248.580 ;
        RECT 681.880 3248.265 688.555 3248.565 ;
        RECT 688.225 3248.250 688.555 3248.265 ;
        RECT 950.000 3232.785 954.600 3233.085 ;
        RECT 941.685 3230.490 942.015 3230.505 ;
        RECT 950.670 3230.490 950.970 3232.785 ;
        RECT 941.685 3230.190 950.970 3230.490 ;
        RECT 941.685 3230.175 942.015 3230.190 ;
        RECT 950.000 3227.145 954.600 3227.445 ;
        RECT 942.145 3225.050 942.475 3225.065 ;
        RECT 950.670 3225.050 950.970 3227.145 ;
        RECT 942.145 3224.750 950.970 3225.050 ;
        RECT 942.145 3224.735 942.475 3224.750 ;
        RECT 950.000 3218.645 954.600 3218.945 ;
        RECT 942.605 3216.210 942.935 3216.225 ;
        RECT 950.670 3216.210 950.970 3218.645 ;
        RECT 942.605 3215.910 950.970 3216.210 ;
        RECT 942.605 3215.895 942.935 3215.910 ;
        RECT 950.000 3213.005 954.600 3213.305 ;
        RECT 943.065 3210.090 943.395 3210.105 ;
        RECT 950.670 3210.090 950.970 3213.005 ;
        RECT 943.065 3209.790 950.970 3210.090 ;
        RECT 943.065 3209.775 943.395 3209.790 ;
        RECT 950.000 3204.505 954.600 3204.805 ;
        RECT 943.525 3201.930 943.855 3201.945 ;
        RECT 950.670 3201.930 950.970 3204.505 ;
        RECT 943.525 3201.630 950.970 3201.930 ;
        RECT 943.525 3201.615 943.855 3201.630 ;
        RECT 950.000 3198.865 954.600 3199.165 ;
        RECT 943.985 3196.490 944.315 3196.505 ;
        RECT 950.670 3196.490 950.970 3198.865 ;
        RECT 943.985 3196.190 950.970 3196.490 ;
        RECT 943.985 3196.175 944.315 3196.190 ;
        RECT 950.000 3190.365 954.600 3190.665 ;
        RECT 944.445 3188.330 944.775 3188.345 ;
        RECT 950.670 3188.330 950.970 3190.365 ;
        RECT 944.445 3188.030 950.970 3188.330 ;
        RECT 944.445 3188.015 944.775 3188.030 ;
        RECT 696.965 2948.290 697.295 2948.305 ;
        RECT 684.790 2947.990 697.295 2948.290 ;
        RECT 684.790 2947.210 685.090 2947.990 ;
        RECT 696.965 2947.975 697.295 2947.990 ;
        RECT 681.880 2946.910 686.480 2947.210 ;
        RECT 684.790 2938.710 685.090 2946.910 ;
        RECT 681.880 2938.410 686.480 2938.710 ;
        RECT 684.790 2933.070 685.090 2938.410 ;
        RECT 681.880 2932.770 686.480 2933.070 ;
        RECT 685.710 2924.570 686.010 2932.770 ;
        RECT 681.880 2924.270 686.480 2924.570 ;
        RECT 685.710 2918.930 686.010 2924.270 ;
        RECT 681.880 2918.630 686.480 2918.930 ;
        RECT 685.710 2910.430 686.010 2918.630 ;
        RECT 681.880 2910.130 686.480 2910.430 ;
        RECT 685.710 2904.790 686.010 2910.130 ;
        RECT 681.880 2904.490 686.480 2904.790 ;
        RECT 950.000 2901.125 954.600 2901.425 ;
        RECT 939.385 2898.650 939.715 2898.665 ;
        RECT 950.670 2898.650 950.970 2901.125 ;
        RECT 939.385 2898.350 950.970 2898.650 ;
        RECT 939.385 2898.335 939.715 2898.350 ;
        RECT 944.190 2895.250 944.570 2895.260 ;
        RECT 944.190 2894.950 950.970 2895.250 ;
        RECT 944.190 2894.940 944.570 2894.950 ;
        RECT 950.670 2892.925 950.970 2894.950 ;
        RECT 950.000 2892.625 954.600 2892.925 ;
      LAYER met3 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met3 ;
        RECT 1332.225 3249.530 1332.555 3249.545 ;
        RECT 1332.225 3249.215 1332.770 3249.530 ;
        RECT 1332.470 3248.565 1332.770 3249.215 ;
        RECT 1331.880 3248.265 1336.480 3248.565 ;
        RECT 1550.000 3232.785 1554.600 3233.085 ;
        RECT 1536.925 3230.490 1537.255 3230.505 ;
        RECT 1550.510 3230.490 1550.810 3232.785 ;
        RECT 1536.925 3230.190 1550.810 3230.490 ;
        RECT 1536.925 3230.175 1537.255 3230.190 ;
        RECT 1550.000 3227.145 1554.600 3227.445 ;
        RECT 1535.545 3225.050 1535.875 3225.065 ;
        RECT 1550.510 3225.050 1550.810 3227.145 ;
        RECT 1535.545 3224.750 1550.810 3225.050 ;
        RECT 1535.545 3224.735 1535.875 3224.750 ;
        RECT 1550.000 3218.645 1554.600 3218.945 ;
        RECT 1535.545 3217.570 1535.875 3217.585 ;
        RECT 1550.510 3217.570 1550.810 3218.645 ;
        RECT 1535.545 3217.270 1550.810 3217.570 ;
        RECT 1535.545 3217.255 1535.875 3217.270 ;
        RECT 1550.000 3213.005 1554.600 3213.305 ;
        RECT 1538.305 3210.770 1538.635 3210.785 ;
        RECT 1550.510 3210.770 1550.810 3213.005 ;
        RECT 1538.305 3210.470 1550.810 3210.770 ;
        RECT 1538.305 3210.455 1538.635 3210.470 ;
        RECT 1550.000 3204.505 1554.600 3204.805 ;
        RECT 1538.305 3202.610 1538.635 3202.625 ;
        RECT 1550.510 3202.610 1550.810 3204.505 ;
        RECT 1538.305 3202.310 1550.810 3202.610 ;
        RECT 1538.305 3202.295 1538.635 3202.310 ;
        RECT 1550.000 3198.865 1554.600 3199.165 ;
        RECT 1533.245 3197.170 1533.575 3197.185 ;
        RECT 1550.510 3197.170 1550.810 3198.865 ;
        RECT 1533.245 3196.870 1550.810 3197.170 ;
        RECT 1533.245 3196.855 1533.575 3196.870 ;
        RECT 1550.000 3190.365 1554.600 3190.665 ;
        RECT 1534.165 3189.690 1534.495 3189.705 ;
        RECT 1550.510 3189.690 1550.810 3190.365 ;
        RECT 1534.165 3189.390 1550.810 3189.690 ;
        RECT 1534.165 3189.375 1534.495 3189.390 ;
        RECT 1331.880 2946.930 1336.480 2947.210 ;
        RECT 1345.565 2946.930 1345.895 2946.945 ;
        RECT 1331.880 2946.910 1345.895 2946.930 ;
        RECT 1336.150 2946.630 1345.895 2946.910 ;
        RECT 1345.565 2946.615 1345.895 2946.630 ;
        RECT 1331.880 2938.410 1336.480 2938.710 ;
        RECT 1336.150 2936.050 1336.450 2938.410 ;
        RECT 1345.565 2936.050 1345.895 2936.065 ;
        RECT 1351.750 2936.050 1352.130 2936.060 ;
        RECT 1336.150 2935.750 1352.130 2936.050 ;
        RECT 1336.150 2933.070 1336.450 2935.750 ;
        RECT 1345.565 2935.735 1345.895 2935.750 ;
        RECT 1351.750 2935.740 1352.130 2935.750 ;
        RECT 1331.880 2932.770 1336.480 2933.070 ;
        RECT 1336.150 2924.570 1336.450 2932.770 ;
        RECT 1331.880 2924.270 1336.480 2924.570 ;
        RECT 1336.150 2918.930 1336.450 2924.270 ;
        RECT 1331.880 2918.630 1336.480 2918.930 ;
        RECT 1336.150 2910.430 1336.450 2918.630 ;
        RECT 1331.880 2910.130 1336.480 2910.430 ;
        RECT 1336.150 2904.790 1336.450 2910.130 ;
        RECT 1331.880 2904.490 1336.480 2904.790 ;
        RECT 1336.150 2902.050 1336.450 2904.490 ;
        RECT 1352.005 2902.050 1352.335 2902.065 ;
        RECT 1336.150 2901.750 1352.335 2902.050 ;
        RECT 1352.005 2901.735 1352.335 2901.750 ;
        RECT 1550.000 2901.125 1554.600 2901.425 ;
        RECT 1538.305 2899.330 1538.635 2899.345 ;
        RECT 1550.510 2899.330 1550.810 2901.125 ;
        RECT 1538.305 2899.030 1550.810 2899.330 ;
        RECT 1538.305 2899.015 1538.635 2899.030 ;
        RECT 1408.125 2895.250 1408.455 2895.265 ;
        RECT 1412.470 2895.250 1412.850 2895.260 ;
        RECT 1408.125 2894.950 1412.850 2895.250 ;
        RECT 1408.125 2894.935 1408.455 2894.950 ;
        RECT 1412.470 2894.940 1412.850 2894.950 ;
        RECT 1551.390 2894.940 1551.770 2895.260 ;
        RECT 1551.430 2892.925 1551.730 2894.940 ;
        RECT 1550.000 2892.625 1554.600 2892.925 ;
      LAYER met3 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met3 ;
        RECT 1935.745 3249.530 1936.075 3249.545 ;
        RECT 1935.745 3249.215 1936.290 3249.530 ;
        RECT 1935.990 3248.565 1936.290 3249.215 ;
        RECT 1931.880 3248.265 1936.480 3248.565 ;
        RECT 2200.000 3232.785 2204.600 3233.085 ;
        RECT 2190.585 3230.490 2190.915 3230.505 ;
        RECT 2200.030 3230.490 2200.330 3232.785 ;
        RECT 2190.585 3230.190 2200.330 3230.490 ;
        RECT 2190.585 3230.175 2190.915 3230.190 ;
        RECT 2200.000 3227.145 2204.600 3227.445 ;
        RECT 2191.045 3225.050 2191.375 3225.065 ;
        RECT 2200.030 3225.050 2200.330 3227.145 ;
        RECT 2191.045 3224.750 2200.330 3225.050 ;
        RECT 2191.045 3224.735 2191.375 3224.750 ;
        RECT 2200.000 3218.645 2204.600 3218.945 ;
        RECT 2191.505 3216.210 2191.835 3216.225 ;
        RECT 2200.030 3216.210 2200.330 3218.645 ;
        RECT 2191.505 3215.910 2200.330 3216.210 ;
        RECT 2191.505 3215.895 2191.835 3215.910 ;
        RECT 2200.000 3213.005 2204.600 3213.305 ;
        RECT 2191.965 3210.090 2192.295 3210.105 ;
        RECT 2200.030 3210.090 2200.330 3213.005 ;
        RECT 2191.965 3209.790 2200.330 3210.090 ;
        RECT 2191.965 3209.775 2192.295 3209.790 ;
        RECT 2200.000 3204.505 2204.600 3204.805 ;
        RECT 2192.425 3201.930 2192.755 3201.945 ;
        RECT 2200.030 3201.930 2200.330 3204.505 ;
        RECT 2192.425 3201.630 2200.330 3201.930 ;
        RECT 2192.425 3201.615 2192.755 3201.630 ;
        RECT 2200.000 3198.865 2204.600 3199.165 ;
        RECT 2192.885 3196.490 2193.215 3196.505 ;
        RECT 2200.030 3196.490 2200.330 3198.865 ;
        RECT 2192.885 3196.190 2200.330 3196.490 ;
        RECT 2192.885 3196.175 2193.215 3196.190 ;
        RECT 2200.000 3190.365 2204.600 3190.665 ;
        RECT 2193.345 3188.330 2193.675 3188.345 ;
        RECT 2200.030 3188.330 2200.330 3190.365 ;
        RECT 2193.345 3188.030 2200.330 3188.330 ;
        RECT 2193.345 3188.015 2193.675 3188.030 ;
        RECT 1931.880 2946.910 1936.480 2947.210 ;
        RECT 1935.990 2938.710 1936.290 2946.910 ;
        RECT 1931.880 2938.410 1936.480 2938.710 ;
        RECT 1935.990 2936.050 1936.290 2938.410 ;
        RECT 1946.070 2936.050 1946.450 2936.060 ;
        RECT 1935.990 2935.750 1946.450 2936.050 ;
        RECT 1935.990 2933.070 1936.290 2935.750 ;
        RECT 1946.070 2935.740 1946.450 2935.750 ;
        RECT 1931.880 2932.770 1936.480 2933.070 ;
        RECT 1935.990 2924.570 1936.290 2932.770 ;
        RECT 1931.880 2924.270 1936.480 2924.570 ;
        RECT 1935.990 2918.930 1936.290 2924.270 ;
        RECT 1931.880 2918.630 1936.480 2918.930 ;
        RECT 1935.990 2910.430 1936.290 2918.630 ;
        RECT 1931.880 2910.130 1936.480 2910.430 ;
        RECT 1935.990 2904.790 1936.290 2910.130 ;
        RECT 1931.880 2904.490 1936.480 2904.790 ;
        RECT 2200.000 2901.125 2204.600 2901.425 ;
        RECT 2193.805 2898.650 2194.135 2898.665 ;
        RECT 2200.030 2898.650 2200.330 2901.125 ;
        RECT 2193.805 2898.350 2200.330 2898.650 ;
        RECT 2193.805 2898.335 2194.135 2898.350 ;
        RECT 2187.110 2895.250 2187.490 2895.260 ;
        RECT 2187.110 2894.950 2200.330 2895.250 ;
        RECT 2187.110 2894.940 2187.490 2894.950 ;
        RECT 2200.030 2892.925 2200.330 2894.950 ;
        RECT 2200.000 2892.625 2204.600 2892.925 ;
      LAYER met3 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met3 ;
        RECT 2582.045 3249.530 2582.375 3249.545 ;
        RECT 2582.045 3249.230 2583.050 3249.530 ;
        RECT 2582.045 3249.215 2582.375 3249.230 ;
        RECT 2582.750 3248.565 2583.050 3249.230 ;
        RECT 2581.880 3248.265 2586.480 3248.565 ;
        RECT 2581.880 2946.930 2586.480 2947.210 ;
        RECT 2594.465 2946.930 2594.795 2946.945 ;
        RECT 2581.880 2946.910 2594.795 2946.930 ;
        RECT 2585.510 2946.630 2594.795 2946.910 ;
        RECT 2594.465 2946.615 2594.795 2946.630 ;
        RECT 2594.465 2938.770 2594.795 2938.785 ;
        RECT 2585.510 2938.710 2594.795 2938.770 ;
        RECT 2581.880 2938.470 2594.795 2938.710 ;
        RECT 2581.880 2938.410 2586.480 2938.470 ;
        RECT 2594.465 2938.455 2594.795 2938.470 ;
        RECT 2585.510 2936.050 2585.810 2938.410 ;
        RECT 2587.310 2936.050 2587.690 2936.060 ;
        RECT 2585.510 2935.750 2587.690 2936.050 ;
        RECT 2585.510 2933.070 2585.810 2935.750 ;
        RECT 2587.310 2935.740 2587.690 2935.750 ;
        RECT 2581.880 2932.770 2586.480 2933.070 ;
        RECT 2585.510 2924.570 2585.810 2932.770 ;
        RECT 2581.880 2924.270 2586.480 2924.570 ;
        RECT 2585.510 2918.930 2585.810 2924.270 ;
        RECT 2581.880 2918.630 2586.480 2918.930 ;
        RECT 2585.510 2910.430 2585.810 2918.630 ;
        RECT 2581.880 2910.130 2586.480 2910.430 ;
        RECT 2585.510 2904.790 2585.810 2910.130 ;
        RECT 2581.880 2904.490 2586.480 2904.790 ;
        RECT 1054.845 2800.050 1055.175 2800.065 ;
        RECT 1055.510 2800.050 1055.890 2800.060 ;
        RECT 1054.845 2799.750 1055.890 2800.050 ;
        RECT 1054.845 2799.735 1055.175 2799.750 ;
        RECT 1055.510 2799.740 1055.890 2799.750 ;
        RECT 1794.830 2799.370 1795.210 2799.380 ;
        RECT 1794.830 2799.070 1796.450 2799.370 ;
        RECT 1794.830 2799.060 1795.210 2799.070 ;
        RECT 1795.190 2798.010 1795.570 2798.020 ;
        RECT 1796.150 2798.010 1796.450 2799.070 ;
        RECT 1795.190 2797.710 1796.450 2798.010 ;
        RECT 1795.190 2797.700 1795.570 2797.710 ;
        RECT 1053.005 2795.980 1053.335 2795.985 ;
        RECT 1732.885 2795.980 1733.215 2795.985 ;
        RECT 1052.750 2795.970 1053.335 2795.980 ;
        RECT 1732.630 2795.970 1733.215 2795.980 ;
        RECT 1052.550 2795.670 1053.335 2795.970 ;
        RECT 1732.430 2795.670 1733.215 2795.970 ;
        RECT 1052.750 2795.660 1053.335 2795.670 ;
        RECT 1732.630 2795.660 1733.215 2795.670 ;
        RECT 1053.005 2795.655 1053.335 2795.660 ;
        RECT 1732.885 2795.655 1733.215 2795.660 ;
        RECT 336.990 2794.610 337.370 2794.620 ;
        RECT 337.705 2794.610 338.035 2794.625 ;
        RECT 336.990 2794.310 338.035 2794.610 ;
        RECT 336.990 2794.300 337.370 2794.310 ;
        RECT 337.705 2794.295 338.035 2794.310 ;
        RECT 342.510 2794.610 342.890 2794.620 ;
        RECT 344.605 2794.610 344.935 2794.625 ;
        RECT 342.510 2794.310 344.935 2794.610 ;
        RECT 342.510 2794.300 342.890 2794.310 ;
        RECT 344.605 2794.295 344.935 2794.310 ;
        RECT 350.790 2794.610 351.170 2794.620 ;
        RECT 351.505 2794.610 351.835 2794.625 ;
        RECT 358.405 2794.620 358.735 2794.625 ;
        RECT 362.085 2794.620 362.415 2794.625 ;
        RECT 350.790 2794.310 351.835 2794.610 ;
        RECT 350.790 2794.300 351.170 2794.310 ;
        RECT 351.505 2794.295 351.835 2794.310 ;
        RECT 358.150 2794.610 358.735 2794.620 ;
        RECT 361.830 2794.610 362.415 2794.620 ;
        RECT 358.150 2794.310 358.960 2794.610 ;
        RECT 361.630 2794.310 362.415 2794.610 ;
        RECT 358.150 2794.300 358.735 2794.310 ;
        RECT 361.830 2794.300 362.415 2794.310 ;
        RECT 364.590 2794.610 364.970 2794.620 ;
        RECT 365.305 2794.610 365.635 2794.625 ;
        RECT 368.525 2794.620 368.855 2794.625 ;
        RECT 371.285 2794.620 371.615 2794.625 ;
        RECT 374.965 2794.620 375.295 2794.625 ;
        RECT 378.645 2794.620 378.975 2794.625 ;
        RECT 368.270 2794.610 368.855 2794.620 ;
        RECT 371.030 2794.610 371.615 2794.620 ;
        RECT 374.710 2794.610 375.295 2794.620 ;
        RECT 378.390 2794.610 378.975 2794.620 ;
        RECT 364.590 2794.310 365.635 2794.610 ;
        RECT 368.070 2794.310 368.855 2794.610 ;
        RECT 370.830 2794.310 371.615 2794.610 ;
        RECT 374.510 2794.310 375.295 2794.610 ;
        RECT 378.190 2794.310 378.975 2794.610 ;
        RECT 364.590 2794.300 364.970 2794.310 ;
        RECT 358.405 2794.295 358.735 2794.300 ;
        RECT 362.085 2794.295 362.415 2794.300 ;
        RECT 365.305 2794.295 365.635 2794.310 ;
        RECT 368.270 2794.300 368.855 2794.310 ;
        RECT 371.030 2794.300 371.615 2794.310 ;
        RECT 374.710 2794.300 375.295 2794.310 ;
        RECT 378.390 2794.300 378.975 2794.310 ;
        RECT 379.310 2794.610 379.690 2794.620 ;
        RECT 380.025 2794.610 380.355 2794.625 ;
        RECT 379.310 2794.310 380.355 2794.610 ;
        RECT 379.310 2794.300 379.690 2794.310 ;
        RECT 368.525 2794.295 368.855 2794.300 ;
        RECT 371.285 2794.295 371.615 2794.300 ;
        RECT 374.965 2794.295 375.295 2794.300 ;
        RECT 378.645 2794.295 378.975 2794.300 ;
        RECT 380.025 2794.295 380.355 2794.310 ;
        RECT 383.910 2794.610 384.290 2794.620 ;
        RECT 384.625 2794.610 384.955 2794.625 ;
        RECT 386.925 2794.620 387.255 2794.625 ;
        RECT 390.605 2794.620 390.935 2794.625 ;
        RECT 392.445 2794.620 392.775 2794.625 ;
        RECT 386.670 2794.610 387.255 2794.620 ;
        RECT 390.350 2794.610 390.935 2794.620 ;
        RECT 392.190 2794.610 392.775 2794.620 ;
        RECT 383.910 2794.310 384.955 2794.610 ;
        RECT 386.470 2794.310 387.255 2794.610 ;
        RECT 390.150 2794.310 390.935 2794.610 ;
        RECT 391.990 2794.310 392.775 2794.610 ;
        RECT 383.910 2794.300 384.290 2794.310 ;
        RECT 384.625 2794.295 384.955 2794.310 ;
        RECT 386.670 2794.300 387.255 2794.310 ;
        RECT 390.350 2794.300 390.935 2794.310 ;
        RECT 392.190 2794.300 392.775 2794.310 ;
        RECT 395.870 2794.610 396.250 2794.620 ;
        RECT 396.585 2794.610 396.915 2794.625 ;
        RECT 399.805 2794.620 400.135 2794.625 ;
        RECT 399.550 2794.610 400.135 2794.620 ;
        RECT 395.870 2794.310 396.915 2794.610 ;
        RECT 399.350 2794.310 400.135 2794.610 ;
        RECT 395.870 2794.300 396.250 2794.310 ;
        RECT 386.925 2794.295 387.255 2794.300 ;
        RECT 390.605 2794.295 390.935 2794.300 ;
        RECT 392.445 2794.295 392.775 2794.300 ;
        RECT 396.585 2794.295 396.915 2794.310 ;
        RECT 399.550 2794.300 400.135 2794.310 ;
        RECT 403.230 2794.610 403.610 2794.620 ;
        RECT 403.945 2794.610 404.275 2794.625 ;
        RECT 406.245 2794.620 406.575 2794.625 ;
        RECT 409.925 2794.620 410.255 2794.625 ;
        RECT 413.605 2794.620 413.935 2794.625 ;
        RECT 414.525 2794.620 414.855 2794.625 ;
        RECT 405.990 2794.610 406.575 2794.620 ;
        RECT 409.670 2794.610 410.255 2794.620 ;
        RECT 413.350 2794.610 413.935 2794.620 ;
        RECT 403.230 2794.310 404.275 2794.610 ;
        RECT 405.790 2794.310 406.575 2794.610 ;
        RECT 409.470 2794.310 410.255 2794.610 ;
        RECT 413.150 2794.310 413.935 2794.610 ;
        RECT 403.230 2794.300 403.610 2794.310 ;
        RECT 399.805 2794.295 400.135 2794.300 ;
        RECT 403.945 2794.295 404.275 2794.310 ;
        RECT 405.990 2794.300 406.575 2794.310 ;
        RECT 409.670 2794.300 410.255 2794.310 ;
        RECT 413.350 2794.300 413.935 2794.310 ;
        RECT 414.270 2794.610 414.855 2794.620 ;
        RECT 417.950 2794.610 418.330 2794.620 ;
        RECT 418.665 2794.610 418.995 2794.625 ;
        RECT 420.965 2794.620 421.295 2794.625 ;
        RECT 414.270 2794.310 415.080 2794.610 ;
        RECT 417.950 2794.310 418.995 2794.610 ;
        RECT 414.270 2794.300 414.855 2794.310 ;
        RECT 417.950 2794.300 418.330 2794.310 ;
        RECT 406.245 2794.295 406.575 2794.300 ;
        RECT 409.925 2794.295 410.255 2794.300 ;
        RECT 413.605 2794.295 413.935 2794.300 ;
        RECT 414.525 2794.295 414.855 2794.300 ;
        RECT 418.665 2794.295 418.995 2794.310 ;
        RECT 420.710 2794.610 421.295 2794.620 ;
        RECT 425.310 2794.610 425.690 2794.620 ;
        RECT 427.405 2794.610 427.735 2794.625 ;
        RECT 432.005 2794.620 432.335 2794.625 ;
        RECT 431.750 2794.610 432.335 2794.620 ;
        RECT 420.710 2794.310 421.520 2794.610 ;
        RECT 425.310 2794.310 427.735 2794.610 ;
        RECT 431.550 2794.310 432.335 2794.610 ;
        RECT 420.710 2794.300 421.295 2794.310 ;
        RECT 425.310 2794.300 425.690 2794.310 ;
        RECT 420.965 2794.295 421.295 2794.300 ;
        RECT 427.405 2794.295 427.735 2794.310 ;
        RECT 431.750 2794.300 432.335 2794.310 ;
        RECT 433.590 2794.610 433.970 2794.620 ;
        RECT 434.305 2794.610 434.635 2794.625 ;
        RECT 439.365 2794.620 439.695 2794.625 ;
        RECT 441.205 2794.620 441.535 2794.625 ;
        RECT 439.110 2794.610 439.695 2794.620 ;
        RECT 433.590 2794.310 434.635 2794.610 ;
        RECT 438.910 2794.310 439.695 2794.610 ;
        RECT 433.590 2794.300 433.970 2794.310 ;
        RECT 432.005 2794.295 432.335 2794.300 ;
        RECT 434.305 2794.295 434.635 2794.310 ;
        RECT 439.110 2794.300 439.695 2794.310 ;
        RECT 440.950 2794.610 441.535 2794.620 ;
        RECT 444.425 2794.620 444.755 2794.625 ;
        RECT 444.425 2794.610 445.010 2794.620 ;
        RECT 440.950 2794.310 441.760 2794.610 ;
        RECT 444.200 2794.310 445.010 2794.610 ;
        RECT 440.950 2794.300 441.535 2794.310 ;
        RECT 439.365 2794.295 439.695 2794.300 ;
        RECT 441.205 2794.295 441.535 2794.300 ;
        RECT 444.425 2794.300 445.010 2794.310 ;
        RECT 445.550 2794.610 445.930 2794.620 ;
        RECT 448.105 2794.610 448.435 2794.625 ;
        RECT 450.405 2794.620 450.735 2794.625 ;
        RECT 455.005 2794.620 455.335 2794.625 ;
        RECT 450.150 2794.610 450.735 2794.620 ;
        RECT 445.550 2794.310 448.435 2794.610 ;
        RECT 449.950 2794.310 450.735 2794.610 ;
        RECT 445.550 2794.300 445.930 2794.310 ;
        RECT 444.425 2794.295 444.755 2794.300 ;
        RECT 448.105 2794.295 448.435 2794.310 ;
        RECT 450.150 2794.300 450.735 2794.310 ;
        RECT 454.750 2794.610 455.335 2794.620 ;
        RECT 460.270 2794.610 460.650 2794.620 ;
        RECT 461.905 2794.610 462.235 2794.625 ;
        RECT 454.750 2794.310 455.560 2794.610 ;
        RECT 460.270 2794.310 462.235 2794.610 ;
        RECT 454.750 2794.300 455.335 2794.310 ;
        RECT 460.270 2794.300 460.650 2794.310 ;
        RECT 450.405 2794.295 450.735 2794.300 ;
        RECT 455.005 2794.295 455.335 2794.300 ;
        RECT 461.905 2794.295 462.235 2794.310 ;
        RECT 466.505 2794.620 466.835 2794.625 ;
        RECT 468.345 2794.620 468.675 2794.625 ;
        RECT 466.505 2794.610 467.090 2794.620 ;
        RECT 468.345 2794.610 468.930 2794.620 ;
        RECT 466.505 2794.310 467.290 2794.610 ;
        RECT 468.120 2794.310 468.930 2794.610 ;
        RECT 466.505 2794.300 467.090 2794.310 ;
        RECT 468.345 2794.300 468.930 2794.310 ;
        RECT 474.990 2794.610 475.370 2794.620 ;
        RECT 475.705 2794.610 476.035 2794.625 ;
        RECT 474.990 2794.310 476.035 2794.610 ;
        RECT 474.990 2794.300 475.370 2794.310 ;
        RECT 466.505 2794.295 466.835 2794.300 ;
        RECT 468.345 2794.295 468.675 2794.300 ;
        RECT 475.705 2794.295 476.035 2794.310 ;
        RECT 478.465 2794.620 478.795 2794.625 ;
        RECT 482.605 2794.620 482.935 2794.625 ;
        RECT 478.465 2794.610 479.050 2794.620 ;
        RECT 482.350 2794.610 482.935 2794.620 ;
        RECT 484.905 2794.620 485.235 2794.625 ;
        RECT 489.045 2794.620 489.375 2794.625 ;
        RECT 484.905 2794.610 485.490 2794.620 ;
        RECT 488.790 2794.610 489.375 2794.620 ;
        RECT 478.465 2794.310 479.250 2794.610 ;
        RECT 482.350 2794.310 483.160 2794.610 ;
        RECT 484.905 2794.310 485.690 2794.610 ;
        RECT 488.590 2794.310 489.375 2794.610 ;
        RECT 478.465 2794.300 479.050 2794.310 ;
        RECT 482.350 2794.300 482.935 2794.310 ;
        RECT 478.465 2794.295 478.795 2794.300 ;
        RECT 482.605 2794.295 482.935 2794.300 ;
        RECT 484.905 2794.300 485.490 2794.310 ;
        RECT 488.790 2794.300 489.375 2794.310 ;
        RECT 491.550 2794.610 491.930 2794.620 ;
        RECT 492.725 2794.610 493.055 2794.625 ;
        RECT 491.550 2794.310 493.055 2794.610 ;
        RECT 491.550 2794.300 491.930 2794.310 ;
        RECT 484.905 2794.295 485.235 2794.300 ;
        RECT 489.045 2794.295 489.375 2794.300 ;
        RECT 492.725 2794.295 493.055 2794.310 ;
        RECT 495.230 2794.610 495.610 2794.620 ;
        RECT 496.405 2794.610 496.735 2794.625 ;
        RECT 495.230 2794.310 496.735 2794.610 ;
        RECT 495.230 2794.300 495.610 2794.310 ;
        RECT 496.405 2794.295 496.735 2794.310 ;
        RECT 500.750 2794.610 501.130 2794.620 ;
        RECT 501.925 2794.610 502.255 2794.625 ;
        RECT 500.750 2794.310 502.255 2794.610 ;
        RECT 500.750 2794.300 501.130 2794.310 ;
        RECT 501.925 2794.295 502.255 2794.310 ;
        RECT 507.190 2794.610 507.570 2794.620 ;
        RECT 509.745 2794.610 510.075 2794.625 ;
        RECT 513.885 2794.620 514.215 2794.625 ;
        RECT 513.630 2794.610 514.215 2794.620 ;
        RECT 507.190 2794.310 510.075 2794.610 ;
        RECT 513.430 2794.310 514.215 2794.610 ;
        RECT 507.190 2794.300 507.570 2794.310 ;
        RECT 509.745 2794.295 510.075 2794.310 ;
        RECT 513.630 2794.300 514.215 2794.310 ;
        RECT 516.390 2794.610 516.770 2794.620 ;
        RECT 517.105 2794.610 517.435 2794.625 ;
        RECT 524.005 2794.620 524.335 2794.625 ;
        RECT 526.765 2794.620 527.095 2794.625 ;
        RECT 523.750 2794.610 524.335 2794.620 ;
        RECT 526.510 2794.610 527.095 2794.620 ;
        RECT 516.390 2794.310 517.435 2794.610 ;
        RECT 523.550 2794.310 524.335 2794.610 ;
        RECT 526.310 2794.310 527.095 2794.610 ;
        RECT 516.390 2794.300 516.770 2794.310 ;
        RECT 513.885 2794.295 514.215 2794.300 ;
        RECT 517.105 2794.295 517.435 2794.310 ;
        RECT 523.750 2794.300 524.335 2794.310 ;
        RECT 526.510 2794.300 527.095 2794.310 ;
        RECT 530.190 2794.610 530.570 2794.620 ;
        RECT 530.905 2794.610 531.235 2794.625 ;
        RECT 530.190 2794.310 531.235 2794.610 ;
        RECT 530.190 2794.300 530.570 2794.310 ;
        RECT 524.005 2794.295 524.335 2794.300 ;
        RECT 526.765 2794.295 527.095 2794.300 ;
        RECT 530.905 2794.295 531.235 2794.310 ;
        RECT 535.710 2794.610 536.090 2794.620 ;
        RECT 537.345 2794.610 537.675 2794.625 ;
        RECT 535.710 2794.310 537.675 2794.610 ;
        RECT 535.710 2794.300 536.090 2794.310 ;
        RECT 537.345 2794.295 537.675 2794.310 ;
        RECT 538.470 2794.610 538.850 2794.620 ;
        RECT 539.185 2794.610 539.515 2794.625 ;
        RECT 538.470 2794.310 539.515 2794.610 ;
        RECT 538.470 2794.300 538.850 2794.310 ;
        RECT 539.185 2794.295 539.515 2794.310 ;
        RECT 542.150 2794.610 542.530 2794.620 ;
        RECT 544.245 2794.610 544.575 2794.625 ;
        RECT 542.150 2794.310 544.575 2794.610 ;
        RECT 542.150 2794.300 542.530 2794.310 ;
        RECT 544.245 2794.295 544.575 2794.310 ;
        RECT 547.670 2794.610 548.050 2794.620 ;
        RECT 551.605 2794.610 551.935 2794.625 ;
        RECT 547.670 2794.310 551.935 2794.610 ;
        RECT 547.670 2794.300 548.050 2794.310 ;
        RECT 551.605 2794.295 551.935 2794.310 ;
        RECT 979.865 2794.610 980.195 2794.625 ;
        RECT 980.990 2794.610 981.370 2794.620 ;
        RECT 979.865 2794.310 981.370 2794.610 ;
        RECT 979.865 2794.295 980.195 2794.310 ;
        RECT 980.990 2794.300 981.370 2794.310 ;
        RECT 1013.190 2794.610 1013.570 2794.620 ;
        RECT 1013.905 2794.610 1014.235 2794.625 ;
        RECT 1018.965 2794.620 1019.295 2794.625 ;
        RECT 1018.710 2794.610 1019.295 2794.620 ;
        RECT 1013.190 2794.310 1014.235 2794.610 ;
        RECT 1018.510 2794.310 1019.295 2794.610 ;
        RECT 1013.190 2794.300 1013.570 2794.310 ;
        RECT 1013.905 2794.295 1014.235 2794.310 ;
        RECT 1018.710 2794.300 1019.295 2794.310 ;
        RECT 1019.630 2794.610 1020.010 2794.620 ;
        RECT 1020.805 2794.610 1021.135 2794.625 ;
        RECT 1019.630 2794.310 1021.135 2794.610 ;
        RECT 1019.630 2794.300 1020.010 2794.310 ;
        RECT 1018.965 2794.295 1019.295 2794.300 ;
        RECT 1020.805 2794.295 1021.135 2794.310 ;
        RECT 1026.990 2794.610 1027.370 2794.620 ;
        RECT 1027.705 2794.610 1028.035 2794.625 ;
        RECT 1026.990 2794.310 1028.035 2794.610 ;
        RECT 1026.990 2794.300 1027.370 2794.310 ;
        RECT 1027.705 2794.295 1028.035 2794.310 ;
        RECT 1030.670 2794.610 1031.050 2794.620 ;
        RECT 1034.605 2794.610 1034.935 2794.625 ;
        RECT 1030.670 2794.310 1034.935 2794.610 ;
        RECT 1030.670 2794.300 1031.050 2794.310 ;
        RECT 1034.605 2794.295 1034.935 2794.310 ;
        RECT 1041.710 2794.610 1042.090 2794.620 ;
        RECT 1042.425 2794.610 1042.755 2794.625 ;
        RECT 1041.710 2794.310 1042.755 2794.610 ;
        RECT 1041.710 2794.300 1042.090 2794.310 ;
        RECT 1042.425 2794.295 1042.755 2794.310 ;
        RECT 1058.985 2794.620 1059.315 2794.625 ;
        RECT 1065.425 2794.620 1065.755 2794.625 ;
        RECT 1058.985 2794.610 1059.570 2794.620 ;
        RECT 1065.425 2794.610 1066.010 2794.620 ;
        RECT 1069.565 2794.610 1069.895 2794.625 ;
        RECT 1070.230 2794.610 1070.610 2794.620 ;
        RECT 1058.985 2794.310 1059.770 2794.610 ;
        RECT 1065.425 2794.310 1066.210 2794.610 ;
        RECT 1069.565 2794.310 1070.610 2794.610 ;
        RECT 1058.985 2794.300 1059.570 2794.310 ;
        RECT 1065.425 2794.300 1066.010 2794.310 ;
        RECT 1058.985 2794.295 1059.315 2794.300 ;
        RECT 1065.425 2794.295 1065.755 2794.300 ;
        RECT 1069.565 2794.295 1069.895 2794.310 ;
        RECT 1070.230 2794.300 1070.610 2794.310 ;
        RECT 1081.270 2794.610 1081.650 2794.620 ;
        RECT 1082.905 2794.610 1083.235 2794.625 ;
        RECT 1081.270 2794.310 1083.235 2794.610 ;
        RECT 1081.270 2794.300 1081.650 2794.310 ;
        RECT 1082.905 2794.295 1083.235 2794.310 ;
        RECT 1087.505 2794.620 1087.835 2794.625 ;
        RECT 1089.805 2794.620 1090.135 2794.625 ;
        RECT 1094.405 2794.620 1094.735 2794.625 ;
        RECT 1087.505 2794.610 1088.090 2794.620 ;
        RECT 1089.550 2794.610 1090.135 2794.620 ;
        RECT 1094.150 2794.610 1094.735 2794.620 ;
        RECT 1087.505 2794.310 1088.290 2794.610 ;
        RECT 1089.550 2794.310 1090.360 2794.610 ;
        RECT 1093.950 2794.310 1094.735 2794.610 ;
        RECT 1087.505 2794.300 1088.090 2794.310 ;
        RECT 1089.550 2794.300 1090.135 2794.310 ;
        RECT 1094.150 2794.300 1094.735 2794.310 ;
        RECT 1095.990 2794.610 1096.370 2794.620 ;
        RECT 1096.705 2794.610 1097.035 2794.625 ;
        RECT 1100.845 2794.620 1101.175 2794.625 ;
        RECT 1103.605 2794.620 1103.935 2794.625 ;
        RECT 1105.445 2794.620 1105.775 2794.625 ;
        RECT 1100.590 2794.610 1101.175 2794.620 ;
        RECT 1095.990 2794.310 1097.035 2794.610 ;
        RECT 1100.390 2794.310 1101.175 2794.610 ;
        RECT 1095.990 2794.300 1096.370 2794.310 ;
        RECT 1087.505 2794.295 1087.835 2794.300 ;
        RECT 1089.805 2794.295 1090.135 2794.300 ;
        RECT 1094.405 2794.295 1094.735 2794.300 ;
        RECT 1096.705 2794.295 1097.035 2794.310 ;
        RECT 1100.590 2794.300 1101.175 2794.310 ;
        RECT 1103.350 2794.610 1103.935 2794.620 ;
        RECT 1105.190 2794.610 1105.775 2794.620 ;
        RECT 1103.350 2794.310 1104.160 2794.610 ;
        RECT 1104.990 2794.310 1105.775 2794.610 ;
        RECT 1103.350 2794.300 1103.935 2794.310 ;
        RECT 1105.190 2794.300 1105.775 2794.310 ;
        RECT 1109.790 2794.610 1110.170 2794.620 ;
        RECT 1110.505 2794.610 1110.835 2794.625 ;
        RECT 1109.790 2794.310 1110.835 2794.610 ;
        RECT 1109.790 2794.300 1110.170 2794.310 ;
        RECT 1100.845 2794.295 1101.175 2794.300 ;
        RECT 1103.605 2794.295 1103.935 2794.300 ;
        RECT 1105.445 2794.295 1105.775 2794.300 ;
        RECT 1110.505 2794.295 1110.835 2794.310 ;
        RECT 1111.425 2794.620 1111.755 2794.625 ;
        RECT 1118.325 2794.620 1118.655 2794.625 ;
        RECT 1111.425 2794.610 1112.010 2794.620 ;
        RECT 1118.070 2794.610 1118.655 2794.620 ;
        RECT 1111.425 2794.310 1112.210 2794.610 ;
        RECT 1117.870 2794.310 1118.655 2794.610 ;
        RECT 1111.425 2794.300 1112.010 2794.310 ;
        RECT 1118.070 2794.300 1118.655 2794.310 ;
        RECT 1121.750 2794.610 1122.130 2794.620 ;
        RECT 1124.305 2794.610 1124.635 2794.625 ;
        RECT 1129.365 2794.620 1129.695 2794.625 ;
        RECT 1131.205 2794.620 1131.535 2794.625 ;
        RECT 1135.805 2794.620 1136.135 2794.625 ;
        RECT 1129.110 2794.610 1129.695 2794.620 ;
        RECT 1121.750 2794.310 1124.635 2794.610 ;
        RECT 1128.910 2794.310 1129.695 2794.610 ;
        RECT 1121.750 2794.300 1122.130 2794.310 ;
        RECT 1111.425 2794.295 1111.755 2794.300 ;
        RECT 1118.325 2794.295 1118.655 2794.300 ;
        RECT 1124.305 2794.295 1124.635 2794.310 ;
        RECT 1129.110 2794.300 1129.695 2794.310 ;
        RECT 1130.950 2794.610 1131.535 2794.620 ;
        RECT 1135.550 2794.610 1136.135 2794.620 ;
        RECT 1130.950 2794.310 1131.760 2794.610 ;
        RECT 1135.350 2794.310 1136.135 2794.610 ;
        RECT 1130.950 2794.300 1131.535 2794.310 ;
        RECT 1135.550 2794.300 1136.135 2794.310 ;
        RECT 1137.390 2794.610 1137.770 2794.620 ;
        RECT 1138.105 2794.610 1138.435 2794.625 ;
        RECT 1137.390 2794.310 1138.435 2794.610 ;
        RECT 1137.390 2794.300 1137.770 2794.310 ;
        RECT 1129.365 2794.295 1129.695 2794.300 ;
        RECT 1131.205 2794.295 1131.535 2794.300 ;
        RECT 1135.805 2794.295 1136.135 2794.300 ;
        RECT 1138.105 2794.295 1138.435 2794.310 ;
        RECT 1139.945 2794.620 1140.275 2794.625 ;
        RECT 1139.945 2794.610 1140.530 2794.620 ;
        RECT 1143.830 2794.610 1144.210 2794.620 ;
        RECT 1145.005 2794.610 1145.335 2794.625 ;
        RECT 1139.945 2794.310 1140.730 2794.610 ;
        RECT 1143.830 2794.310 1145.335 2794.610 ;
        RECT 1139.945 2794.300 1140.530 2794.310 ;
        RECT 1143.830 2794.300 1144.210 2794.310 ;
        RECT 1139.945 2794.295 1140.275 2794.300 ;
        RECT 1145.005 2794.295 1145.335 2794.310 ;
        RECT 1146.385 2794.620 1146.715 2794.625 ;
        RECT 1146.385 2794.610 1146.970 2794.620 ;
        RECT 1151.190 2794.610 1151.570 2794.620 ;
        RECT 1151.905 2794.610 1152.235 2794.625 ;
        RECT 1146.385 2794.310 1147.170 2794.610 ;
        RECT 1151.190 2794.310 1152.235 2794.610 ;
        RECT 1146.385 2794.300 1146.970 2794.310 ;
        RECT 1151.190 2794.300 1151.570 2794.310 ;
        RECT 1146.385 2794.295 1146.715 2794.300 ;
        RECT 1151.905 2794.295 1152.235 2794.310 ;
        RECT 1153.950 2794.610 1154.330 2794.620 ;
        RECT 1158.805 2794.610 1159.135 2794.625 ;
        RECT 1165.245 2794.620 1165.575 2794.625 ;
        RECT 1172.605 2794.620 1172.935 2794.625 ;
        RECT 1153.950 2794.310 1159.135 2794.610 ;
        RECT 1153.950 2794.300 1154.330 2794.310 ;
        RECT 1158.805 2794.295 1159.135 2794.310 ;
        RECT 1164.990 2794.610 1165.575 2794.620 ;
        RECT 1172.350 2794.610 1172.935 2794.620 ;
        RECT 1178.790 2794.610 1179.170 2794.620 ;
        RECT 1179.505 2794.610 1179.835 2794.625 ;
        RECT 1186.405 2794.620 1186.735 2794.625 ;
        RECT 1164.990 2794.310 1165.800 2794.610 ;
        RECT 1172.350 2794.310 1173.160 2794.610 ;
        RECT 1178.790 2794.310 1179.835 2794.610 ;
        RECT 1164.990 2794.300 1165.575 2794.310 ;
        RECT 1172.350 2794.300 1172.935 2794.310 ;
        RECT 1178.790 2794.300 1179.170 2794.310 ;
        RECT 1165.245 2794.295 1165.575 2794.300 ;
        RECT 1172.605 2794.295 1172.935 2794.300 ;
        RECT 1179.505 2794.295 1179.835 2794.310 ;
        RECT 1186.150 2794.610 1186.735 2794.620 ;
        RECT 1198.110 2794.610 1198.490 2794.620 ;
        RECT 1200.205 2794.610 1200.535 2794.625 ;
        RECT 1613.285 2794.620 1613.615 2794.625 ;
        RECT 1642.725 2794.620 1643.055 2794.625 ;
        RECT 1652.845 2794.620 1653.175 2794.625 ;
        RECT 1659.285 2794.620 1659.615 2794.625 ;
        RECT 1613.030 2794.610 1613.615 2794.620 ;
        RECT 1642.470 2794.610 1643.055 2794.620 ;
        RECT 1652.590 2794.610 1653.175 2794.620 ;
        RECT 1659.030 2794.610 1659.615 2794.620 ;
        RECT 1186.150 2794.310 1186.960 2794.610 ;
        RECT 1198.110 2794.310 1200.535 2794.610 ;
        RECT 1612.830 2794.310 1613.615 2794.610 ;
        RECT 1642.270 2794.310 1643.055 2794.610 ;
        RECT 1652.390 2794.310 1653.175 2794.610 ;
        RECT 1658.830 2794.310 1659.615 2794.610 ;
        RECT 1186.150 2794.300 1186.735 2794.310 ;
        RECT 1198.110 2794.300 1198.490 2794.310 ;
        RECT 1186.405 2794.295 1186.735 2794.300 ;
        RECT 1200.205 2794.295 1200.535 2794.310 ;
        RECT 1613.030 2794.300 1613.615 2794.310 ;
        RECT 1642.470 2794.300 1643.055 2794.310 ;
        RECT 1652.590 2794.300 1653.175 2794.310 ;
        RECT 1659.030 2794.300 1659.615 2794.310 ;
        RECT 1665.470 2794.610 1665.850 2794.620 ;
        RECT 1669.405 2794.610 1669.735 2794.625 ;
        RECT 1670.325 2794.620 1670.655 2794.625 ;
        RECT 1665.470 2794.310 1669.735 2794.610 ;
        RECT 1665.470 2794.300 1665.850 2794.310 ;
        RECT 1613.285 2794.295 1613.615 2794.300 ;
        RECT 1642.725 2794.295 1643.055 2794.300 ;
        RECT 1652.845 2794.295 1653.175 2794.300 ;
        RECT 1659.285 2794.295 1659.615 2794.300 ;
        RECT 1669.405 2794.295 1669.735 2794.310 ;
        RECT 1670.070 2794.610 1670.655 2794.620 ;
        RECT 1677.225 2794.620 1677.555 2794.625 ;
        RECT 1695.165 2794.620 1695.495 2794.625 ;
        RECT 1677.225 2794.610 1677.810 2794.620 ;
        RECT 1694.910 2794.610 1695.495 2794.620 ;
        RECT 1670.070 2794.310 1670.880 2794.610 ;
        RECT 1677.225 2794.310 1678.010 2794.610 ;
        RECT 1694.710 2794.310 1695.495 2794.610 ;
        RECT 1670.070 2794.300 1670.655 2794.310 ;
        RECT 1670.325 2794.295 1670.655 2794.300 ;
        RECT 1677.225 2794.300 1677.810 2794.310 ;
        RECT 1694.910 2794.300 1695.495 2794.310 ;
        RECT 1677.225 2794.295 1677.555 2794.300 ;
        RECT 1695.165 2794.295 1695.495 2794.300 ;
        RECT 1699.305 2794.620 1699.635 2794.625 ;
        RECT 1706.205 2794.620 1706.535 2794.625 ;
        RECT 1712.645 2794.620 1712.975 2794.625 ;
        RECT 1718.165 2794.620 1718.495 2794.625 ;
        RECT 1723.685 2794.620 1724.015 2794.625 ;
        RECT 1699.305 2794.610 1699.890 2794.620 ;
        RECT 1705.950 2794.610 1706.535 2794.620 ;
        RECT 1712.390 2794.610 1712.975 2794.620 ;
        RECT 1717.910 2794.610 1718.495 2794.620 ;
        RECT 1723.430 2794.610 1724.015 2794.620 ;
        RECT 1699.305 2794.310 1700.090 2794.610 ;
        RECT 1705.750 2794.310 1706.535 2794.610 ;
        RECT 1712.190 2794.310 1712.975 2794.610 ;
        RECT 1717.710 2794.310 1718.495 2794.610 ;
        RECT 1723.230 2794.310 1724.015 2794.610 ;
        RECT 1699.305 2794.300 1699.890 2794.310 ;
        RECT 1705.950 2794.300 1706.535 2794.310 ;
        RECT 1712.390 2794.300 1712.975 2794.310 ;
        RECT 1717.910 2794.300 1718.495 2794.310 ;
        RECT 1723.430 2794.300 1724.015 2794.310 ;
        RECT 1699.305 2794.295 1699.635 2794.300 ;
        RECT 1706.205 2794.295 1706.535 2794.300 ;
        RECT 1712.645 2794.295 1712.975 2794.300 ;
        RECT 1718.165 2794.295 1718.495 2794.300 ;
        RECT 1723.685 2794.295 1724.015 2794.300 ;
        RECT 1728.745 2794.620 1729.075 2794.625 ;
        RECT 1741.165 2794.620 1741.495 2794.625 ;
        RECT 1747.605 2794.620 1747.935 2794.625 ;
        RECT 1728.745 2794.610 1729.330 2794.620 ;
        RECT 1740.910 2794.610 1741.495 2794.620 ;
        RECT 1747.350 2794.610 1747.935 2794.620 ;
        RECT 1728.745 2794.310 1729.530 2794.610 ;
        RECT 1740.710 2794.310 1741.495 2794.610 ;
        RECT 1747.150 2794.310 1747.935 2794.610 ;
        RECT 1728.745 2794.300 1729.330 2794.310 ;
        RECT 1740.910 2794.300 1741.495 2794.310 ;
        RECT 1747.350 2794.300 1747.935 2794.310 ;
        RECT 1728.745 2794.295 1729.075 2794.300 ;
        RECT 1741.165 2794.295 1741.495 2794.300 ;
        RECT 1747.605 2794.295 1747.935 2794.300 ;
        RECT 1760.025 2794.610 1760.355 2794.625 ;
        RECT 1762.070 2794.610 1762.450 2794.620 ;
        RECT 1760.025 2794.310 1762.450 2794.610 ;
        RECT 1760.025 2794.295 1760.355 2794.310 ;
        RECT 1762.070 2794.300 1762.450 2794.310 ;
        RECT 2242.565 2794.610 2242.895 2794.625 ;
        RECT 2243.230 2794.610 2243.610 2794.620 ;
        RECT 2242.565 2794.310 2243.610 2794.610 ;
        RECT 2242.565 2794.295 2242.895 2794.310 ;
        RECT 2243.230 2794.300 2243.610 2794.310 ;
        RECT 2256.365 2794.610 2256.695 2794.625 ;
        RECT 2257.030 2794.610 2257.410 2794.620 ;
        RECT 2256.365 2794.310 2257.410 2794.610 ;
        RECT 2256.365 2794.295 2256.695 2794.310 ;
        RECT 2257.030 2794.300 2257.410 2794.310 ;
        RECT 2263.265 2794.610 2263.595 2794.625 ;
        RECT 2268.325 2794.620 2268.655 2794.625 ;
        RECT 2264.390 2794.610 2264.770 2794.620 ;
        RECT 2268.070 2794.610 2268.655 2794.620 ;
        RECT 2263.265 2794.310 2264.770 2794.610 ;
        RECT 2267.870 2794.310 2268.655 2794.610 ;
        RECT 2263.265 2794.295 2263.595 2794.310 ;
        RECT 2264.390 2794.300 2264.770 2794.310 ;
        RECT 2268.070 2794.300 2268.655 2794.310 ;
        RECT 2268.325 2794.295 2268.655 2794.300 ;
        RECT 2270.165 2794.610 2270.495 2794.625 ;
        RECT 2276.350 2794.610 2276.730 2794.620 ;
        RECT 2270.165 2794.310 2276.730 2794.610 ;
        RECT 2270.165 2794.295 2270.495 2794.310 ;
        RECT 2276.350 2794.300 2276.730 2794.310 ;
        RECT 2277.065 2794.610 2277.395 2794.625 ;
        RECT 2282.790 2794.610 2283.170 2794.620 ;
        RECT 2277.065 2794.310 2283.170 2794.610 ;
        RECT 2277.065 2794.295 2277.395 2794.310 ;
        RECT 2282.790 2794.300 2283.170 2794.310 ;
        RECT 2283.965 2794.610 2284.295 2794.625 ;
        RECT 2287.390 2794.610 2287.770 2794.620 ;
        RECT 2283.965 2794.310 2287.770 2794.610 ;
        RECT 2283.965 2794.295 2284.295 2794.310 ;
        RECT 2287.390 2794.300 2287.770 2794.310 ;
        RECT 2290.865 2794.610 2291.195 2794.625 ;
        RECT 2293.830 2794.610 2294.210 2794.620 ;
        RECT 2290.865 2794.310 2294.210 2794.610 ;
        RECT 2290.865 2794.295 2291.195 2794.310 ;
        RECT 2293.830 2794.300 2294.210 2794.310 ;
        RECT 2297.765 2794.610 2298.095 2794.625 ;
        RECT 2304.665 2794.620 2304.995 2794.625 ;
        RECT 2308.805 2794.620 2309.135 2794.625 ;
        RECT 2300.270 2794.610 2300.650 2794.620 ;
        RECT 2297.765 2794.310 2300.650 2794.610 ;
        RECT 2297.765 2794.295 2298.095 2794.310 ;
        RECT 2300.270 2794.300 2300.650 2794.310 ;
        RECT 2304.665 2794.610 2305.250 2794.620 ;
        RECT 2308.550 2794.610 2309.135 2794.620 ;
        RECT 2304.665 2794.310 2305.450 2794.610 ;
        RECT 2308.350 2794.310 2309.135 2794.610 ;
        RECT 2304.665 2794.300 2305.250 2794.310 ;
        RECT 2308.550 2794.300 2309.135 2794.310 ;
        RECT 2304.665 2794.295 2304.995 2794.300 ;
        RECT 2308.805 2794.295 2309.135 2794.300 ;
        RECT 2311.565 2794.610 2311.895 2794.625 ;
        RECT 2316.830 2794.610 2317.210 2794.620 ;
        RECT 2311.565 2794.310 2317.210 2794.610 ;
        RECT 2311.565 2794.295 2311.895 2794.310 ;
        RECT 2316.830 2794.300 2317.210 2794.310 ;
        RECT 2318.465 2794.610 2318.795 2794.625 ;
        RECT 2322.350 2794.610 2322.730 2794.620 ;
        RECT 2318.465 2794.310 2322.730 2794.610 ;
        RECT 2318.465 2794.295 2318.795 2794.310 ;
        RECT 2322.350 2794.300 2322.730 2794.310 ;
        RECT 2325.365 2794.610 2325.695 2794.625 ;
        RECT 2328.790 2794.610 2329.170 2794.620 ;
        RECT 2325.365 2794.310 2329.170 2794.610 ;
        RECT 2325.365 2794.295 2325.695 2794.310 ;
        RECT 2328.790 2794.300 2329.170 2794.310 ;
        RECT 2332.265 2794.610 2332.595 2794.625 ;
        RECT 2339.625 2794.620 2339.955 2794.625 ;
        RECT 2343.765 2794.620 2344.095 2794.625 ;
        RECT 2334.310 2794.610 2334.690 2794.620 ;
        RECT 2339.625 2794.610 2340.210 2794.620 ;
        RECT 2343.510 2794.610 2344.095 2794.620 ;
        RECT 2332.265 2794.310 2334.690 2794.610 ;
        RECT 2339.400 2794.310 2340.210 2794.610 ;
        RECT 2343.310 2794.310 2344.095 2794.610 ;
        RECT 2332.265 2794.295 2332.595 2794.310 ;
        RECT 2334.310 2794.300 2334.690 2794.310 ;
        RECT 2339.625 2794.300 2340.210 2794.310 ;
        RECT 2343.510 2794.300 2344.095 2794.310 ;
        RECT 2339.625 2794.295 2339.955 2794.300 ;
        RECT 2343.765 2794.295 2344.095 2794.300 ;
        RECT 2346.065 2794.610 2346.395 2794.625 ;
        RECT 2351.790 2794.610 2352.170 2794.620 ;
        RECT 2346.065 2794.310 2352.170 2794.610 ;
        RECT 2346.065 2794.295 2346.395 2794.310 ;
        RECT 2351.790 2794.300 2352.170 2794.310 ;
        RECT 2352.965 2794.610 2353.295 2794.625 ;
        RECT 2357.310 2794.610 2357.690 2794.620 ;
        RECT 2352.965 2794.310 2357.690 2794.610 ;
        RECT 2352.965 2794.295 2353.295 2794.310 ;
        RECT 2357.310 2794.300 2357.690 2794.310 ;
        RECT 2359.865 2794.610 2360.195 2794.625 ;
        RECT 2363.750 2794.610 2364.130 2794.620 ;
        RECT 2359.865 2794.310 2364.130 2794.610 ;
        RECT 2359.865 2794.295 2360.195 2794.310 ;
        RECT 2363.750 2794.300 2364.130 2794.310 ;
        RECT 2366.765 2794.610 2367.095 2794.625 ;
        RECT 2374.125 2794.620 2374.455 2794.625 ;
        RECT 2370.190 2794.610 2370.570 2794.620 ;
        RECT 2373.870 2794.610 2374.455 2794.620 ;
        RECT 2366.765 2794.310 2370.570 2794.610 ;
        RECT 2373.670 2794.310 2374.455 2794.610 ;
        RECT 2366.765 2794.295 2367.095 2794.310 ;
        RECT 2370.190 2794.300 2370.570 2794.310 ;
        RECT 2373.870 2794.300 2374.455 2794.310 ;
        RECT 2374.125 2794.295 2374.455 2794.300 ;
        RECT 2385.625 2794.620 2385.955 2794.625 ;
        RECT 2391.605 2794.620 2391.935 2794.625 ;
        RECT 2385.625 2794.610 2386.210 2794.620 ;
        RECT 2391.350 2794.610 2391.935 2794.620 ;
        RECT 2385.625 2794.310 2386.410 2794.610 ;
        RECT 2391.150 2794.310 2391.935 2794.610 ;
        RECT 2385.625 2794.300 2386.210 2794.310 ;
        RECT 2391.350 2794.300 2391.935 2794.310 ;
        RECT 2385.625 2794.295 2385.955 2794.300 ;
        RECT 2391.605 2794.295 2391.935 2794.300 ;
        RECT 2394.825 2794.620 2395.155 2794.625 ;
        RECT 2394.825 2794.610 2395.410 2794.620 ;
        RECT 2415.065 2794.610 2415.395 2794.625 ;
        RECT 2420.790 2794.610 2421.170 2794.620 ;
        RECT 2394.825 2794.310 2395.610 2794.610 ;
        RECT 2415.065 2794.310 2421.170 2794.610 ;
        RECT 2394.825 2794.300 2395.410 2794.310 ;
        RECT 2394.825 2794.295 2395.155 2794.300 ;
        RECT 2415.065 2794.295 2415.395 2794.310 ;
        RECT 2420.790 2794.300 2421.170 2794.310 ;
        RECT 2428.865 2794.610 2429.195 2794.625 ;
        RECT 2429.990 2794.610 2430.370 2794.620 ;
        RECT 2428.865 2794.310 2430.370 2794.610 ;
        RECT 2428.865 2794.295 2429.195 2794.310 ;
        RECT 2429.990 2794.300 2430.370 2794.310 ;
        RECT 397.045 2793.940 397.375 2793.945 ;
        RECT 396.790 2793.930 397.375 2793.940 ;
        RECT 396.590 2793.630 397.375 2793.930 ;
        RECT 396.790 2793.620 397.375 2793.630 ;
        RECT 397.045 2793.615 397.375 2793.620 ;
        RECT 426.945 2793.940 427.275 2793.945 ;
        RECT 426.945 2793.930 427.530 2793.940 ;
        RECT 430.830 2793.930 431.210 2793.940 ;
        RECT 433.845 2793.930 434.175 2793.945 ;
        RECT 426.945 2793.630 427.730 2793.930 ;
        RECT 430.830 2793.630 434.175 2793.930 ;
        RECT 426.945 2793.620 427.530 2793.630 ;
        RECT 430.830 2793.620 431.210 2793.630 ;
        RECT 426.945 2793.615 427.275 2793.620 ;
        RECT 433.845 2793.615 434.175 2793.630 ;
        RECT 455.465 2793.940 455.795 2793.945 ;
        RECT 462.365 2793.940 462.695 2793.945 ;
        RECT 455.465 2793.930 456.050 2793.940 ;
        RECT 462.110 2793.930 462.695 2793.940 ;
        RECT 455.465 2793.630 456.250 2793.930 ;
        RECT 461.910 2793.630 462.695 2793.930 ;
        RECT 455.465 2793.620 456.050 2793.630 ;
        RECT 462.110 2793.620 462.695 2793.630 ;
        RECT 465.790 2793.930 466.170 2793.940 ;
        RECT 468.805 2793.930 469.135 2793.945 ;
        RECT 465.790 2793.630 469.135 2793.930 ;
        RECT 465.790 2793.620 466.170 2793.630 ;
        RECT 455.465 2793.615 455.795 2793.620 ;
        RECT 462.365 2793.615 462.695 2793.620 ;
        RECT 468.805 2793.615 469.135 2793.630 ;
        RECT 474.070 2793.930 474.450 2793.940 ;
        RECT 475.245 2793.930 475.575 2793.945 ;
        RECT 474.070 2793.630 475.575 2793.930 ;
        RECT 474.070 2793.620 474.450 2793.630 ;
        RECT 475.245 2793.615 475.575 2793.630 ;
        RECT 497.990 2793.930 498.370 2793.940 ;
        RECT 501.005 2793.930 501.335 2793.945 ;
        RECT 508.825 2793.940 509.155 2793.945 ;
        RECT 510.205 2793.940 510.535 2793.945 ;
        RECT 508.825 2793.930 509.410 2793.940 ;
        RECT 509.950 2793.930 510.535 2793.940 ;
        RECT 497.990 2793.630 501.335 2793.930 ;
        RECT 508.600 2793.630 509.410 2793.930 ;
        RECT 509.750 2793.630 510.535 2793.930 ;
        RECT 497.990 2793.620 498.370 2793.630 ;
        RECT 501.005 2793.615 501.335 2793.630 ;
        RECT 508.825 2793.620 509.410 2793.630 ;
        RECT 509.950 2793.620 510.535 2793.630 ;
        RECT 531.110 2793.930 531.490 2793.940 ;
        RECT 534.585 2793.930 534.915 2793.945 ;
        RECT 531.110 2793.630 534.915 2793.930 ;
        RECT 531.110 2793.620 531.490 2793.630 ;
        RECT 508.825 2793.615 509.155 2793.620 ;
        RECT 510.205 2793.615 510.535 2793.620 ;
        RECT 534.585 2793.615 534.915 2793.630 ;
        RECT 986.765 2793.930 987.095 2793.945 ;
        RECT 1001.025 2793.940 1001.355 2793.945 ;
        RECT 1076.465 2793.940 1076.795 2793.945 ;
        RECT 1083.365 2793.940 1083.695 2793.945 ;
        RECT 987.430 2793.930 987.810 2793.940 ;
        RECT 1001.025 2793.930 1001.610 2793.940 ;
        RECT 986.765 2793.630 987.810 2793.930 ;
        RECT 1000.800 2793.630 1001.610 2793.930 ;
        RECT 986.765 2793.615 987.095 2793.630 ;
        RECT 987.430 2793.620 987.810 2793.630 ;
        RECT 1001.025 2793.620 1001.610 2793.630 ;
        RECT 1076.465 2793.930 1077.050 2793.940 ;
        RECT 1083.110 2793.930 1083.695 2793.940 ;
        RECT 1076.465 2793.630 1077.250 2793.930 ;
        RECT 1082.910 2793.630 1083.695 2793.930 ;
        RECT 1076.465 2793.620 1077.050 2793.630 ;
        RECT 1083.110 2793.620 1083.695 2793.630 ;
        RECT 1086.790 2793.930 1087.170 2793.940 ;
        RECT 1089.345 2793.930 1089.675 2793.945 ;
        RECT 1086.790 2793.630 1089.675 2793.930 ;
        RECT 1086.790 2793.620 1087.170 2793.630 ;
        RECT 1001.025 2793.615 1001.355 2793.620 ;
        RECT 1076.465 2793.615 1076.795 2793.620 ;
        RECT 1083.365 2793.615 1083.695 2793.620 ;
        RECT 1089.345 2793.615 1089.675 2793.630 ;
        RECT 1122.005 2793.930 1122.335 2793.945 ;
        RECT 1122.670 2793.930 1123.050 2793.940 ;
        RECT 1122.005 2793.630 1123.050 2793.930 ;
        RECT 1122.005 2793.615 1122.335 2793.630 ;
        RECT 1122.670 2793.620 1123.050 2793.630 ;
        RECT 1128.190 2793.930 1128.570 2793.940 ;
        RECT 1130.745 2793.930 1131.075 2793.945 ;
        RECT 1128.190 2793.630 1131.075 2793.930 ;
        RECT 1128.190 2793.620 1128.570 2793.630 ;
        RECT 1130.745 2793.615 1131.075 2793.630 ;
        RECT 1163.150 2793.930 1163.530 2793.940 ;
        RECT 1165.705 2793.930 1166.035 2793.945 ;
        RECT 1173.065 2793.940 1173.395 2793.945 ;
        RECT 1173.065 2793.930 1173.650 2793.940 ;
        RECT 1163.150 2793.630 1166.035 2793.930 ;
        RECT 1172.840 2793.630 1173.650 2793.930 ;
        RECT 1163.150 2793.620 1163.530 2793.630 ;
        RECT 1165.705 2793.615 1166.035 2793.630 ;
        RECT 1173.065 2793.620 1173.650 2793.630 ;
        RECT 1179.965 2793.930 1180.295 2793.945 ;
        RECT 1186.865 2793.940 1187.195 2793.945 ;
        RECT 1688.725 2793.940 1689.055 2793.945 ;
        RECT 1180.630 2793.930 1181.010 2793.940 ;
        RECT 1186.865 2793.930 1187.450 2793.940 ;
        RECT 1688.470 2793.930 1689.055 2793.940 ;
        RECT 1179.965 2793.630 1181.010 2793.930 ;
        RECT 1186.640 2793.630 1187.450 2793.930 ;
        RECT 1688.270 2793.630 1689.055 2793.930 ;
        RECT 1173.065 2793.615 1173.395 2793.620 ;
        RECT 1179.965 2793.615 1180.295 2793.630 ;
        RECT 1180.630 2793.620 1181.010 2793.630 ;
        RECT 1186.865 2793.620 1187.450 2793.630 ;
        RECT 1688.470 2793.620 1689.055 2793.630 ;
        RECT 1186.865 2793.615 1187.195 2793.620 ;
        RECT 1688.725 2793.615 1689.055 2793.620 ;
        RECT 1766.465 2793.930 1766.795 2793.945 ;
        RECT 1780.265 2793.940 1780.595 2793.945 ;
        RECT 1767.590 2793.930 1767.970 2793.940 ;
        RECT 1780.265 2793.930 1780.850 2793.940 ;
        RECT 1766.465 2793.630 1767.970 2793.930 ;
        RECT 1780.040 2793.630 1780.850 2793.930 ;
        RECT 1766.465 2793.615 1766.795 2793.630 ;
        RECT 1767.590 2793.620 1767.970 2793.630 ;
        RECT 1780.265 2793.620 1780.850 2793.630 ;
        RECT 2263.725 2793.930 2264.055 2793.945 ;
        RECT 2273.385 2793.940 2273.715 2793.945 ;
        RECT 2279.825 2793.940 2280.155 2793.945 ;
        RECT 2284.425 2793.940 2284.755 2793.945 ;
        RECT 2268.990 2793.930 2269.370 2793.940 ;
        RECT 2263.725 2793.630 2269.370 2793.930 ;
        RECT 1780.265 2793.615 1780.595 2793.620 ;
        RECT 2263.725 2793.615 2264.055 2793.630 ;
        RECT 2268.990 2793.620 2269.370 2793.630 ;
        RECT 2273.385 2793.930 2273.970 2793.940 ;
        RECT 2279.825 2793.930 2280.410 2793.940 ;
        RECT 2284.425 2793.930 2285.010 2793.940 ;
        RECT 2297.510 2793.930 2297.890 2793.940 ;
        RECT 2298.225 2793.930 2298.555 2793.945 ;
        RECT 2304.205 2793.940 2304.535 2793.945 ;
        RECT 2303.950 2793.930 2304.535 2793.940 ;
        RECT 2273.385 2793.630 2274.170 2793.930 ;
        RECT 2279.825 2793.630 2280.610 2793.930 ;
        RECT 2284.425 2793.630 2285.210 2793.930 ;
        RECT 2297.510 2793.630 2298.555 2793.930 ;
        RECT 2303.750 2793.630 2304.535 2793.930 ;
        RECT 2273.385 2793.620 2273.970 2793.630 ;
        RECT 2279.825 2793.620 2280.410 2793.630 ;
        RECT 2284.425 2793.620 2285.010 2793.630 ;
        RECT 2297.510 2793.620 2297.890 2793.630 ;
        RECT 2273.385 2793.615 2273.715 2793.620 ;
        RECT 2279.825 2793.615 2280.155 2793.620 ;
        RECT 2284.425 2793.615 2284.755 2793.620 ;
        RECT 2298.225 2793.615 2298.555 2793.630 ;
        RECT 2303.950 2793.620 2304.535 2793.630 ;
        RECT 2304.205 2793.615 2304.535 2793.620 ;
        RECT 2305.125 2793.930 2305.455 2793.945 ;
        RECT 2315.245 2793.940 2315.575 2793.945 ;
        RECT 2321.685 2793.940 2322.015 2793.945 ;
        RECT 2310.390 2793.930 2310.770 2793.940 ;
        RECT 2314.990 2793.930 2315.575 2793.940 ;
        RECT 2321.430 2793.930 2322.015 2793.940 ;
        RECT 2305.125 2793.630 2310.770 2793.930 ;
        RECT 2314.790 2793.630 2315.575 2793.930 ;
        RECT 2321.230 2793.630 2322.015 2793.930 ;
        RECT 2305.125 2793.615 2305.455 2793.630 ;
        RECT 2310.390 2793.620 2310.770 2793.630 ;
        RECT 2314.990 2793.620 2315.575 2793.630 ;
        RECT 2321.430 2793.620 2322.015 2793.630 ;
        RECT 2326.030 2793.930 2326.410 2793.940 ;
        RECT 2326.745 2793.930 2327.075 2793.945 ;
        RECT 2326.030 2793.630 2327.075 2793.930 ;
        RECT 2326.030 2793.620 2326.410 2793.630 ;
        RECT 2315.245 2793.615 2315.575 2793.620 ;
        RECT 2321.685 2793.615 2322.015 2793.620 ;
        RECT 2326.745 2793.615 2327.075 2793.630 ;
        RECT 2332.470 2793.930 2332.850 2793.940 ;
        RECT 2333.645 2793.930 2333.975 2793.945 ;
        RECT 2332.470 2793.630 2333.975 2793.930 ;
        RECT 2332.470 2793.620 2332.850 2793.630 ;
        RECT 2333.645 2793.615 2333.975 2793.630 ;
        RECT 2339.165 2793.930 2339.495 2793.945 ;
        RECT 2345.350 2793.930 2345.730 2793.940 ;
        RECT 2339.165 2793.630 2345.730 2793.930 ;
        RECT 2339.165 2793.615 2339.495 2793.630 ;
        RECT 2345.350 2793.620 2345.730 2793.630 ;
        RECT 2347.445 2793.930 2347.775 2793.945 ;
        RECT 2356.645 2793.940 2356.975 2793.945 ;
        RECT 2361.245 2793.940 2361.575 2793.945 ;
        RECT 2348.110 2793.930 2348.490 2793.940 ;
        RECT 2356.390 2793.930 2356.975 2793.940 ;
        RECT 2360.990 2793.930 2361.575 2793.940 ;
        RECT 2347.445 2793.630 2348.490 2793.930 ;
        RECT 2356.190 2793.630 2356.975 2793.930 ;
        RECT 2360.790 2793.630 2361.575 2793.930 ;
        RECT 2347.445 2793.615 2347.775 2793.630 ;
        RECT 2348.110 2793.620 2348.490 2793.630 ;
        RECT 2356.390 2793.620 2356.975 2793.630 ;
        RECT 2360.990 2793.620 2361.575 2793.630 ;
        RECT 2356.645 2793.615 2356.975 2793.620 ;
        RECT 2361.245 2793.615 2361.575 2793.620 ;
        RECT 2367.225 2793.940 2367.555 2793.945 ;
        RECT 2377.345 2793.940 2377.675 2793.945 ;
        RECT 2367.225 2793.930 2367.810 2793.940 ;
        RECT 2377.345 2793.930 2377.930 2793.940 ;
        RECT 2402.645 2793.930 2402.975 2793.945 ;
        RECT 2403.310 2793.930 2403.690 2793.940 ;
        RECT 2367.225 2793.630 2368.010 2793.930 ;
        RECT 2377.345 2793.630 2378.130 2793.930 ;
        RECT 2402.645 2793.630 2403.690 2793.930 ;
        RECT 2367.225 2793.620 2367.810 2793.630 ;
        RECT 2377.345 2793.620 2377.930 2793.630 ;
        RECT 2367.225 2793.615 2367.555 2793.620 ;
        RECT 2377.345 2793.615 2377.675 2793.620 ;
        RECT 2402.645 2793.615 2402.975 2793.630 ;
        RECT 2403.310 2793.620 2403.690 2793.630 ;
        RECT 2421.965 2793.930 2422.295 2793.945 ;
        RECT 2423.550 2793.930 2423.930 2793.940 ;
        RECT 2421.965 2793.630 2423.930 2793.930 ;
        RECT 2421.965 2793.615 2422.295 2793.630 ;
        RECT 2423.550 2793.620 2423.930 2793.630 ;
        RECT 2435.765 2793.930 2436.095 2793.945 ;
        RECT 2436.430 2793.930 2436.810 2793.940 ;
        RECT 2435.765 2793.630 2436.810 2793.930 ;
        RECT 2435.765 2793.615 2436.095 2793.630 ;
        RECT 2436.430 2793.620 2436.810 2793.630 ;
        RECT 500.085 2793.250 500.415 2793.265 ;
        RECT 501.670 2793.250 502.050 2793.260 ;
        RECT 500.085 2792.950 502.050 2793.250 ;
        RECT 500.085 2792.935 500.415 2792.950 ;
        RECT 501.670 2792.940 502.050 2792.950 ;
        RECT 520.070 2793.250 520.450 2793.260 ;
        RECT 520.785 2793.250 521.115 2793.265 ;
        RECT 520.070 2792.950 521.115 2793.250 ;
        RECT 520.070 2792.940 520.450 2792.950 ;
        RECT 520.785 2792.935 521.115 2792.950 ;
        RECT 541.485 2793.250 541.815 2793.265 ;
        RECT 543.070 2793.250 543.450 2793.260 ;
        RECT 541.485 2792.950 543.450 2793.250 ;
        RECT 541.485 2792.935 541.815 2792.950 ;
        RECT 543.070 2792.940 543.450 2792.950 ;
        RECT 1010.685 2793.250 1011.015 2793.265 ;
        RECT 1024.485 2793.260 1024.815 2793.265 ;
        RECT 1012.270 2793.250 1012.650 2793.260 ;
        RECT 1024.230 2793.250 1024.815 2793.260 ;
        RECT 1010.685 2792.950 1012.650 2793.250 ;
        RECT 1024.030 2792.950 1024.815 2793.250 ;
        RECT 1010.685 2792.935 1011.015 2792.950 ;
        RECT 1012.270 2792.940 1012.650 2792.950 ;
        RECT 1024.230 2792.940 1024.815 2792.950 ;
        RECT 1024.485 2792.935 1024.815 2792.940 ;
        RECT 1045.185 2793.250 1045.515 2793.265 ;
        RECT 1048.150 2793.250 1048.530 2793.260 ;
        RECT 1045.185 2792.950 1048.530 2793.250 ;
        RECT 1045.185 2792.935 1045.515 2792.950 ;
        RECT 1048.150 2792.940 1048.530 2792.950 ;
        RECT 1166.165 2793.250 1166.495 2793.265 ;
        RECT 1636.745 2793.260 1637.075 2793.265 ;
        RECT 1167.750 2793.250 1168.130 2793.260 ;
        RECT 1166.165 2792.950 1168.130 2793.250 ;
        RECT 1166.165 2792.935 1166.495 2792.950 ;
        RECT 1167.750 2792.940 1168.130 2792.950 ;
        RECT 1636.745 2793.250 1637.330 2793.260 ;
        RECT 1681.110 2793.250 1681.490 2793.260 ;
        RECT 1682.285 2793.250 1682.615 2793.265 ;
        RECT 1636.745 2792.950 1682.615 2793.250 ;
        RECT 1636.745 2792.940 1637.330 2792.950 ;
        RECT 1681.110 2792.940 1681.490 2792.950 ;
        RECT 1636.745 2792.935 1637.075 2792.940 ;
        RECT 1682.285 2792.935 1682.615 2792.950 ;
        RECT 1787.165 2793.250 1787.495 2793.265 ;
        RECT 1787.830 2793.250 1788.210 2793.260 ;
        RECT 1787.165 2792.950 1788.210 2793.250 ;
        RECT 1787.165 2792.935 1787.495 2792.950 ;
        RECT 1787.830 2792.940 1788.210 2792.950 ;
        RECT 2263.470 2793.250 2263.850 2793.260 ;
        RECT 2266.485 2793.250 2266.815 2793.265 ;
        RECT 2263.470 2792.950 2266.815 2793.250 ;
        RECT 2263.470 2792.940 2263.850 2792.950 ;
        RECT 2266.485 2792.935 2266.815 2792.950 ;
        RECT 2291.990 2793.250 2292.370 2793.260 ;
        RECT 2294.085 2793.250 2294.415 2793.265 ;
        RECT 2291.990 2792.950 2294.415 2793.250 ;
        RECT 2291.990 2792.940 2292.370 2792.950 ;
        RECT 2294.085 2792.935 2294.415 2792.950 ;
        RECT 2338.910 2793.250 2339.290 2793.260 ;
        RECT 2340.085 2793.250 2340.415 2793.265 ;
        RECT 2338.910 2792.950 2340.415 2793.250 ;
        RECT 2338.910 2792.940 2339.290 2792.950 ;
        RECT 2340.085 2792.935 2340.415 2792.950 ;
        RECT 2373.665 2793.250 2373.995 2793.265 ;
        RECT 2374.790 2793.250 2375.170 2793.260 ;
        RECT 2373.665 2792.950 2375.170 2793.250 ;
        RECT 2373.665 2792.935 2373.995 2792.950 ;
        RECT 2374.790 2792.940 2375.170 2792.950 ;
        RECT 2402.645 2793.250 2402.975 2793.265 ;
        RECT 2408.165 2793.260 2408.495 2793.265 ;
        RECT 2404.230 2793.250 2404.610 2793.260 ;
        RECT 2402.645 2792.950 2404.610 2793.250 ;
        RECT 2402.645 2792.935 2402.975 2792.950 ;
        RECT 2404.230 2792.940 2404.610 2792.950 ;
        RECT 2407.910 2793.250 2408.495 2793.260 ;
        RECT 2415.065 2793.260 2415.395 2793.265 ;
        RECT 2442.665 2793.260 2442.995 2793.265 ;
        RECT 2415.065 2793.250 2415.650 2793.260 ;
        RECT 2442.665 2793.250 2443.250 2793.260 ;
        RECT 2407.910 2792.950 2408.720 2793.250 ;
        RECT 2414.840 2792.950 2415.650 2793.250 ;
        RECT 2442.440 2792.950 2443.250 2793.250 ;
        RECT 2407.910 2792.940 2408.495 2792.950 ;
        RECT 2408.165 2792.935 2408.495 2792.940 ;
        RECT 2415.065 2792.940 2415.650 2792.950 ;
        RECT 2442.665 2792.940 2443.250 2792.950 ;
        RECT 2415.065 2792.935 2415.395 2792.940 ;
        RECT 2442.665 2792.935 2442.995 2792.940 ;
        RECT 348.950 2792.570 349.330 2792.580 ;
        RECT 351.045 2792.570 351.375 2792.585 ;
        RECT 348.950 2792.270 351.375 2792.570 ;
        RECT 348.950 2792.260 349.330 2792.270 ;
        RECT 351.045 2792.255 351.375 2792.270 ;
        RECT 1116.230 2792.570 1116.610 2792.580 ;
        RECT 1117.405 2792.570 1117.735 2792.585 ;
        RECT 1116.230 2792.270 1117.735 2792.570 ;
        RECT 1116.230 2792.260 1116.610 2792.270 ;
        RECT 1117.405 2792.255 1117.735 2792.270 ;
        RECT 1152.365 2792.570 1152.695 2792.585 ;
        RECT 1153.030 2792.570 1153.410 2792.580 ;
        RECT 1152.365 2792.270 1153.410 2792.570 ;
        RECT 1152.365 2792.255 1152.695 2792.270 ;
        RECT 1153.030 2792.260 1153.410 2792.270 ;
        RECT 1596.265 2792.570 1596.595 2792.585 ;
        RECT 1752.665 2792.580 1752.995 2792.585 ;
        RECT 1637.870 2792.570 1638.250 2792.580 ;
        RECT 1596.265 2792.270 1638.250 2792.570 ;
        RECT 1596.265 2792.255 1596.595 2792.270 ;
        RECT 1637.870 2792.260 1638.250 2792.270 ;
        RECT 1752.665 2792.570 1753.250 2792.580 ;
        RECT 2415.065 2792.570 2415.395 2792.585 ;
        RECT 2418.030 2792.570 2418.410 2792.580 ;
        RECT 1752.665 2792.270 1753.450 2792.570 ;
        RECT 2415.065 2792.270 2418.410 2792.570 ;
        RECT 1752.665 2792.260 1753.250 2792.270 ;
        RECT 1752.665 2792.255 1752.995 2792.260 ;
        RECT 2415.065 2792.255 2415.395 2792.270 ;
        RECT 2418.030 2792.260 2418.410 2792.270 ;
        RECT 1159.265 2791.900 1159.595 2791.905 ;
        RECT 1193.765 2791.900 1194.095 2791.905 ;
        RECT 1159.265 2791.890 1159.850 2791.900 ;
        RECT 1159.040 2791.590 1159.850 2791.890 ;
        RECT 1159.265 2791.580 1159.850 2791.590 ;
        RECT 1193.510 2791.890 1194.095 2791.900 ;
        RECT 1587.065 2791.900 1587.395 2791.905 ;
        RECT 1587.065 2791.890 1587.650 2791.900 ;
        RECT 1193.510 2791.590 1194.320 2791.890 ;
        RECT 1586.840 2791.590 1587.650 2791.890 ;
        RECT 1193.510 2791.580 1194.095 2791.590 ;
        RECT 1159.265 2791.575 1159.595 2791.580 ;
        RECT 1193.765 2791.575 1194.095 2791.580 ;
        RECT 1587.065 2791.580 1587.650 2791.590 ;
        RECT 1600.865 2791.890 1601.195 2791.905 ;
        RECT 1759.565 2791.900 1759.895 2791.905 ;
        RECT 1602.910 2791.890 1603.290 2791.900 ;
        RECT 1600.865 2791.590 1603.290 2791.890 ;
        RECT 1587.065 2791.575 1587.395 2791.580 ;
        RECT 1600.865 2791.575 1601.195 2791.590 ;
        RECT 1602.910 2791.580 1603.290 2791.590 ;
        RECT 1759.310 2791.890 1759.895 2791.900 ;
        RECT 1773.365 2791.890 1773.695 2791.905 ;
        RECT 1794.065 2791.900 1794.395 2791.905 ;
        RECT 1774.030 2791.890 1774.410 2791.900 ;
        RECT 1794.065 2791.890 1794.650 2791.900 ;
        RECT 1759.310 2791.590 1760.120 2791.890 ;
        RECT 1773.365 2791.590 1774.410 2791.890 ;
        RECT 1793.840 2791.590 1794.650 2791.890 ;
        RECT 1759.310 2791.580 1759.895 2791.590 ;
        RECT 1759.565 2791.575 1759.895 2791.580 ;
        RECT 1773.365 2791.575 1773.695 2791.590 ;
        RECT 1774.030 2791.580 1774.410 2791.590 ;
        RECT 1794.065 2791.580 1794.650 2791.590 ;
        RECT 2387.465 2791.890 2387.795 2791.905 ;
        RECT 2392.270 2791.890 2392.650 2791.900 ;
        RECT 2387.465 2791.590 2392.650 2791.890 ;
        RECT 1794.065 2791.575 1794.395 2791.580 ;
        RECT 2387.465 2791.575 2387.795 2791.590 ;
        RECT 2392.270 2791.580 2392.650 2791.590 ;
        RECT 2428.865 2791.890 2429.195 2791.905 ;
        RECT 2433.670 2791.890 2434.050 2791.900 ;
        RECT 2428.865 2791.590 2434.050 2791.890 ;
        RECT 2428.865 2791.575 2429.195 2791.590 ;
        RECT 2433.670 2791.580 2434.050 2791.590 ;
        RECT 2435.765 2791.890 2436.095 2791.905 ;
        RECT 2439.190 2791.890 2439.570 2791.900 ;
        RECT 2435.765 2791.590 2439.570 2791.890 ;
        RECT 2435.765 2791.575 2436.095 2791.590 ;
        RECT 2439.190 2791.580 2439.570 2791.590 ;
        RECT 410.385 2791.210 410.715 2791.225 ;
        RECT 993.870 2791.210 994.250 2791.220 ;
        RECT 410.385 2790.910 994.250 2791.210 ;
        RECT 410.385 2790.895 410.715 2790.910 ;
        RECT 993.870 2790.900 994.250 2790.910 ;
        RECT 1159.265 2791.210 1159.595 2791.225 ;
        RECT 1164.070 2791.210 1164.450 2791.220 ;
        RECT 1159.265 2790.910 1164.450 2791.210 ;
        RECT 1159.265 2790.895 1159.595 2790.910 ;
        RECT 1164.070 2790.900 1164.450 2790.910 ;
        RECT 1417.070 2791.210 1417.450 2791.220 ;
        RECT 2249.670 2791.210 2250.050 2791.220 ;
        RECT 1417.070 2790.910 2250.050 2791.210 ;
        RECT 1417.070 2790.900 1417.450 2790.910 ;
        RECT 2249.670 2790.900 2250.050 2790.910 ;
        RECT 2307.885 2791.210 2308.215 2791.225 ;
        RECT 2408.165 2791.210 2408.495 2791.225 ;
        RECT 2410.670 2791.210 2411.050 2791.220 ;
        RECT 2307.885 2790.910 2407.330 2791.210 ;
        RECT 2307.885 2790.895 2308.215 2790.910 ;
        RECT 1191.670 2790.530 1192.050 2790.540 ;
        RECT 1193.305 2790.530 1193.635 2790.545 ;
        RECT 1191.670 2790.230 1193.635 2790.530 ;
        RECT 1191.670 2790.220 1192.050 2790.230 ;
        RECT 1193.305 2790.215 1193.635 2790.230 ;
        RECT 1642.265 2790.530 1642.595 2790.545 ;
        RECT 1644.310 2790.530 1644.690 2790.540 ;
        RECT 1642.265 2790.230 1644.690 2790.530 ;
        RECT 1642.265 2790.215 1642.595 2790.230 ;
        RECT 1644.310 2790.220 1644.690 2790.230 ;
        RECT 2380.565 2790.530 2380.895 2790.545 ;
        RECT 2386.750 2790.530 2387.130 2790.540 ;
        RECT 2380.565 2790.230 2387.130 2790.530 ;
        RECT 2380.565 2790.215 2380.895 2790.230 ;
        RECT 2386.750 2790.220 2387.130 2790.230 ;
        RECT 2394.365 2790.530 2394.695 2790.545 ;
        RECT 2398.710 2790.530 2399.090 2790.540 ;
        RECT 2394.365 2790.230 2399.090 2790.530 ;
        RECT 2407.030 2790.530 2407.330 2790.910 ;
        RECT 2408.165 2790.910 2411.050 2791.210 ;
        RECT 2408.165 2790.895 2408.495 2790.910 ;
        RECT 2410.670 2790.900 2411.050 2790.910 ;
        RECT 2445.630 2790.530 2446.010 2790.540 ;
        RECT 2407.030 2790.230 2446.010 2790.530 ;
        RECT 2394.365 2790.215 2394.695 2790.230 ;
        RECT 2398.710 2790.220 2399.090 2790.230 ;
        RECT 2445.630 2790.220 2446.010 2790.230 ;
        RECT 1648.245 2789.860 1648.575 2789.865 ;
        RECT 1647.990 2789.850 1648.575 2789.860 ;
        RECT 1647.790 2789.550 1648.575 2789.850 ;
        RECT 1647.990 2789.540 1648.575 2789.550 ;
        RECT 1648.245 2789.535 1648.575 2789.540 ;
        RECT 2380.565 2789.850 2380.895 2789.865 ;
        RECT 2381.230 2789.850 2381.610 2789.860 ;
        RECT 2380.565 2789.550 2381.610 2789.850 ;
        RECT 2380.565 2789.535 2380.895 2789.550 ;
        RECT 2381.230 2789.540 2381.610 2789.550 ;
        RECT 2235.665 2789.170 2235.995 2789.185 ;
        RECT 2236.790 2789.170 2237.170 2789.180 ;
        RECT 2235.665 2788.870 2237.170 2789.170 ;
        RECT 2235.665 2788.855 2235.995 2788.870 ;
        RECT 2236.790 2788.860 2237.170 2788.870 ;
        RECT 2415.065 2789.170 2415.395 2789.185 ;
        RECT 2417.110 2789.170 2417.490 2789.180 ;
        RECT 2415.065 2788.870 2417.490 2789.170 ;
        RECT 2415.065 2788.855 2415.395 2788.870 ;
        RECT 2417.110 2788.860 2417.490 2788.870 ;
        RECT 1007.465 2788.500 1007.795 2788.505 ;
        RECT 1007.465 2788.490 1008.050 2788.500 ;
        RECT 1007.240 2788.190 1008.050 2788.490 ;
        RECT 1007.465 2788.180 1008.050 2788.190 ;
        RECT 1035.270 2788.490 1035.650 2788.500 ;
        RECT 1038.285 2788.490 1038.615 2788.505 ;
        RECT 1035.270 2788.190 1038.615 2788.490 ;
        RECT 1035.270 2788.180 1035.650 2788.190 ;
        RECT 1007.465 2788.175 1007.795 2788.180 ;
        RECT 1038.285 2788.175 1038.615 2788.190 ;
        RECT 1051.830 2788.490 1052.210 2788.500 ;
        RECT 1055.305 2788.490 1055.635 2788.505 ;
        RECT 1051.830 2788.190 1055.635 2788.490 ;
        RECT 1051.830 2788.180 1052.210 2788.190 ;
        RECT 1055.305 2788.175 1055.635 2788.190 ;
        RECT 1617.885 2788.490 1618.215 2788.505 ;
        RECT 1618.550 2788.490 1618.930 2788.500 ;
        RECT 1617.885 2788.190 1618.930 2788.490 ;
        RECT 1617.885 2788.175 1618.215 2788.190 ;
        RECT 1618.550 2788.180 1618.930 2788.190 ;
        RECT 1624.070 2788.490 1624.450 2788.500 ;
        RECT 1624.785 2788.490 1625.115 2788.505 ;
        RECT 1624.070 2788.190 1625.115 2788.490 ;
        RECT 1624.070 2788.180 1624.450 2788.190 ;
        RECT 1624.785 2788.175 1625.115 2788.190 ;
        RECT 1628.465 2788.490 1628.795 2788.505 ;
        RECT 1631.430 2788.490 1631.810 2788.500 ;
        RECT 1628.465 2788.190 1631.810 2788.490 ;
        RECT 1628.465 2788.175 1628.795 2788.190 ;
        RECT 1631.430 2788.180 1631.810 2788.190 ;
        RECT 1649.625 2788.490 1649.955 2788.505 ;
        RECT 1655.350 2788.490 1655.730 2788.500 ;
        RECT 1649.625 2788.190 1655.730 2788.490 ;
        RECT 1649.625 2788.175 1649.955 2788.190 ;
        RECT 1655.350 2788.180 1655.730 2788.190 ;
        RECT 1683.665 2788.490 1683.995 2788.505 ;
        RECT 1689.390 2788.490 1689.770 2788.500 ;
        RECT 1683.665 2788.190 1689.770 2788.490 ;
        RECT 1683.665 2788.175 1683.995 2788.190 ;
        RECT 1689.390 2788.180 1689.770 2788.190 ;
        RECT 1718.165 2788.490 1718.495 2788.505 ;
        RECT 1724.350 2788.490 1724.730 2788.500 ;
        RECT 1718.165 2788.190 1724.730 2788.490 ;
        RECT 1718.165 2788.175 1718.495 2788.190 ;
        RECT 1724.350 2788.180 1724.730 2788.190 ;
        RECT 1760.485 2788.490 1760.815 2788.505 ;
        RECT 1765.750 2788.490 1766.130 2788.500 ;
        RECT 1760.485 2788.190 1766.130 2788.490 ;
        RECT 1760.485 2788.175 1760.815 2788.190 ;
        RECT 1765.750 2788.180 1766.130 2788.190 ;
        RECT 2421.965 2788.490 2422.295 2788.505 ;
        RECT 2428.150 2788.490 2428.530 2788.500 ;
        RECT 2421.965 2788.190 2428.530 2788.490 ;
        RECT 2421.965 2788.175 2422.295 2788.190 ;
        RECT 2428.150 2788.180 2428.530 2788.190 ;
        RECT 1034.605 2787.820 1034.935 2787.825 ;
        RECT 1034.350 2787.810 1034.935 2787.820 ;
        RECT 1039.870 2787.810 1040.250 2787.820 ;
        RECT 1041.505 2787.810 1041.835 2787.825 ;
        RECT 1034.350 2787.510 1035.160 2787.810 ;
        RECT 1039.870 2787.510 1041.835 2787.810 ;
        RECT 1034.350 2787.500 1034.935 2787.510 ;
        RECT 1039.870 2787.500 1040.250 2787.510 ;
        RECT 1034.605 2787.495 1034.935 2787.500 ;
        RECT 1041.505 2787.495 1041.835 2787.510 ;
        RECT 1046.310 2787.810 1046.690 2787.820 ;
        RECT 1048.405 2787.810 1048.735 2787.825 ;
        RECT 1062.205 2787.820 1062.535 2787.825 ;
        RECT 1046.310 2787.510 1048.735 2787.810 ;
        RECT 1046.310 2787.500 1046.690 2787.510 ;
        RECT 1048.405 2787.495 1048.735 2787.510 ;
        RECT 1061.950 2787.810 1062.535 2787.820 ;
        RECT 1067.470 2787.810 1067.850 2787.820 ;
        RECT 1069.105 2787.810 1069.435 2787.825 ;
        RECT 1061.950 2787.510 1062.760 2787.810 ;
        RECT 1067.470 2787.510 1069.435 2787.810 ;
        RECT 1061.950 2787.500 1062.535 2787.510 ;
        RECT 1067.470 2787.500 1067.850 2787.510 ;
        RECT 1062.205 2787.495 1062.535 2787.500 ;
        RECT 1069.105 2787.495 1069.435 2787.510 ;
        RECT 1073.910 2787.810 1074.290 2787.820 ;
        RECT 1076.005 2787.810 1076.335 2787.825 ;
        RECT 1073.910 2787.510 1076.335 2787.810 ;
        RECT 1073.910 2787.500 1074.290 2787.510 ;
        RECT 1076.005 2787.495 1076.335 2787.510 ;
        RECT 1580.165 2787.810 1580.495 2787.825 ;
        RECT 1580.830 2787.810 1581.210 2787.820 ;
        RECT 1580.165 2787.510 1581.210 2787.810 ;
        RECT 1580.165 2787.495 1580.495 2787.510 ;
        RECT 1580.830 2787.500 1581.210 2787.510 ;
        RECT 1593.965 2787.810 1594.295 2787.825 ;
        RECT 1594.630 2787.810 1595.010 2787.820 ;
        RECT 1593.965 2787.510 1595.010 2787.810 ;
        RECT 1593.965 2787.495 1594.295 2787.510 ;
        RECT 1594.630 2787.500 1595.010 2787.510 ;
        RECT 1601.325 2787.810 1601.655 2787.825 ;
        RECT 1604.750 2787.810 1605.130 2787.820 ;
        RECT 1601.325 2787.510 1605.130 2787.810 ;
        RECT 1601.325 2787.495 1601.655 2787.510 ;
        RECT 1604.750 2787.500 1605.130 2787.510 ;
        RECT 1607.765 2787.810 1608.095 2787.825 ;
        RECT 1613.950 2787.810 1614.330 2787.820 ;
        RECT 1607.765 2787.510 1614.330 2787.810 ;
        RECT 1607.765 2787.495 1608.095 2787.510 ;
        RECT 1613.950 2787.500 1614.330 2787.510 ;
        RECT 1614.665 2787.810 1614.995 2787.825 ;
        RECT 1620.390 2787.810 1620.770 2787.820 ;
        RECT 1614.665 2787.510 1620.770 2787.810 ;
        RECT 1614.665 2787.495 1614.995 2787.510 ;
        RECT 1620.390 2787.500 1620.770 2787.510 ;
        RECT 1621.565 2787.810 1621.895 2787.825 ;
        RECT 1626.830 2787.810 1627.210 2787.820 ;
        RECT 1621.565 2787.510 1627.210 2787.810 ;
        RECT 1621.565 2787.495 1621.895 2787.510 ;
        RECT 1626.830 2787.500 1627.210 2787.510 ;
        RECT 1630.510 2787.810 1630.890 2787.820 ;
        RECT 1631.685 2787.810 1632.015 2787.825 ;
        RECT 1649.165 2787.820 1649.495 2787.825 ;
        RECT 1630.510 2787.510 1632.015 2787.810 ;
        RECT 1630.510 2787.500 1630.890 2787.510 ;
        RECT 1631.685 2787.495 1632.015 2787.510 ;
        RECT 1648.910 2787.810 1649.495 2787.820 ;
        RECT 1656.065 2787.810 1656.395 2787.825 ;
        RECT 1660.870 2787.810 1661.250 2787.820 ;
        RECT 1648.910 2787.510 1649.720 2787.810 ;
        RECT 1656.065 2787.510 1661.250 2787.810 ;
        RECT 1648.910 2787.500 1649.495 2787.510 ;
        RECT 1649.165 2787.495 1649.495 2787.500 ;
        RECT 1656.065 2787.495 1656.395 2787.510 ;
        RECT 1660.870 2787.500 1661.250 2787.510 ;
        RECT 1662.965 2787.810 1663.295 2787.825 ;
        RECT 1666.390 2787.810 1666.770 2787.820 ;
        RECT 1662.965 2787.510 1666.770 2787.810 ;
        RECT 1662.965 2787.495 1663.295 2787.510 ;
        RECT 1666.390 2787.500 1666.770 2787.510 ;
        RECT 1669.865 2787.810 1670.195 2787.825 ;
        RECT 1672.830 2787.810 1673.210 2787.820 ;
        RECT 1669.865 2787.510 1673.210 2787.810 ;
        RECT 1669.865 2787.495 1670.195 2787.510 ;
        RECT 1672.830 2787.500 1673.210 2787.510 ;
        RECT 1676.765 2787.810 1677.095 2787.825 ;
        RECT 1684.125 2787.820 1684.455 2787.825 ;
        RECT 1678.350 2787.810 1678.730 2787.820 ;
        RECT 1676.765 2787.510 1678.730 2787.810 ;
        RECT 1676.765 2787.495 1677.095 2787.510 ;
        RECT 1678.350 2787.500 1678.730 2787.510 ;
        RECT 1683.870 2787.810 1684.455 2787.820 ;
        RECT 1690.565 2787.810 1690.895 2787.825 ;
        RECT 1695.830 2787.810 1696.210 2787.820 ;
        RECT 1683.870 2787.510 1684.680 2787.810 ;
        RECT 1690.565 2787.510 1696.210 2787.810 ;
        RECT 1683.870 2787.500 1684.455 2787.510 ;
        RECT 1684.125 2787.495 1684.455 2787.500 ;
        RECT 1690.565 2787.495 1690.895 2787.510 ;
        RECT 1695.830 2787.500 1696.210 2787.510 ;
        RECT 1697.465 2787.810 1697.795 2787.825 ;
        RECT 1702.270 2787.810 1702.650 2787.820 ;
        RECT 1697.465 2787.510 1702.650 2787.810 ;
        RECT 1697.465 2787.495 1697.795 2787.510 ;
        RECT 1702.270 2787.500 1702.650 2787.510 ;
        RECT 1704.365 2787.810 1704.695 2787.825 ;
        RECT 1708.710 2787.810 1709.090 2787.820 ;
        RECT 1704.365 2787.510 1709.090 2787.810 ;
        RECT 1704.365 2787.495 1704.695 2787.510 ;
        RECT 1708.710 2787.500 1709.090 2787.510 ;
        RECT 1711.265 2787.810 1711.595 2787.825 ;
        RECT 1713.310 2787.810 1713.690 2787.820 ;
        RECT 1711.265 2787.510 1713.690 2787.810 ;
        RECT 1711.265 2787.495 1711.595 2787.510 ;
        RECT 1713.310 2787.500 1713.690 2787.510 ;
        RECT 1718.625 2787.810 1718.955 2787.825 ;
        RECT 1719.750 2787.810 1720.130 2787.820 ;
        RECT 1718.625 2787.510 1720.130 2787.810 ;
        RECT 1718.625 2787.495 1718.955 2787.510 ;
        RECT 1719.750 2787.500 1720.130 2787.510 ;
        RECT 1725.065 2787.810 1725.395 2787.825 ;
        RECT 1730.790 2787.810 1731.170 2787.820 ;
        RECT 1725.065 2787.510 1731.170 2787.810 ;
        RECT 1725.065 2787.495 1725.395 2787.510 ;
        RECT 1730.790 2787.500 1731.170 2787.510 ;
        RECT 1731.965 2787.810 1732.295 2787.825 ;
        RECT 1737.230 2787.810 1737.610 2787.820 ;
        RECT 1731.965 2787.510 1737.610 2787.810 ;
        RECT 1731.965 2787.495 1732.295 2787.510 ;
        RECT 1737.230 2787.500 1737.610 2787.510 ;
        RECT 1738.865 2787.810 1739.195 2787.825 ;
        RECT 1743.670 2787.810 1744.050 2787.820 ;
        RECT 1738.865 2787.510 1744.050 2787.810 ;
        RECT 1738.865 2787.495 1739.195 2787.510 ;
        RECT 1743.670 2787.500 1744.050 2787.510 ;
        RECT 1745.765 2787.810 1746.095 2787.825 ;
        RECT 1748.270 2787.810 1748.650 2787.820 ;
        RECT 1745.765 2787.510 1748.650 2787.810 ;
        RECT 1745.765 2787.495 1746.095 2787.510 ;
        RECT 1748.270 2787.500 1748.650 2787.510 ;
        RECT 1752.665 2787.810 1752.995 2787.825 ;
        RECT 1760.025 2787.820 1760.355 2787.825 ;
        RECT 1754.710 2787.810 1755.090 2787.820 ;
        RECT 1760.025 2787.810 1760.610 2787.820 ;
        RECT 1752.665 2787.510 1755.090 2787.810 ;
        RECT 1759.800 2787.510 1760.610 2787.810 ;
        RECT 1752.665 2787.495 1752.995 2787.510 ;
        RECT 1754.710 2787.500 1755.090 2787.510 ;
        RECT 1760.025 2787.500 1760.610 2787.510 ;
        RECT 1766.465 2787.810 1766.795 2787.825 ;
        RECT 1772.190 2787.810 1772.570 2787.820 ;
        RECT 1766.465 2787.510 1772.570 2787.810 ;
        RECT 1760.025 2787.495 1760.355 2787.500 ;
        RECT 1766.465 2787.495 1766.795 2787.510 ;
        RECT 1772.190 2787.500 1772.570 2787.510 ;
        RECT 1773.825 2787.810 1774.155 2787.825 ;
        RECT 1777.710 2787.810 1778.090 2787.820 ;
        RECT 1773.825 2787.510 1778.090 2787.810 ;
        RECT 1773.825 2787.495 1774.155 2787.510 ;
        RECT 1777.710 2787.500 1778.090 2787.510 ;
        RECT 1780.265 2787.810 1780.595 2787.825 ;
        RECT 1783.230 2787.810 1783.610 2787.820 ;
        RECT 1780.265 2787.510 1783.610 2787.810 ;
        RECT 1780.265 2787.495 1780.595 2787.510 ;
        RECT 1783.230 2787.500 1783.610 2787.510 ;
        RECT 1787.165 2787.810 1787.495 2787.825 ;
        RECT 1789.670 2787.810 1790.050 2787.820 ;
        RECT 1787.165 2787.510 1790.050 2787.810 ;
        RECT 1787.165 2787.495 1787.495 2787.510 ;
        RECT 1789.670 2787.500 1790.050 2787.510 ;
        RECT 1794.525 2787.810 1794.855 2787.825 ;
        RECT 1795.190 2787.810 1795.570 2787.820 ;
        RECT 1794.525 2787.510 1795.570 2787.810 ;
        RECT 1794.525 2787.495 1794.855 2787.510 ;
        RECT 1795.190 2787.500 1795.570 2787.510 ;
        RECT 1828.105 2787.810 1828.435 2787.825 ;
        RECT 1869.505 2787.810 1869.835 2787.825 ;
        RECT 1828.105 2787.510 1869.835 2787.810 ;
        RECT 1828.105 2787.495 1828.435 2787.510 ;
        RECT 1869.505 2787.495 1869.835 2787.510 ;
        RECT 2228.765 2787.810 2229.095 2787.825 ;
        RECT 2231.270 2787.810 2231.650 2787.820 ;
        RECT 2228.765 2787.510 2231.650 2787.810 ;
        RECT 2228.765 2787.495 2229.095 2787.510 ;
        RECT 2231.270 2787.500 2231.650 2787.510 ;
        RECT 305.045 2715.050 305.375 2715.065 ;
        RECT 686.385 2715.050 686.715 2715.065 ;
        RECT 305.045 2714.750 686.715 2715.050 ;
        RECT 305.045 2714.735 305.375 2714.750 ;
        RECT 686.385 2714.735 686.715 2714.750 ;
      LAYER met3 ;
        RECT 305.055 2696.480 1395.530 2697.345 ;
      LAYER met3 ;
        RECT 1395.930 2696.880 1399.930 2697.480 ;
      LAYER met3 ;
        RECT 305.055 2693.120 1395.930 2696.480 ;
        RECT 305.055 2691.720 1395.530 2693.120 ;
      LAYER met3 ;
        RECT 1395.930 2692.120 1399.930 2692.720 ;
      LAYER met3 ;
        RECT 305.055 2687.680 1395.930 2691.720 ;
        RECT 305.055 2686.280 1395.530 2687.680 ;
      LAYER met3 ;
        RECT 1395.930 2686.680 1399.930 2687.280 ;
      LAYER met3 ;
        RECT 305.055 2682.920 1395.930 2686.280 ;
        RECT 305.055 2681.520 1395.530 2682.920 ;
      LAYER met3 ;
        RECT 1395.930 2681.920 1399.930 2682.520 ;
      LAYER met3 ;
        RECT 305.055 2677.480 1395.930 2681.520 ;
        RECT 305.055 2676.080 1395.530 2677.480 ;
      LAYER met3 ;
        RECT 1395.930 2676.480 1399.930 2677.080 ;
      LAYER met3 ;
        RECT 305.055 2672.720 1395.930 2676.080 ;
        RECT 305.055 2671.320 1395.530 2672.720 ;
      LAYER met3 ;
        RECT 1395.930 2671.720 1399.930 2672.320 ;
      LAYER met3 ;
        RECT 305.055 2667.960 1395.930 2671.320 ;
        RECT 305.055 2666.560 1395.530 2667.960 ;
      LAYER met3 ;
        RECT 1395.930 2666.960 1399.930 2667.560 ;
      LAYER met3 ;
        RECT 305.055 2662.520 1395.930 2666.560 ;
        RECT 305.055 2661.120 1395.530 2662.520 ;
      LAYER met3 ;
        RECT 1395.930 2661.520 1399.930 2662.120 ;
      LAYER met3 ;
        RECT 305.055 2657.760 1395.930 2661.120 ;
        RECT 305.055 2656.360 1395.530 2657.760 ;
      LAYER met3 ;
        RECT 1395.930 2656.760 1399.930 2657.360 ;
      LAYER met3 ;
        RECT 305.055 2652.320 1395.930 2656.360 ;
        RECT 305.055 2650.920 1395.530 2652.320 ;
      LAYER met3 ;
        RECT 1395.930 2651.320 1399.930 2651.920 ;
      LAYER met3 ;
        RECT 305.055 2647.560 1395.930 2650.920 ;
        RECT 305.055 2646.160 1395.530 2647.560 ;
      LAYER met3 ;
        RECT 1395.930 2646.560 1399.930 2647.160 ;
      LAYER met3 ;
        RECT 305.055 2642.120 1395.930 2646.160 ;
        RECT 305.055 2640.720 1395.530 2642.120 ;
      LAYER met3 ;
        RECT 1395.930 2641.120 1399.930 2641.720 ;
      LAYER met3 ;
        RECT 305.055 2637.360 1395.930 2640.720 ;
        RECT 305.055 2635.960 1395.530 2637.360 ;
      LAYER met3 ;
        RECT 1395.930 2636.360 1399.930 2636.960 ;
      LAYER met3 ;
        RECT 305.055 2632.600 1395.930 2635.960 ;
        RECT 305.055 2631.200 1395.530 2632.600 ;
      LAYER met3 ;
        RECT 1395.930 2631.600 1399.930 2632.200 ;
      LAYER met3 ;
        RECT 305.055 2627.160 1395.930 2631.200 ;
        RECT 305.055 2625.760 1395.530 2627.160 ;
      LAYER met3 ;
        RECT 1395.930 2626.160 1399.930 2626.760 ;
      LAYER met3 ;
        RECT 305.055 2622.400 1395.930 2625.760 ;
        RECT 305.055 2621.000 1395.530 2622.400 ;
      LAYER met3 ;
        RECT 1395.930 2621.400 1399.930 2622.000 ;
      LAYER met3 ;
        RECT 305.055 2616.960 1395.930 2621.000 ;
        RECT 305.055 2615.560 1395.530 2616.960 ;
      LAYER met3 ;
        RECT 1395.930 2615.960 1399.930 2616.560 ;
      LAYER met3 ;
        RECT 305.055 2612.200 1395.930 2615.560 ;
        RECT 305.055 2610.800 1395.530 2612.200 ;
      LAYER met3 ;
        RECT 1395.930 2611.200 1399.930 2611.800 ;
      LAYER met3 ;
        RECT 305.055 2606.760 1395.930 2610.800 ;
        RECT 305.055 2605.360 1395.530 2606.760 ;
      LAYER met3 ;
        RECT 1395.930 2605.760 1399.930 2606.360 ;
      LAYER met3 ;
        RECT 305.055 2602.000 1395.930 2605.360 ;
        RECT 305.055 2600.600 1395.530 2602.000 ;
      LAYER met3 ;
        RECT 1395.930 2601.000 1399.930 2601.600 ;
      LAYER met3 ;
        RECT 305.055 2597.240 1395.930 2600.600 ;
        RECT 305.055 2595.840 1395.530 2597.240 ;
      LAYER met3 ;
        RECT 1395.930 2596.240 1399.930 2596.840 ;
      LAYER met3 ;
        RECT 305.055 2591.800 1395.930 2595.840 ;
        RECT 305.055 2590.400 1395.530 2591.800 ;
      LAYER met3 ;
        RECT 1395.930 2590.800 1399.930 2591.400 ;
      LAYER met3 ;
        RECT 305.055 2587.040 1395.930 2590.400 ;
        RECT 305.055 2585.640 1395.530 2587.040 ;
      LAYER met3 ;
        RECT 1395.930 2586.040 1399.930 2586.640 ;
      LAYER met3 ;
        RECT 305.055 2581.600 1395.930 2585.640 ;
        RECT 305.055 2580.200 1395.530 2581.600 ;
      LAYER met3 ;
        RECT 1395.930 2580.600 1399.930 2581.200 ;
      LAYER met3 ;
        RECT 305.055 2576.840 1395.930 2580.200 ;
        RECT 305.055 2575.440 1395.530 2576.840 ;
      LAYER met3 ;
        RECT 1395.930 2575.840 1399.930 2576.440 ;
      LAYER met3 ;
        RECT 305.055 2572.080 1395.930 2575.440 ;
        RECT 305.055 2570.680 1395.530 2572.080 ;
      LAYER met3 ;
        RECT 1395.930 2571.080 1399.930 2571.680 ;
      LAYER met3 ;
        RECT 305.055 2566.640 1395.930 2570.680 ;
        RECT 305.055 2565.240 1395.530 2566.640 ;
      LAYER met3 ;
        RECT 1395.930 2565.640 1399.930 2566.240 ;
      LAYER met3 ;
        RECT 305.055 2561.880 1395.930 2565.240 ;
        RECT 305.055 2560.480 1395.530 2561.880 ;
      LAYER met3 ;
        RECT 1395.930 2560.880 1399.930 2561.480 ;
      LAYER met3 ;
        RECT 305.055 2556.440 1395.930 2560.480 ;
        RECT 305.055 2555.040 1395.530 2556.440 ;
      LAYER met3 ;
        RECT 1395.930 2555.440 1399.930 2556.040 ;
      LAYER met3 ;
        RECT 305.055 2551.680 1395.930 2555.040 ;
        RECT 305.055 2550.280 1395.530 2551.680 ;
      LAYER met3 ;
        RECT 1395.930 2550.680 1399.930 2551.280 ;
      LAYER met3 ;
        RECT 305.055 2546.240 1395.930 2550.280 ;
        RECT 305.055 2544.840 1395.530 2546.240 ;
      LAYER met3 ;
        RECT 1395.930 2545.240 1399.930 2545.840 ;
      LAYER met3 ;
        RECT 305.055 2541.480 1395.930 2544.840 ;
        RECT 305.055 2540.080 1395.530 2541.480 ;
      LAYER met3 ;
        RECT 1395.930 2540.480 1399.930 2541.080 ;
      LAYER met3 ;
        RECT 305.055 2536.720 1395.930 2540.080 ;
        RECT 305.055 2535.320 1395.530 2536.720 ;
      LAYER met3 ;
        RECT 1395.930 2535.720 1399.930 2536.320 ;
      LAYER met3 ;
        RECT 305.055 2531.280 1395.930 2535.320 ;
        RECT 305.055 2529.880 1395.530 2531.280 ;
      LAYER met3 ;
        RECT 1395.930 2530.280 1399.930 2530.880 ;
      LAYER met3 ;
        RECT 305.055 2526.520 1395.930 2529.880 ;
        RECT 305.055 2525.120 1395.530 2526.520 ;
      LAYER met3 ;
        RECT 1395.930 2525.520 1399.930 2526.120 ;
      LAYER met3 ;
        RECT 305.055 2521.080 1395.930 2525.120 ;
        RECT 305.055 2519.680 1395.530 2521.080 ;
      LAYER met3 ;
        RECT 1395.930 2520.080 1399.930 2520.680 ;
      LAYER met3 ;
        RECT 305.055 2516.320 1395.930 2519.680 ;
        RECT 305.055 2514.920 1395.530 2516.320 ;
      LAYER met3 ;
        RECT 1395.930 2515.320 1399.930 2515.920 ;
      LAYER met3 ;
        RECT 305.055 2510.880 1395.930 2514.920 ;
        RECT 305.055 2509.480 1395.530 2510.880 ;
      LAYER met3 ;
        RECT 1395.930 2509.880 1399.930 2510.480 ;
      LAYER met3 ;
        RECT 305.055 2506.120 1395.930 2509.480 ;
        RECT 305.055 2504.720 1395.530 2506.120 ;
      LAYER met3 ;
        RECT 1395.930 2505.120 1399.930 2505.720 ;
      LAYER met3 ;
        RECT 305.055 2501.360 1395.930 2504.720 ;
        RECT 305.055 2499.960 1395.530 2501.360 ;
      LAYER met3 ;
        RECT 1395.930 2500.360 1399.930 2500.960 ;
      LAYER met3 ;
        RECT 305.055 2495.920 1395.930 2499.960 ;
        RECT 305.055 2494.520 1395.530 2495.920 ;
      LAYER met3 ;
        RECT 1395.930 2494.920 1399.930 2495.520 ;
      LAYER met3 ;
        RECT 305.055 2491.160 1395.930 2494.520 ;
        RECT 305.055 2489.760 1395.530 2491.160 ;
      LAYER met3 ;
        RECT 1395.930 2490.160 1399.930 2490.760 ;
      LAYER met3 ;
        RECT 305.055 2485.720 1395.930 2489.760 ;
        RECT 305.055 2484.320 1395.530 2485.720 ;
      LAYER met3 ;
        RECT 1395.930 2484.720 1399.930 2485.320 ;
      LAYER met3 ;
        RECT 305.055 2480.960 1395.930 2484.320 ;
        RECT 305.055 2479.560 1395.530 2480.960 ;
      LAYER met3 ;
        RECT 1395.930 2479.960 1399.930 2480.560 ;
      LAYER met3 ;
        RECT 305.055 2476.200 1395.930 2479.560 ;
        RECT 305.055 2474.800 1395.530 2476.200 ;
      LAYER met3 ;
        RECT 1395.930 2475.200 1399.930 2475.800 ;
      LAYER met3 ;
        RECT 305.055 2470.760 1395.930 2474.800 ;
        RECT 305.055 2469.360 1395.530 2470.760 ;
      LAYER met3 ;
        RECT 1395.930 2469.760 1399.930 2470.360 ;
      LAYER met3 ;
        RECT 305.055 2466.000 1395.930 2469.360 ;
        RECT 305.055 2464.600 1395.530 2466.000 ;
      LAYER met3 ;
        RECT 1395.930 2465.000 1399.930 2465.600 ;
      LAYER met3 ;
        RECT 305.055 2460.560 1395.930 2464.600 ;
        RECT 305.055 2459.160 1395.530 2460.560 ;
      LAYER met3 ;
        RECT 1395.930 2459.560 1399.930 2460.160 ;
      LAYER met3 ;
        RECT 305.055 2455.800 1395.930 2459.160 ;
        RECT 305.055 2454.400 1395.530 2455.800 ;
      LAYER met3 ;
        RECT 1395.930 2454.800 1399.930 2455.400 ;
      LAYER met3 ;
        RECT 305.055 2450.360 1395.930 2454.400 ;
        RECT 305.055 2448.960 1395.530 2450.360 ;
      LAYER met3 ;
        RECT 1395.930 2449.360 1399.930 2449.960 ;
      LAYER met3 ;
        RECT 305.055 2445.600 1395.930 2448.960 ;
        RECT 305.055 2444.200 1395.530 2445.600 ;
      LAYER met3 ;
        RECT 1395.930 2444.600 1399.930 2445.200 ;
      LAYER met3 ;
        RECT 305.055 2440.840 1395.930 2444.200 ;
        RECT 305.055 2439.440 1395.530 2440.840 ;
      LAYER met3 ;
        RECT 1395.930 2439.840 1399.930 2440.440 ;
      LAYER met3 ;
        RECT 305.055 2435.400 1395.930 2439.440 ;
        RECT 305.055 2434.000 1395.530 2435.400 ;
      LAYER met3 ;
        RECT 1395.930 2434.400 1399.930 2435.000 ;
      LAYER met3 ;
        RECT 305.055 2430.640 1395.930 2434.000 ;
        RECT 305.055 2429.240 1395.530 2430.640 ;
      LAYER met3 ;
        RECT 1395.930 2429.640 1399.930 2430.240 ;
      LAYER met3 ;
        RECT 305.055 2425.200 1395.930 2429.240 ;
        RECT 305.055 2423.800 1395.530 2425.200 ;
      LAYER met3 ;
        RECT 1395.930 2424.200 1399.930 2424.800 ;
      LAYER met3 ;
        RECT 305.055 2420.440 1395.930 2423.800 ;
        RECT 305.055 2419.040 1395.530 2420.440 ;
      LAYER met3 ;
        RECT 1395.930 2419.440 1399.930 2420.040 ;
      LAYER met3 ;
        RECT 305.055 2415.000 1395.930 2419.040 ;
        RECT 305.055 2413.600 1395.530 2415.000 ;
      LAYER met3 ;
        RECT 1395.930 2414.000 1399.930 2414.600 ;
      LAYER met3 ;
        RECT 305.055 2410.240 1395.930 2413.600 ;
        RECT 305.055 2408.840 1395.530 2410.240 ;
      LAYER met3 ;
        RECT 1395.930 2409.240 1399.930 2409.840 ;
      LAYER met3 ;
        RECT 305.055 2405.480 1395.930 2408.840 ;
        RECT 305.055 2404.080 1395.530 2405.480 ;
      LAYER met3 ;
        RECT 1395.930 2404.480 1399.930 2405.080 ;
      LAYER met3 ;
        RECT 305.055 2400.040 1395.930 2404.080 ;
        RECT 305.055 2398.640 1395.530 2400.040 ;
      LAYER met3 ;
        RECT 1395.930 2399.040 1399.930 2399.640 ;
      LAYER met3 ;
        RECT 305.055 2395.280 1395.930 2398.640 ;
        RECT 305.055 2393.880 1395.530 2395.280 ;
      LAYER met3 ;
        RECT 1395.930 2394.280 1399.930 2394.880 ;
      LAYER met3 ;
        RECT 305.055 2389.840 1395.930 2393.880 ;
        RECT 305.055 2388.440 1395.530 2389.840 ;
      LAYER met3 ;
        RECT 1395.930 2388.840 1399.930 2389.440 ;
      LAYER met3 ;
        RECT 305.055 2385.080 1395.930 2388.440 ;
        RECT 305.055 2383.680 1395.530 2385.080 ;
      LAYER met3 ;
        RECT 1395.930 2384.080 1399.930 2384.680 ;
      LAYER met3 ;
        RECT 305.055 2379.640 1395.930 2383.680 ;
        RECT 305.055 2378.240 1395.530 2379.640 ;
      LAYER met3 ;
        RECT 1395.930 2378.640 1399.930 2379.240 ;
      LAYER met3 ;
        RECT 305.055 2374.880 1395.930 2378.240 ;
        RECT 305.055 2373.480 1395.530 2374.880 ;
      LAYER met3 ;
        RECT 1395.930 2373.880 1399.930 2374.480 ;
      LAYER met3 ;
        RECT 305.055 2370.120 1395.930 2373.480 ;
        RECT 305.055 2368.720 1395.530 2370.120 ;
      LAYER met3 ;
        RECT 1395.930 2369.120 1399.930 2369.720 ;
      LAYER met3 ;
        RECT 305.055 2364.680 1395.930 2368.720 ;
        RECT 305.055 2363.280 1395.530 2364.680 ;
      LAYER met3 ;
        RECT 1395.930 2363.680 1399.930 2364.280 ;
      LAYER met3 ;
        RECT 305.055 2359.920 1395.930 2363.280 ;
        RECT 305.055 2358.520 1395.530 2359.920 ;
      LAYER met3 ;
        RECT 1395.930 2358.920 1399.930 2359.520 ;
      LAYER met3 ;
        RECT 305.055 2354.480 1395.930 2358.520 ;
        RECT 305.055 2353.080 1395.530 2354.480 ;
      LAYER met3 ;
        RECT 1395.930 2353.480 1399.930 2354.080 ;
      LAYER met3 ;
        RECT 305.055 2349.720 1395.930 2353.080 ;
        RECT 305.055 2348.320 1395.530 2349.720 ;
      LAYER met3 ;
        RECT 1395.930 2348.720 1399.930 2349.320 ;
      LAYER met3 ;
        RECT 305.055 2344.960 1395.930 2348.320 ;
        RECT 305.055 2343.560 1395.530 2344.960 ;
      LAYER met3 ;
        RECT 1395.930 2343.960 1399.930 2344.560 ;
      LAYER met3 ;
        RECT 305.055 2339.520 1395.930 2343.560 ;
        RECT 305.055 2338.120 1395.530 2339.520 ;
      LAYER met3 ;
        RECT 1395.930 2338.520 1399.930 2339.120 ;
      LAYER met3 ;
        RECT 305.055 2334.760 1395.930 2338.120 ;
        RECT 305.055 2333.360 1395.530 2334.760 ;
      LAYER met3 ;
        RECT 1395.930 2333.760 1399.930 2334.360 ;
      LAYER met3 ;
        RECT 305.055 2329.320 1395.930 2333.360 ;
        RECT 305.055 2327.920 1395.530 2329.320 ;
      LAYER met3 ;
        RECT 1395.930 2328.320 1399.930 2328.920 ;
      LAYER met3 ;
        RECT 305.055 2324.560 1395.930 2327.920 ;
        RECT 305.055 2323.160 1395.530 2324.560 ;
      LAYER met3 ;
        RECT 1395.930 2323.560 1399.930 2324.160 ;
      LAYER met3 ;
        RECT 305.055 2319.120 1395.930 2323.160 ;
        RECT 305.055 2317.720 1395.530 2319.120 ;
      LAYER met3 ;
        RECT 1395.930 2318.120 1399.930 2318.720 ;
      LAYER met3 ;
        RECT 305.055 2314.360 1395.930 2317.720 ;
        RECT 305.055 2312.960 1395.530 2314.360 ;
      LAYER met3 ;
        RECT 1395.930 2313.360 1399.930 2313.960 ;
      LAYER met3 ;
        RECT 305.055 2309.600 1395.930 2312.960 ;
        RECT 305.055 2308.200 1395.530 2309.600 ;
      LAYER met3 ;
        RECT 1395.930 2308.600 1399.930 2309.200 ;
      LAYER met3 ;
        RECT 305.055 2304.160 1395.930 2308.200 ;
        RECT 305.055 2302.760 1395.530 2304.160 ;
      LAYER met3 ;
        RECT 1395.930 2303.160 1399.930 2303.760 ;
      LAYER met3 ;
        RECT 305.055 2299.400 1395.930 2302.760 ;
        RECT 305.055 2298.000 1395.530 2299.400 ;
      LAYER met3 ;
        RECT 1395.930 2298.400 1399.930 2299.000 ;
      LAYER met3 ;
        RECT 305.055 2293.960 1395.930 2298.000 ;
        RECT 305.055 2292.560 1395.530 2293.960 ;
      LAYER met3 ;
        RECT 1395.930 2292.960 1399.930 2293.560 ;
      LAYER met3 ;
        RECT 305.055 2289.200 1395.930 2292.560 ;
        RECT 305.055 2287.800 1395.530 2289.200 ;
      LAYER met3 ;
        RECT 1395.930 2288.200 1399.930 2288.800 ;
      LAYER met3 ;
        RECT 305.055 2283.760 1395.930 2287.800 ;
        RECT 305.055 2282.360 1395.530 2283.760 ;
      LAYER met3 ;
        RECT 1395.930 2282.760 1399.930 2283.360 ;
      LAYER met3 ;
        RECT 305.055 2279.000 1395.930 2282.360 ;
        RECT 305.055 2277.600 1395.530 2279.000 ;
      LAYER met3 ;
        RECT 1395.930 2278.000 1399.930 2278.600 ;
      LAYER met3 ;
        RECT 305.055 2274.240 1395.930 2277.600 ;
        RECT 305.055 2272.840 1395.530 2274.240 ;
      LAYER met3 ;
        RECT 1395.930 2273.240 1399.930 2273.840 ;
      LAYER met3 ;
        RECT 305.055 2268.800 1395.930 2272.840 ;
        RECT 305.055 2267.400 1395.530 2268.800 ;
      LAYER met3 ;
        RECT 1395.930 2267.800 1399.930 2268.400 ;
      LAYER met3 ;
        RECT 305.055 2264.040 1395.930 2267.400 ;
        RECT 305.055 2262.640 1395.530 2264.040 ;
      LAYER met3 ;
        RECT 1395.930 2263.040 1399.930 2263.640 ;
      LAYER met3 ;
        RECT 305.055 2258.600 1395.930 2262.640 ;
        RECT 305.055 2257.200 1395.530 2258.600 ;
      LAYER met3 ;
        RECT 1395.930 2257.600 1399.930 2258.200 ;
      LAYER met3 ;
        RECT 305.055 2253.840 1395.930 2257.200 ;
        RECT 305.055 2252.440 1395.530 2253.840 ;
      LAYER met3 ;
        RECT 1395.930 2252.840 1399.930 2253.440 ;
      LAYER met3 ;
        RECT 305.055 2249.080 1395.930 2252.440 ;
        RECT 305.055 2247.680 1395.530 2249.080 ;
      LAYER met3 ;
        RECT 1395.930 2248.080 1399.930 2248.680 ;
      LAYER met3 ;
        RECT 305.055 2243.640 1395.930 2247.680 ;
        RECT 305.055 2242.240 1395.530 2243.640 ;
      LAYER met3 ;
        RECT 1395.930 2242.640 1399.930 2243.240 ;
      LAYER met3 ;
        RECT 305.055 2238.880 1395.930 2242.240 ;
        RECT 305.055 2237.480 1395.530 2238.880 ;
      LAYER met3 ;
        RECT 1395.930 2237.880 1399.930 2238.480 ;
      LAYER met3 ;
        RECT 305.055 2233.440 1395.930 2237.480 ;
        RECT 305.055 2232.040 1395.530 2233.440 ;
      LAYER met3 ;
        RECT 1395.930 2232.440 1399.930 2233.040 ;
      LAYER met3 ;
        RECT 305.055 2228.680 1395.930 2232.040 ;
        RECT 305.055 2227.280 1395.530 2228.680 ;
      LAYER met3 ;
        RECT 1395.930 2227.680 1399.930 2228.280 ;
      LAYER met3 ;
        RECT 305.055 2223.240 1395.930 2227.280 ;
        RECT 305.055 2221.840 1395.530 2223.240 ;
      LAYER met3 ;
        RECT 1395.930 2222.240 1399.930 2222.840 ;
      LAYER met3 ;
        RECT 305.055 2218.480 1395.930 2221.840 ;
        RECT 305.055 2217.080 1395.530 2218.480 ;
      LAYER met3 ;
        RECT 1395.930 2217.480 1399.930 2218.080 ;
      LAYER met3 ;
        RECT 305.055 2213.720 1395.930 2217.080 ;
        RECT 305.055 2212.320 1395.530 2213.720 ;
      LAYER met3 ;
        RECT 1395.930 2212.720 1399.930 2213.320 ;
      LAYER met3 ;
        RECT 305.055 2208.280 1395.930 2212.320 ;
        RECT 305.055 2206.880 1395.530 2208.280 ;
      LAYER met3 ;
        RECT 1395.930 2207.280 1399.930 2207.880 ;
      LAYER met3 ;
        RECT 305.055 2203.520 1395.930 2206.880 ;
        RECT 305.055 2202.120 1395.530 2203.520 ;
      LAYER met3 ;
        RECT 1395.930 2202.520 1399.930 2203.120 ;
      LAYER met3 ;
        RECT 305.055 2198.080 1395.930 2202.120 ;
        RECT 305.055 2196.680 1395.530 2198.080 ;
      LAYER met3 ;
        RECT 1395.930 2197.080 1399.930 2197.680 ;
      LAYER met3 ;
        RECT 305.055 2193.320 1395.930 2196.680 ;
        RECT 305.055 2191.920 1395.530 2193.320 ;
      LAYER met3 ;
        RECT 1395.930 2192.320 1399.930 2192.920 ;
      LAYER met3 ;
        RECT 305.055 2187.880 1395.930 2191.920 ;
        RECT 305.055 2186.480 1395.530 2187.880 ;
      LAYER met3 ;
        RECT 1395.930 2186.880 1399.930 2187.480 ;
      LAYER met3 ;
        RECT 305.055 2183.120 1395.930 2186.480 ;
        RECT 305.055 2181.720 1395.530 2183.120 ;
      LAYER met3 ;
        RECT 1395.930 2182.120 1399.930 2182.720 ;
      LAYER met3 ;
        RECT 305.055 2178.360 1395.930 2181.720 ;
        RECT 305.055 2176.960 1395.530 2178.360 ;
      LAYER met3 ;
        RECT 1395.930 2177.360 1399.930 2177.960 ;
      LAYER met3 ;
        RECT 305.055 2172.920 1395.930 2176.960 ;
        RECT 305.055 2171.520 1395.530 2172.920 ;
      LAYER met3 ;
        RECT 1395.930 2171.920 1399.930 2172.520 ;
      LAYER met3 ;
        RECT 305.055 2168.160 1395.930 2171.520 ;
        RECT 305.055 2166.760 1395.530 2168.160 ;
      LAYER met3 ;
        RECT 1395.930 2167.160 1399.930 2167.760 ;
      LAYER met3 ;
        RECT 305.055 2162.720 1395.930 2166.760 ;
        RECT 305.055 2161.320 1395.530 2162.720 ;
      LAYER met3 ;
        RECT 1395.930 2161.720 1399.930 2162.320 ;
      LAYER met3 ;
        RECT 305.055 2157.960 1395.930 2161.320 ;
        RECT 305.055 2156.560 1395.530 2157.960 ;
      LAYER met3 ;
        RECT 1395.930 2156.960 1399.930 2157.560 ;
      LAYER met3 ;
        RECT 305.055 2153.200 1395.930 2156.560 ;
        RECT 305.055 2151.800 1395.530 2153.200 ;
      LAYER met3 ;
        RECT 1395.930 2152.200 1399.930 2152.800 ;
      LAYER met3 ;
        RECT 305.055 2147.760 1395.930 2151.800 ;
        RECT 305.055 2146.360 1395.530 2147.760 ;
      LAYER met3 ;
        RECT 1395.930 2147.250 1399.930 2147.360 ;
        RECT 1410.425 2147.250 1410.755 2147.265 ;
        RECT 1395.930 2146.950 1410.755 2147.250 ;
        RECT 1395.930 2146.760 1399.930 2146.950 ;
        RECT 1410.425 2146.935 1410.755 2146.950 ;
      LAYER met3 ;
        RECT 305.055 2143.000 1395.930 2146.360 ;
        RECT 305.055 2141.600 1395.530 2143.000 ;
      LAYER met3 ;
        RECT 1395.930 2142.490 1399.930 2142.600 ;
        RECT 1414.105 2142.490 1414.435 2142.505 ;
        RECT 1395.930 2142.190 1414.435 2142.490 ;
        RECT 1395.930 2142.000 1399.930 2142.190 ;
        RECT 1414.105 2142.175 1414.435 2142.190 ;
      LAYER met3 ;
        RECT 305.055 2137.560 1395.930 2141.600 ;
        RECT 305.055 2136.160 1395.530 2137.560 ;
      LAYER met3 ;
        RECT 1395.930 2137.050 1399.930 2137.160 ;
        RECT 1414.105 2137.050 1414.435 2137.065 ;
        RECT 1395.930 2136.750 1414.435 2137.050 ;
        RECT 1395.930 2136.560 1399.930 2136.750 ;
        RECT 1414.105 2136.735 1414.435 2136.750 ;
      LAYER met3 ;
        RECT 305.055 2132.800 1395.930 2136.160 ;
        RECT 305.055 2131.400 1395.530 2132.800 ;
      LAYER met3 ;
        RECT 1395.930 2132.290 1399.930 2132.400 ;
        RECT 1413.645 2132.290 1413.975 2132.305 ;
        RECT 1395.930 2131.990 1413.975 2132.290 ;
        RECT 1395.930 2131.800 1399.930 2131.990 ;
        RECT 1413.645 2131.975 1413.975 2131.990 ;
      LAYER met3 ;
        RECT 305.055 2127.360 1395.930 2131.400 ;
        RECT 305.055 2125.960 1395.530 2127.360 ;
      LAYER met3 ;
        RECT 1395.930 2126.850 1399.930 2126.960 ;
        RECT 1410.425 2126.850 1410.755 2126.865 ;
        RECT 1395.930 2126.550 1410.755 2126.850 ;
        RECT 1395.930 2126.360 1399.930 2126.550 ;
        RECT 1410.425 2126.535 1410.755 2126.550 ;
      LAYER met3 ;
        RECT 305.055 2122.600 1395.930 2125.960 ;
        RECT 305.055 2121.200 1395.530 2122.600 ;
      LAYER met3 ;
        RECT 1395.930 2122.090 1399.930 2122.200 ;
        RECT 1414.105 2122.090 1414.435 2122.105 ;
        RECT 1395.930 2121.790 1414.435 2122.090 ;
        RECT 1395.930 2121.600 1399.930 2121.790 ;
        RECT 1414.105 2121.775 1414.435 2121.790 ;
      LAYER met3 ;
        RECT 305.055 2117.840 1395.930 2121.200 ;
        RECT 305.055 2116.440 1395.530 2117.840 ;
      LAYER met3 ;
        RECT 1395.930 2117.330 1399.930 2117.440 ;
        RECT 1414.105 2117.330 1414.435 2117.345 ;
        RECT 1395.930 2117.030 1414.435 2117.330 ;
        RECT 1395.930 2116.840 1399.930 2117.030 ;
        RECT 1414.105 2117.015 1414.435 2117.030 ;
      LAYER met3 ;
        RECT 305.055 2112.400 1395.930 2116.440 ;
        RECT 305.055 2111.000 1395.530 2112.400 ;
      LAYER met3 ;
        RECT 1395.930 2111.890 1399.930 2112.000 ;
        RECT 1410.425 2111.890 1410.755 2111.905 ;
        RECT 1395.930 2111.590 1410.755 2111.890 ;
        RECT 1395.930 2111.400 1399.930 2111.590 ;
        RECT 1410.425 2111.575 1410.755 2111.590 ;
      LAYER met3 ;
        RECT 305.055 2107.640 1395.930 2111.000 ;
        RECT 305.055 2106.240 1395.530 2107.640 ;
      LAYER met3 ;
        RECT 1395.930 2107.130 1399.930 2107.240 ;
        RECT 1414.105 2107.130 1414.435 2107.145 ;
        RECT 1395.930 2106.830 1414.435 2107.130 ;
        RECT 1395.930 2106.640 1399.930 2106.830 ;
        RECT 1414.105 2106.815 1414.435 2106.830 ;
      LAYER met3 ;
        RECT 305.055 2102.200 1395.930 2106.240 ;
        RECT 305.055 2100.800 1395.530 2102.200 ;
      LAYER met3 ;
        RECT 1395.930 2101.690 1399.930 2101.800 ;
        RECT 1414.105 2101.690 1414.435 2101.705 ;
        RECT 1395.930 2101.390 1414.435 2101.690 ;
        RECT 1395.930 2101.200 1399.930 2101.390 ;
        RECT 1414.105 2101.375 1414.435 2101.390 ;
      LAYER met3 ;
        RECT 305.055 2097.440 1395.930 2100.800 ;
        RECT 305.055 2096.040 1395.530 2097.440 ;
      LAYER met3 ;
        RECT 1395.930 2096.930 1399.930 2097.040 ;
        RECT 1414.105 2096.930 1414.435 2096.945 ;
        RECT 1395.930 2096.630 1414.435 2096.930 ;
        RECT 1395.930 2096.440 1399.930 2096.630 ;
        RECT 1414.105 2096.615 1414.435 2096.630 ;
      LAYER met3 ;
        RECT 305.055 2092.000 1395.930 2096.040 ;
        RECT 305.055 2090.600 1395.530 2092.000 ;
      LAYER met3 ;
        RECT 1395.930 2091.490 1399.930 2091.600 ;
        RECT 1410.425 2091.490 1410.755 2091.505 ;
        RECT 1395.930 2091.190 1410.755 2091.490 ;
        RECT 1395.930 2091.000 1399.930 2091.190 ;
        RECT 1410.425 2091.175 1410.755 2091.190 ;
      LAYER met3 ;
        RECT 305.055 2087.240 1395.930 2090.600 ;
      LAYER met3 ;
        RECT 1410.630 2087.410 1411.010 2087.420 ;
        RECT 2193.805 2087.410 2194.135 2087.425 ;
      LAYER met3 ;
        RECT 305.055 2085.840 1395.530 2087.240 ;
      LAYER met3 ;
        RECT 1410.630 2087.110 2194.135 2087.410 ;
        RECT 1410.630 2087.100 1411.010 2087.110 ;
        RECT 2193.805 2087.095 2194.135 2087.110 ;
        RECT 1395.930 2086.730 1399.930 2086.840 ;
        RECT 1409.505 2086.730 1409.835 2086.745 ;
        RECT 1395.930 2086.430 1409.835 2086.730 ;
        RECT 1395.930 2086.240 1399.930 2086.430 ;
        RECT 1409.505 2086.415 1409.835 2086.430 ;
      LAYER met3 ;
        RECT 305.055 2082.480 1395.930 2085.840 ;
        RECT 305.055 2081.080 1395.530 2082.480 ;
      LAYER met3 ;
        RECT 1395.930 2081.970 1399.930 2082.080 ;
        RECT 1414.105 2081.970 1414.435 2081.985 ;
        RECT 1395.930 2081.670 1414.435 2081.970 ;
        RECT 1395.930 2081.480 1399.930 2081.670 ;
        RECT 1414.105 2081.655 1414.435 2081.670 ;
      LAYER met3 ;
        RECT 305.055 2077.040 1395.930 2081.080 ;
        RECT 305.055 2075.640 1395.530 2077.040 ;
      LAYER met3 ;
        RECT 1395.930 2076.530 1399.930 2076.640 ;
        RECT 1414.105 2076.530 1414.435 2076.545 ;
        RECT 1395.930 2076.230 1414.435 2076.530 ;
        RECT 1395.930 2076.040 1399.930 2076.230 ;
        RECT 1414.105 2076.215 1414.435 2076.230 ;
      LAYER met3 ;
        RECT 305.055 2072.280 1395.930 2075.640 ;
        RECT 305.055 2070.880 1395.530 2072.280 ;
      LAYER met3 ;
        RECT 1395.930 2071.770 1399.930 2071.880 ;
        RECT 1413.645 2071.770 1413.975 2071.785 ;
        RECT 1395.930 2071.470 1413.975 2071.770 ;
        RECT 1395.930 2071.280 1399.930 2071.470 ;
        RECT 1413.645 2071.455 1413.975 2071.470 ;
      LAYER met3 ;
        RECT 305.055 2066.840 1395.930 2070.880 ;
        RECT 305.055 2065.440 1395.530 2066.840 ;
      LAYER met3 ;
        RECT 1395.930 2066.330 1399.930 2066.440 ;
        RECT 1414.105 2066.330 1414.435 2066.345 ;
        RECT 1395.930 2066.030 1414.435 2066.330 ;
        RECT 1395.930 2065.840 1399.930 2066.030 ;
        RECT 1414.105 2066.015 1414.435 2066.030 ;
      LAYER met3 ;
        RECT 305.055 2062.080 1395.930 2065.440 ;
        RECT 305.055 2060.680 1395.530 2062.080 ;
      LAYER met3 ;
        RECT 1395.930 2061.570 1399.930 2061.680 ;
        RECT 1414.105 2061.570 1414.435 2061.585 ;
        RECT 1395.930 2061.270 1414.435 2061.570 ;
        RECT 1395.930 2061.080 1399.930 2061.270 ;
        RECT 1414.105 2061.255 1414.435 2061.270 ;
      LAYER met3 ;
        RECT 305.055 2056.640 1395.930 2060.680 ;
        RECT 305.055 2055.240 1395.530 2056.640 ;
      LAYER met3 ;
        RECT 1395.930 2056.130 1399.930 2056.240 ;
        RECT 1409.045 2056.130 1409.375 2056.145 ;
        RECT 1395.930 2055.830 1409.375 2056.130 ;
        RECT 1395.930 2055.640 1399.930 2055.830 ;
        RECT 1409.045 2055.815 1409.375 2055.830 ;
      LAYER met3 ;
        RECT 305.055 2051.880 1395.930 2055.240 ;
        RECT 305.055 2050.480 1395.530 2051.880 ;
      LAYER met3 ;
        RECT 1395.930 2051.370 1399.930 2051.480 ;
        RECT 1408.585 2051.370 1408.915 2051.385 ;
        RECT 1395.930 2051.070 1408.915 2051.370 ;
        RECT 2559.280 2051.235 2561.020 2052.140 ;
        RECT 1395.930 2050.880 1399.930 2051.070 ;
        RECT 1408.585 2051.055 1408.915 2051.070 ;
      LAYER met3 ;
        RECT 305.055 2047.120 1395.930 2050.480 ;
        RECT 305.055 2045.720 1395.530 2047.120 ;
      LAYER met3 ;
        RECT 1395.930 2046.610 1399.930 2046.720 ;
        RECT 1409.045 2046.610 1409.375 2046.625 ;
        RECT 1395.930 2046.310 1409.375 2046.610 ;
        RECT 1395.930 2046.120 1399.930 2046.310 ;
        RECT 1409.045 2046.295 1409.375 2046.310 ;
      LAYER met3 ;
        RECT 305.055 2041.680 1395.930 2045.720 ;
        RECT 305.055 2040.280 1395.530 2041.680 ;
      LAYER met3 ;
        RECT 1395.930 2041.170 1399.930 2041.280 ;
        RECT 1414.565 2041.170 1414.895 2041.185 ;
        RECT 1395.930 2040.870 1414.895 2041.170 ;
        RECT 1395.930 2040.680 1399.930 2040.870 ;
        RECT 1414.565 2040.855 1414.895 2040.870 ;
      LAYER met3 ;
        RECT 305.055 2036.920 1395.930 2040.280 ;
        RECT 305.055 2035.520 1395.530 2036.920 ;
      LAYER met3 ;
        RECT 1395.930 2036.410 1399.930 2036.520 ;
        RECT 1409.505 2036.410 1409.835 2036.425 ;
        RECT 1395.930 2036.110 1409.835 2036.410 ;
        RECT 1395.930 2035.920 1399.930 2036.110 ;
        RECT 1409.505 2036.095 1409.835 2036.110 ;
      LAYER met3 ;
        RECT 305.055 2031.480 1395.930 2035.520 ;
        RECT 305.055 2030.080 1395.530 2031.480 ;
      LAYER met3 ;
        RECT 1395.930 2030.970 1399.930 2031.080 ;
        RECT 1414.105 2030.970 1414.435 2030.985 ;
        RECT 1395.930 2030.670 1414.435 2030.970 ;
        RECT 1395.930 2030.480 1399.930 2030.670 ;
        RECT 1414.105 2030.655 1414.435 2030.670 ;
      LAYER met3 ;
        RECT 305.055 2026.720 1395.930 2030.080 ;
        RECT 305.055 2025.320 1395.530 2026.720 ;
      LAYER met3 ;
        RECT 1395.930 2026.210 1399.930 2026.320 ;
        RECT 1413.185 2026.210 1413.515 2026.225 ;
        RECT 1395.930 2025.910 1413.515 2026.210 ;
        RECT 1395.930 2025.720 1399.930 2025.910 ;
        RECT 1413.185 2025.895 1413.515 2025.910 ;
      LAYER met3 ;
        RECT 305.055 2021.960 1395.930 2025.320 ;
        RECT 305.055 2020.560 1395.530 2021.960 ;
      LAYER met3 ;
        RECT 1395.930 2021.450 1399.930 2021.560 ;
        RECT 1409.045 2021.450 1409.375 2021.465 ;
        RECT 1395.930 2021.150 1409.375 2021.450 ;
        RECT 1395.930 2020.960 1399.930 2021.150 ;
        RECT 1409.045 2021.135 1409.375 2021.150 ;
      LAYER met3 ;
        RECT 305.055 2016.520 1395.930 2020.560 ;
        RECT 305.055 2015.120 1395.530 2016.520 ;
      LAYER met3 ;
        RECT 1395.930 2016.010 1399.930 2016.120 ;
        RECT 1410.425 2016.010 1410.755 2016.025 ;
        RECT 1395.930 2015.710 1410.755 2016.010 ;
        RECT 1395.930 2015.520 1399.930 2015.710 ;
        RECT 1410.425 2015.695 1410.755 2015.710 ;
      LAYER met3 ;
        RECT 305.055 2011.760 1395.930 2015.120 ;
        RECT 305.055 2010.360 1395.530 2011.760 ;
      LAYER met3 ;
        RECT 1395.930 2011.250 1399.930 2011.360 ;
        RECT 1410.425 2011.250 1410.755 2011.265 ;
        RECT 1395.930 2010.950 1410.755 2011.250 ;
        RECT 1395.930 2010.760 1399.930 2010.950 ;
        RECT 1410.425 2010.935 1410.755 2010.950 ;
      LAYER met3 ;
        RECT 305.055 2006.320 1395.930 2010.360 ;
        RECT 305.055 2004.920 1395.530 2006.320 ;
      LAYER met3 ;
        RECT 1395.930 2005.810 1399.930 2005.920 ;
        RECT 1414.105 2005.810 1414.435 2005.825 ;
        RECT 1395.930 2005.510 1414.435 2005.810 ;
        RECT 1395.930 2005.320 1399.930 2005.510 ;
        RECT 1414.105 2005.495 1414.435 2005.510 ;
      LAYER met3 ;
        RECT 305.055 2001.560 1395.930 2004.920 ;
        RECT 305.055 2000.160 1395.530 2001.560 ;
      LAYER met3 ;
        RECT 1395.930 2001.050 1399.930 2001.160 ;
        RECT 1413.645 2001.050 1413.975 2001.065 ;
        RECT 1395.930 2000.750 1413.975 2001.050 ;
        RECT 1395.930 2000.560 1399.930 2000.750 ;
        RECT 1413.645 2000.735 1413.975 2000.750 ;
      LAYER met3 ;
        RECT 305.055 1996.120 1395.930 2000.160 ;
        RECT 305.055 1994.720 1395.530 1996.120 ;
      LAYER met3 ;
        RECT 1395.930 1995.610 1399.930 1995.720 ;
        RECT 1414.105 1995.610 1414.435 1995.625 ;
        RECT 1395.930 1995.310 1414.435 1995.610 ;
        RECT 1395.930 1995.120 1399.930 1995.310 ;
        RECT 1414.105 1995.295 1414.435 1995.310 ;
      LAYER met3 ;
        RECT 305.055 1991.360 1395.930 1994.720 ;
        RECT 305.055 1989.960 1395.530 1991.360 ;
      LAYER met3 ;
        RECT 1395.930 1990.850 1399.930 1990.960 ;
        RECT 1414.105 1990.850 1414.435 1990.865 ;
        RECT 1395.930 1990.550 1414.435 1990.850 ;
        RECT 1395.930 1990.360 1399.930 1990.550 ;
        RECT 1414.105 1990.535 1414.435 1990.550 ;
      LAYER met3 ;
        RECT 305.055 1986.600 1395.930 1989.960 ;
        RECT 305.055 1985.200 1395.530 1986.600 ;
      LAYER met3 ;
        RECT 1395.930 1986.090 1399.930 1986.200 ;
        RECT 1414.105 1986.090 1414.435 1986.105 ;
        RECT 1395.930 1985.790 1414.435 1986.090 ;
        RECT 1395.930 1985.600 1399.930 1985.790 ;
        RECT 1414.105 1985.775 1414.435 1985.790 ;
      LAYER met3 ;
        RECT 305.055 1981.160 1395.930 1985.200 ;
        RECT 305.055 1979.760 1395.530 1981.160 ;
      LAYER met3 ;
        RECT 1395.930 1980.650 1399.930 1980.760 ;
        RECT 1414.105 1980.650 1414.435 1980.665 ;
        RECT 1395.930 1980.350 1414.435 1980.650 ;
        RECT 1395.930 1980.160 1399.930 1980.350 ;
        RECT 1414.105 1980.335 1414.435 1980.350 ;
      LAYER met3 ;
        RECT 305.055 1976.400 1395.930 1979.760 ;
        RECT 305.055 1975.000 1395.530 1976.400 ;
      LAYER met3 ;
        RECT 1395.930 1975.890 1399.930 1976.000 ;
        RECT 1414.105 1975.890 1414.435 1975.905 ;
        RECT 1395.930 1975.590 1414.435 1975.890 ;
        RECT 1395.930 1975.400 1399.930 1975.590 ;
        RECT 1414.105 1975.575 1414.435 1975.590 ;
      LAYER met3 ;
        RECT 305.055 1970.960 1395.930 1975.000 ;
        RECT 305.055 1969.560 1395.530 1970.960 ;
      LAYER met3 ;
        RECT 1395.930 1970.450 1399.930 1970.560 ;
        RECT 1414.105 1970.450 1414.435 1970.465 ;
        RECT 1395.930 1970.150 1414.435 1970.450 ;
        RECT 1395.930 1969.960 1399.930 1970.150 ;
        RECT 1414.105 1970.135 1414.435 1970.150 ;
      LAYER met3 ;
        RECT 305.055 1966.200 1395.930 1969.560 ;
        RECT 305.055 1964.800 1395.530 1966.200 ;
      LAYER met3 ;
        RECT 1395.930 1965.690 1399.930 1965.800 ;
        RECT 1409.505 1965.690 1409.835 1965.705 ;
        RECT 1395.930 1965.390 1409.835 1965.690 ;
        RECT 1395.930 1965.200 1399.930 1965.390 ;
        RECT 1409.505 1965.375 1409.835 1965.390 ;
      LAYER met3 ;
        RECT 305.055 1960.760 1395.930 1964.800 ;
        RECT 305.055 1959.360 1395.530 1960.760 ;
      LAYER met3 ;
        RECT 1395.930 1960.250 1399.930 1960.360 ;
        RECT 1414.105 1960.250 1414.435 1960.265 ;
        RECT 1395.930 1959.950 1414.435 1960.250 ;
        RECT 1395.930 1959.760 1399.930 1959.950 ;
        RECT 1414.105 1959.935 1414.435 1959.950 ;
      LAYER met3 ;
        RECT 305.055 1956.000 1395.930 1959.360 ;
        RECT 305.055 1954.600 1395.530 1956.000 ;
      LAYER met3 ;
        RECT 1395.930 1955.490 1399.930 1955.600 ;
        RECT 1410.425 1955.490 1410.755 1955.505 ;
        RECT 1395.930 1955.190 1410.755 1955.490 ;
        RECT 1395.930 1955.000 1399.930 1955.190 ;
        RECT 1410.425 1955.175 1410.755 1955.190 ;
      LAYER met3 ;
        RECT 305.055 1951.240 1395.930 1954.600 ;
      LAYER met3 ;
        RECT 1550.000 1951.445 1554.600 1951.745 ;
      LAYER met3 ;
        RECT 305.055 1949.840 1395.530 1951.240 ;
      LAYER met3 ;
        RECT 1395.930 1950.730 1399.930 1950.840 ;
        RECT 1413.645 1950.730 1413.975 1950.745 ;
        RECT 1395.930 1950.430 1413.975 1950.730 ;
        RECT 1395.930 1950.240 1399.930 1950.430 ;
        RECT 1413.645 1950.415 1413.975 1950.430 ;
      LAYER met3 ;
        RECT 305.055 1945.800 1395.930 1949.840 ;
      LAYER met3 ;
        RECT 1550.000 1945.805 1554.600 1946.105 ;
      LAYER met3 ;
        RECT 305.055 1944.400 1395.530 1945.800 ;
      LAYER met3 ;
        RECT 1395.930 1945.290 1399.930 1945.400 ;
        RECT 1413.645 1945.290 1413.975 1945.305 ;
        RECT 1395.930 1944.990 1413.975 1945.290 ;
        RECT 1395.930 1944.800 1399.930 1944.990 ;
        RECT 1413.645 1944.975 1413.975 1944.990 ;
      LAYER met3 ;
        RECT 305.055 1941.040 1395.930 1944.400 ;
        RECT 305.055 1939.640 1395.530 1941.040 ;
      LAYER met3 ;
        RECT 1395.930 1940.530 1399.930 1940.640 ;
        RECT 1413.645 1940.530 1413.975 1940.545 ;
        RECT 1395.930 1940.230 1413.975 1940.530 ;
        RECT 1395.930 1940.040 1399.930 1940.230 ;
        RECT 1413.645 1940.215 1413.975 1940.230 ;
      LAYER met3 ;
        RECT 305.055 1935.600 1395.930 1939.640 ;
      LAYER met3 ;
        RECT 1550.000 1937.305 1554.600 1937.605 ;
      LAYER met3 ;
        RECT 305.055 1934.200 1395.530 1935.600 ;
      LAYER met3 ;
        RECT 1395.930 1935.090 1399.930 1935.200 ;
        RECT 1413.645 1935.090 1413.975 1935.105 ;
        RECT 1395.930 1934.790 1413.975 1935.090 ;
        RECT 1395.930 1934.600 1399.930 1934.790 ;
        RECT 1413.645 1934.775 1413.975 1934.790 ;
      LAYER met3 ;
        RECT 305.055 1930.840 1395.930 1934.200 ;
      LAYER met3 ;
        RECT 1550.000 1931.665 1554.600 1931.965 ;
      LAYER met3 ;
        RECT 305.055 1929.440 1395.530 1930.840 ;
      LAYER met3 ;
        RECT 1395.930 1930.330 1399.930 1930.440 ;
        RECT 1413.645 1930.330 1413.975 1930.345 ;
        RECT 1395.930 1930.030 1413.975 1930.330 ;
        RECT 1395.930 1929.840 1399.930 1930.030 ;
        RECT 1413.645 1930.015 1413.975 1930.030 ;
      LAYER met3 ;
        RECT 305.055 1926.080 1395.930 1929.440 ;
        RECT 305.055 1924.680 1395.530 1926.080 ;
      LAYER met3 ;
        RECT 1395.930 1925.570 1399.930 1925.680 ;
        RECT 1413.645 1925.570 1413.975 1925.585 ;
        RECT 1395.930 1925.270 1413.975 1925.570 ;
        RECT 1395.930 1925.080 1399.930 1925.270 ;
        RECT 1413.645 1925.255 1413.975 1925.270 ;
      LAYER met3 ;
        RECT 305.055 1920.640 1395.930 1924.680 ;
      LAYER met3 ;
        RECT 1550.000 1923.165 1554.600 1923.465 ;
        RECT 1414.105 1922.850 1414.435 1922.865 ;
        RECT 1399.630 1922.550 1414.435 1922.850 ;
      LAYER met3 ;
        RECT 305.055 1919.240 1395.530 1920.640 ;
      LAYER met3 ;
        RECT 1399.630 1920.240 1399.930 1922.550 ;
        RECT 1414.105 1922.535 1414.435 1922.550 ;
        RECT 1395.930 1919.640 1399.930 1920.240 ;
      LAYER met3 ;
        RECT 305.055 1915.880 1395.930 1919.240 ;
      LAYER met3 ;
        RECT 1550.000 1917.525 1554.600 1917.825 ;
      LAYER met3 ;
        RECT 305.055 1914.480 1395.530 1915.880 ;
      LAYER met3 ;
        RECT 1395.930 1915.370 1399.930 1915.480 ;
        RECT 1414.105 1915.370 1414.435 1915.385 ;
        RECT 1395.930 1915.070 1414.435 1915.370 ;
        RECT 1395.930 1914.880 1399.930 1915.070 ;
        RECT 1414.105 1915.055 1414.435 1915.070 ;
      LAYER met3 ;
        RECT 305.055 1910.440 1395.930 1914.480 ;
      LAYER met3 ;
        RECT 1414.105 1910.610 1414.435 1910.625 ;
      LAYER met3 ;
        RECT 305.055 1909.040 1395.530 1910.440 ;
      LAYER met3 ;
        RECT 1399.630 1910.310 1414.435 1910.610 ;
        RECT 1399.630 1910.040 1399.930 1910.310 ;
        RECT 1414.105 1910.295 1414.435 1910.310 ;
        RECT 1395.930 1909.440 1399.930 1910.040 ;
      LAYER met3 ;
        RECT 305.055 1905.680 1395.930 1909.040 ;
      LAYER met3 ;
        RECT 1550.000 1909.025 1554.600 1909.325 ;
      LAYER met3 ;
        RECT 305.055 1904.280 1395.530 1905.680 ;
      LAYER met3 ;
        RECT 1395.930 1905.170 1399.930 1905.280 ;
        RECT 1414.105 1905.170 1414.435 1905.185 ;
        RECT 1395.930 1904.870 1414.435 1905.170 ;
        RECT 1395.930 1904.680 1399.930 1904.870 ;
        RECT 1414.105 1904.855 1414.435 1904.870 ;
      LAYER met3 ;
        RECT 305.055 1900.240 1395.930 1904.280 ;
      LAYER met3 ;
        RECT 1414.105 1901.090 1414.435 1901.105 ;
        RECT 1399.630 1900.790 1414.435 1901.090 ;
      LAYER met3 ;
        RECT 305.055 1898.840 1395.530 1900.240 ;
      LAYER met3 ;
        RECT 1399.630 1899.840 1399.930 1900.790 ;
        RECT 1414.105 1900.775 1414.435 1900.790 ;
        RECT 1395.930 1899.240 1399.930 1899.840 ;
      LAYER met3 ;
        RECT 305.055 1895.480 1395.930 1898.840 ;
        RECT 305.055 1894.080 1395.530 1895.480 ;
      LAYER met3 ;
        RECT 1395.930 1894.970 1399.930 1895.080 ;
        RECT 1408.585 1894.970 1408.915 1894.985 ;
        RECT 1395.930 1894.670 1408.915 1894.970 ;
        RECT 1395.930 1894.480 1399.930 1894.670 ;
        RECT 1408.585 1894.655 1408.915 1894.670 ;
      LAYER met3 ;
        RECT 305.055 1890.720 1395.930 1894.080 ;
        RECT 305.055 1889.320 1395.530 1890.720 ;
      LAYER met3 ;
        RECT 1395.930 1890.210 1399.930 1890.320 ;
        RECT 1414.105 1890.210 1414.435 1890.225 ;
        RECT 1395.930 1889.910 1414.435 1890.210 ;
        RECT 1395.930 1889.720 1399.930 1889.910 ;
        RECT 1414.105 1889.895 1414.435 1889.910 ;
      LAYER met3 ;
        RECT 305.055 1885.280 1395.930 1889.320 ;
        RECT 305.055 1883.880 1395.530 1885.280 ;
      LAYER met3 ;
        RECT 1395.930 1884.770 1399.930 1884.880 ;
        RECT 1414.105 1884.770 1414.435 1884.785 ;
        RECT 1395.930 1884.470 1414.435 1884.770 ;
        RECT 1395.930 1884.280 1399.930 1884.470 ;
        RECT 1414.105 1884.455 1414.435 1884.470 ;
      LAYER met3 ;
        RECT 305.055 1880.520 1395.930 1883.880 ;
        RECT 305.055 1879.120 1395.530 1880.520 ;
      LAYER met3 ;
        RECT 1395.930 1880.010 1399.930 1880.120 ;
        RECT 1414.105 1880.010 1414.435 1880.025 ;
        RECT 1395.930 1879.710 1414.435 1880.010 ;
        RECT 1395.930 1879.520 1399.930 1879.710 ;
        RECT 1414.105 1879.695 1414.435 1879.710 ;
      LAYER met3 ;
        RECT 305.055 1875.080 1395.930 1879.120 ;
        RECT 305.055 1873.680 1395.530 1875.080 ;
      LAYER met3 ;
        RECT 1395.930 1874.570 1399.930 1874.680 ;
        RECT 1414.105 1874.570 1414.435 1874.585 ;
        RECT 1395.930 1874.270 1414.435 1874.570 ;
        RECT 1395.930 1874.080 1399.930 1874.270 ;
        RECT 1414.105 1874.255 1414.435 1874.270 ;
      LAYER met3 ;
        RECT 305.055 1870.320 1395.930 1873.680 ;
        RECT 305.055 1868.920 1395.530 1870.320 ;
      LAYER met3 ;
        RECT 1395.930 1869.810 1399.930 1869.920 ;
        RECT 1414.105 1869.810 1414.435 1869.825 ;
        RECT 1395.930 1869.510 1414.435 1869.810 ;
        RECT 1395.930 1869.320 1399.930 1869.510 ;
        RECT 1414.105 1869.495 1414.435 1869.510 ;
      LAYER met3 ;
        RECT 305.055 1864.880 1395.930 1868.920 ;
        RECT 305.055 1863.480 1395.530 1864.880 ;
      LAYER met3 ;
        RECT 1395.930 1864.370 1399.930 1864.480 ;
        RECT 1413.645 1864.370 1413.975 1864.385 ;
        RECT 1395.930 1864.070 1413.975 1864.370 ;
        RECT 1395.930 1863.880 1399.930 1864.070 ;
        RECT 1413.645 1864.055 1413.975 1864.070 ;
      LAYER met3 ;
        RECT 305.055 1860.120 1395.930 1863.480 ;
        RECT 305.055 1858.720 1395.530 1860.120 ;
      LAYER met3 ;
        RECT 1395.930 1859.610 1399.930 1859.720 ;
        RECT 1414.105 1859.610 1414.435 1859.625 ;
        RECT 1395.930 1859.310 1414.435 1859.610 ;
        RECT 1395.930 1859.120 1399.930 1859.310 ;
        RECT 1414.105 1859.295 1414.435 1859.310 ;
      LAYER met3 ;
        RECT 305.055 1855.360 1395.930 1858.720 ;
        RECT 305.055 1853.960 1395.530 1855.360 ;
      LAYER met3 ;
        RECT 1395.930 1854.850 1399.930 1854.960 ;
        RECT 1414.105 1854.850 1414.435 1854.865 ;
        RECT 1395.930 1854.550 1414.435 1854.850 ;
        RECT 1395.930 1854.360 1399.930 1854.550 ;
        RECT 1414.105 1854.535 1414.435 1854.550 ;
      LAYER met3 ;
        RECT 305.055 1849.920 1395.930 1853.960 ;
        RECT 305.055 1848.520 1395.530 1849.920 ;
      LAYER met3 ;
        RECT 1395.930 1849.410 1399.930 1849.520 ;
        RECT 1413.645 1849.410 1413.975 1849.425 ;
        RECT 1395.930 1849.110 1413.975 1849.410 ;
        RECT 1395.930 1848.920 1399.930 1849.110 ;
        RECT 1413.645 1849.095 1413.975 1849.110 ;
      LAYER met3 ;
        RECT 305.055 1845.160 1395.930 1848.520 ;
        RECT 305.055 1843.760 1395.530 1845.160 ;
      LAYER met3 ;
        RECT 1395.930 1844.650 1399.930 1844.760 ;
        RECT 1414.105 1844.650 1414.435 1844.665 ;
        RECT 1395.930 1844.350 1414.435 1844.650 ;
        RECT 1395.930 1844.160 1399.930 1844.350 ;
        RECT 1414.105 1844.335 1414.435 1844.350 ;
      LAYER met3 ;
        RECT 305.055 1839.720 1395.930 1843.760 ;
        RECT 305.055 1838.320 1395.530 1839.720 ;
      LAYER met3 ;
        RECT 1395.930 1839.210 1399.930 1839.320 ;
        RECT 1414.105 1839.210 1414.435 1839.225 ;
        RECT 1395.930 1838.910 1414.435 1839.210 ;
        RECT 1395.930 1838.720 1399.930 1838.910 ;
        RECT 1414.105 1838.895 1414.435 1838.910 ;
      LAYER met3 ;
        RECT 305.055 1834.960 1395.930 1838.320 ;
        RECT 305.055 1833.560 1395.530 1834.960 ;
      LAYER met3 ;
        RECT 1395.930 1834.450 1399.930 1834.560 ;
        RECT 1414.105 1834.450 1414.435 1834.465 ;
        RECT 1395.930 1834.150 1414.435 1834.450 ;
        RECT 1395.930 1833.960 1399.930 1834.150 ;
        RECT 1414.105 1834.135 1414.435 1834.150 ;
      LAYER met3 ;
        RECT 305.055 1829.520 1395.930 1833.560 ;
        RECT 305.055 1828.120 1395.530 1829.520 ;
      LAYER met3 ;
        RECT 1395.930 1829.010 1399.930 1829.120 ;
        RECT 1414.105 1829.010 1414.435 1829.025 ;
        RECT 1395.930 1828.710 1414.435 1829.010 ;
        RECT 1395.930 1828.520 1399.930 1828.710 ;
        RECT 1414.105 1828.695 1414.435 1828.710 ;
      LAYER met3 ;
        RECT 305.055 1824.760 1395.930 1828.120 ;
        RECT 305.055 1823.360 1395.530 1824.760 ;
      LAYER met3 ;
        RECT 1395.930 1824.250 1399.930 1824.360 ;
        RECT 1408.585 1824.250 1408.915 1824.265 ;
        RECT 1395.930 1823.950 1408.915 1824.250 ;
        RECT 1395.930 1823.760 1399.930 1823.950 ;
        RECT 1408.585 1823.935 1408.915 1823.950 ;
      LAYER met3 ;
        RECT 305.055 1820.000 1395.930 1823.360 ;
        RECT 305.055 1818.600 1395.530 1820.000 ;
      LAYER met3 ;
        RECT 1395.930 1819.490 1399.930 1819.600 ;
        RECT 1408.585 1819.490 1408.915 1819.505 ;
        RECT 1395.930 1819.190 1408.915 1819.490 ;
        RECT 1395.930 1819.000 1399.930 1819.190 ;
        RECT 1408.585 1819.175 1408.915 1819.190 ;
      LAYER met3 ;
        RECT 305.055 1814.560 1395.930 1818.600 ;
        RECT 305.055 1813.160 1395.530 1814.560 ;
      LAYER met3 ;
        RECT 1395.930 1814.050 1399.930 1814.160 ;
        RECT 1408.585 1814.050 1408.915 1814.065 ;
        RECT 1395.930 1813.750 1408.915 1814.050 ;
        RECT 1395.930 1813.560 1399.930 1813.750 ;
        RECT 1408.585 1813.735 1408.915 1813.750 ;
      LAYER met3 ;
        RECT 305.055 1809.800 1395.930 1813.160 ;
        RECT 305.055 1808.400 1395.530 1809.800 ;
      LAYER met3 ;
        RECT 1395.930 1809.290 1399.930 1809.400 ;
        RECT 1408.585 1809.290 1408.915 1809.305 ;
        RECT 1395.930 1808.990 1408.915 1809.290 ;
        RECT 1395.930 1808.800 1399.930 1808.990 ;
        RECT 1408.585 1808.975 1408.915 1808.990 ;
      LAYER met3 ;
        RECT 305.055 1804.360 1395.930 1808.400 ;
        RECT 305.055 1802.960 1395.530 1804.360 ;
      LAYER met3 ;
        RECT 1395.930 1803.850 1399.930 1803.960 ;
        RECT 1414.105 1803.850 1414.435 1803.865 ;
        RECT 1395.930 1803.550 1414.435 1803.850 ;
        RECT 1395.930 1803.360 1399.930 1803.550 ;
        RECT 1414.105 1803.535 1414.435 1803.550 ;
      LAYER met3 ;
        RECT 305.055 1799.600 1395.930 1802.960 ;
        RECT 305.055 1798.200 1395.530 1799.600 ;
      LAYER met3 ;
        RECT 1395.930 1799.090 1399.930 1799.200 ;
        RECT 1408.585 1799.090 1408.915 1799.105 ;
        RECT 1395.930 1798.790 1408.915 1799.090 ;
        RECT 1395.930 1798.600 1399.930 1798.790 ;
        RECT 1408.585 1798.775 1408.915 1798.790 ;
      LAYER met3 ;
        RECT 305.055 1794.840 1395.930 1798.200 ;
        RECT 305.055 1793.440 1395.530 1794.840 ;
      LAYER met3 ;
        RECT 1395.930 1794.330 1399.930 1794.440 ;
        RECT 1409.045 1794.330 1409.375 1794.345 ;
        RECT 1395.930 1794.030 1409.375 1794.330 ;
        RECT 1395.930 1793.840 1399.930 1794.030 ;
        RECT 1409.045 1794.015 1409.375 1794.030 ;
      LAYER met3 ;
        RECT 305.055 1789.400 1395.930 1793.440 ;
        RECT 305.055 1788.000 1395.530 1789.400 ;
      LAYER met3 ;
        RECT 1395.930 1788.890 1399.930 1789.000 ;
        RECT 1411.805 1788.890 1412.135 1788.905 ;
        RECT 1395.930 1788.590 1412.135 1788.890 ;
        RECT 1395.930 1788.400 1399.930 1788.590 ;
        RECT 1411.805 1788.575 1412.135 1788.590 ;
      LAYER met3 ;
        RECT 305.055 1784.640 1395.930 1788.000 ;
        RECT 305.055 1783.240 1395.530 1784.640 ;
      LAYER met3 ;
        RECT 1395.930 1784.130 1399.930 1784.240 ;
        RECT 1414.105 1784.130 1414.435 1784.145 ;
        RECT 1395.930 1783.830 1414.435 1784.130 ;
        RECT 1395.930 1783.640 1399.930 1783.830 ;
        RECT 1414.105 1783.815 1414.435 1783.830 ;
      LAYER met3 ;
        RECT 305.055 1779.200 1395.930 1783.240 ;
        RECT 305.055 1777.800 1395.530 1779.200 ;
      LAYER met3 ;
        RECT 1395.930 1778.690 1399.930 1778.800 ;
        RECT 1408.585 1778.690 1408.915 1778.705 ;
        RECT 1395.930 1778.390 1408.915 1778.690 ;
        RECT 1395.930 1778.200 1399.930 1778.390 ;
        RECT 1408.585 1778.375 1408.915 1778.390 ;
      LAYER met3 ;
        RECT 305.055 1774.440 1395.930 1777.800 ;
        RECT 305.055 1773.040 1395.530 1774.440 ;
      LAYER met3 ;
        RECT 1395.930 1773.930 1399.930 1774.040 ;
        RECT 1408.585 1773.930 1408.915 1773.945 ;
        RECT 1395.930 1773.630 1408.915 1773.930 ;
        RECT 1395.930 1773.440 1399.930 1773.630 ;
        RECT 1408.585 1773.615 1408.915 1773.630 ;
      LAYER met3 ;
        RECT 305.055 1769.000 1395.930 1773.040 ;
        RECT 305.055 1767.600 1395.530 1769.000 ;
      LAYER met3 ;
        RECT 1395.930 1768.490 1399.930 1768.600 ;
        RECT 1408.585 1768.490 1408.915 1768.505 ;
        RECT 1395.930 1768.190 1408.915 1768.490 ;
        RECT 1395.930 1768.000 1399.930 1768.190 ;
        RECT 1408.585 1768.175 1408.915 1768.190 ;
      LAYER met3 ;
        RECT 305.055 1764.240 1395.930 1767.600 ;
        RECT 305.055 1762.840 1395.530 1764.240 ;
      LAYER met3 ;
        RECT 1395.930 1763.730 1399.930 1763.840 ;
        RECT 1408.585 1763.730 1408.915 1763.745 ;
        RECT 1395.930 1763.430 1408.915 1763.730 ;
        RECT 1395.930 1763.240 1399.930 1763.430 ;
        RECT 1408.585 1763.415 1408.915 1763.430 ;
      LAYER met3 ;
        RECT 305.055 1759.480 1395.930 1762.840 ;
        RECT 305.055 1758.080 1395.530 1759.480 ;
      LAYER met3 ;
        RECT 1395.930 1758.970 1399.930 1759.080 ;
        RECT 1413.185 1758.970 1413.515 1758.985 ;
        RECT 1395.930 1758.670 1413.515 1758.970 ;
        RECT 1395.930 1758.480 1399.930 1758.670 ;
        RECT 1413.185 1758.655 1413.515 1758.670 ;
      LAYER met3 ;
        RECT 305.055 1754.040 1395.930 1758.080 ;
        RECT 305.055 1752.640 1395.530 1754.040 ;
      LAYER met3 ;
        RECT 1395.930 1753.530 1399.930 1753.640 ;
        RECT 1408.585 1753.530 1408.915 1753.545 ;
        RECT 1395.930 1753.230 1408.915 1753.530 ;
        RECT 1395.930 1753.040 1399.930 1753.230 ;
        RECT 1408.585 1753.215 1408.915 1753.230 ;
      LAYER met3 ;
        RECT 305.055 1749.280 1395.930 1752.640 ;
        RECT 305.055 1747.880 1395.530 1749.280 ;
      LAYER met3 ;
        RECT 1395.930 1748.770 1399.930 1748.880 ;
        RECT 1412.725 1748.770 1413.055 1748.785 ;
        RECT 1395.930 1748.470 1413.055 1748.770 ;
        RECT 1395.930 1748.280 1399.930 1748.470 ;
        RECT 1412.725 1748.455 1413.055 1748.470 ;
      LAYER met3 ;
        RECT 305.055 1743.840 1395.930 1747.880 ;
        RECT 305.055 1742.440 1395.530 1743.840 ;
      LAYER met3 ;
        RECT 1395.930 1743.330 1399.930 1743.440 ;
        RECT 1414.105 1743.330 1414.435 1743.345 ;
        RECT 1395.930 1743.030 1414.435 1743.330 ;
        RECT 1395.930 1742.840 1399.930 1743.030 ;
        RECT 1414.105 1743.015 1414.435 1743.030 ;
      LAYER met3 ;
        RECT 305.055 1739.080 1395.930 1742.440 ;
        RECT 305.055 1737.680 1395.530 1739.080 ;
      LAYER met3 ;
        RECT 1395.930 1738.570 1399.930 1738.680 ;
        RECT 1414.105 1738.570 1414.435 1738.585 ;
        RECT 1395.930 1738.270 1414.435 1738.570 ;
        RECT 1395.930 1738.080 1399.930 1738.270 ;
        RECT 1414.105 1738.255 1414.435 1738.270 ;
      LAYER met3 ;
        RECT 305.055 1733.640 1395.930 1737.680 ;
        RECT 305.055 1732.240 1395.530 1733.640 ;
      LAYER met3 ;
        RECT 1395.930 1733.130 1399.930 1733.240 ;
        RECT 1409.965 1733.130 1410.295 1733.145 ;
        RECT 1395.930 1732.830 1410.295 1733.130 ;
        RECT 1395.930 1732.640 1399.930 1732.830 ;
        RECT 1409.965 1732.815 1410.295 1732.830 ;
      LAYER met3 ;
        RECT 305.055 1728.880 1395.930 1732.240 ;
        RECT 305.055 1727.480 1395.530 1728.880 ;
      LAYER met3 ;
        RECT 1395.930 1728.370 1399.930 1728.480 ;
        RECT 1414.105 1728.370 1414.435 1728.385 ;
        RECT 1395.930 1728.070 1414.435 1728.370 ;
        RECT 1395.930 1727.880 1399.930 1728.070 ;
        RECT 1414.105 1728.055 1414.435 1728.070 ;
      LAYER met3 ;
        RECT 305.055 1724.120 1395.930 1727.480 ;
        RECT 305.055 1722.720 1395.530 1724.120 ;
      LAYER met3 ;
        RECT 1395.930 1723.610 1399.930 1723.720 ;
        RECT 1413.645 1723.610 1413.975 1723.625 ;
        RECT 1395.930 1723.310 1413.975 1723.610 ;
        RECT 1395.930 1723.120 1399.930 1723.310 ;
        RECT 1413.645 1723.295 1413.975 1723.310 ;
      LAYER met3 ;
        RECT 305.055 1718.680 1395.930 1722.720 ;
        RECT 305.055 1717.280 1395.530 1718.680 ;
      LAYER met3 ;
        RECT 1395.930 1718.170 1399.930 1718.280 ;
        RECT 1410.425 1718.170 1410.755 1718.185 ;
        RECT 1395.930 1717.870 1410.755 1718.170 ;
        RECT 1395.930 1717.680 1399.930 1717.870 ;
        RECT 1410.425 1717.855 1410.755 1717.870 ;
      LAYER met3 ;
        RECT 305.055 1713.920 1395.930 1717.280 ;
        RECT 305.055 1712.520 1395.530 1713.920 ;
      LAYER met3 ;
        RECT 1395.930 1713.410 1399.930 1713.520 ;
        RECT 1409.965 1713.410 1410.295 1713.425 ;
        RECT 1395.930 1713.110 1410.295 1713.410 ;
        RECT 1395.930 1712.920 1399.930 1713.110 ;
        RECT 1409.965 1713.095 1410.295 1713.110 ;
      LAYER met3 ;
        RECT 305.055 1708.480 1395.930 1712.520 ;
        RECT 305.055 1707.080 1395.530 1708.480 ;
      LAYER met3 ;
        RECT 1395.930 1707.970 1399.930 1708.080 ;
        RECT 1414.105 1707.970 1414.435 1707.985 ;
        RECT 1395.930 1707.670 1414.435 1707.970 ;
        RECT 1395.930 1707.480 1399.930 1707.670 ;
        RECT 1414.105 1707.655 1414.435 1707.670 ;
      LAYER met3 ;
        RECT 305.055 1703.720 1395.930 1707.080 ;
        RECT 305.055 1702.320 1395.530 1703.720 ;
      LAYER met3 ;
        RECT 1395.930 1703.210 1399.930 1703.320 ;
        RECT 1409.505 1703.210 1409.835 1703.225 ;
        RECT 1395.930 1702.910 1409.835 1703.210 ;
        RECT 1395.930 1702.720 1399.930 1702.910 ;
        RECT 1409.505 1702.895 1409.835 1702.910 ;
      LAYER met3 ;
        RECT 305.055 1698.960 1395.930 1702.320 ;
        RECT 305.055 1697.560 1395.530 1698.960 ;
      LAYER met3 ;
        RECT 1395.930 1698.450 1399.930 1698.560 ;
        RECT 1409.045 1698.450 1409.375 1698.465 ;
        RECT 1395.930 1698.150 1409.375 1698.450 ;
        RECT 1395.930 1697.960 1399.930 1698.150 ;
        RECT 1409.045 1698.135 1409.375 1698.150 ;
      LAYER met3 ;
        RECT 305.055 1693.520 1395.930 1697.560 ;
        RECT 305.055 1692.120 1395.530 1693.520 ;
      LAYER met3 ;
        RECT 1395.930 1693.010 1399.930 1693.120 ;
        RECT 1409.505 1693.010 1409.835 1693.025 ;
        RECT 1395.930 1692.710 1409.835 1693.010 ;
        RECT 1395.930 1692.520 1399.930 1692.710 ;
        RECT 1409.505 1692.695 1409.835 1692.710 ;
      LAYER met3 ;
        RECT 305.055 1688.760 1395.930 1692.120 ;
        RECT 305.055 1687.360 1395.530 1688.760 ;
      LAYER met3 ;
        RECT 1395.930 1688.250 1399.930 1688.360 ;
        RECT 1409.505 1688.250 1409.835 1688.265 ;
        RECT 1395.930 1687.950 1409.835 1688.250 ;
        RECT 1395.930 1687.760 1399.930 1687.950 ;
        RECT 1409.505 1687.935 1409.835 1687.950 ;
      LAYER met3 ;
        RECT 305.055 1683.320 1395.930 1687.360 ;
        RECT 305.055 1681.920 1395.530 1683.320 ;
      LAYER met3 ;
        RECT 1395.930 1682.810 1399.930 1682.920 ;
        RECT 1411.805 1682.810 1412.135 1682.825 ;
        RECT 1395.930 1682.510 1412.135 1682.810 ;
        RECT 1395.930 1682.320 1399.930 1682.510 ;
        RECT 1411.805 1682.495 1412.135 1682.510 ;
      LAYER met3 ;
        RECT 305.055 1678.560 1395.930 1681.920 ;
        RECT 305.055 1677.160 1395.530 1678.560 ;
      LAYER met3 ;
        RECT 1395.930 1678.050 1399.930 1678.160 ;
        RECT 1411.805 1678.050 1412.135 1678.065 ;
        RECT 1395.930 1677.750 1412.135 1678.050 ;
        RECT 1395.930 1677.560 1399.930 1677.750 ;
        RECT 1411.805 1677.735 1412.135 1677.750 ;
      LAYER met3 ;
        RECT 305.055 1673.120 1395.930 1677.160 ;
        RECT 305.055 1671.720 1395.530 1673.120 ;
      LAYER met3 ;
        RECT 1395.930 1672.610 1399.930 1672.720 ;
        RECT 1410.425 1672.610 1410.755 1672.625 ;
        RECT 1395.930 1672.310 1410.755 1672.610 ;
        RECT 1395.930 1672.120 1399.930 1672.310 ;
        RECT 1410.425 1672.295 1410.755 1672.310 ;
      LAYER met3 ;
        RECT 305.055 1668.360 1395.930 1671.720 ;
        RECT 305.055 1666.960 1395.530 1668.360 ;
      LAYER met3 ;
        RECT 1395.930 1667.850 1399.930 1667.960 ;
        RECT 1409.505 1667.850 1409.835 1667.865 ;
        RECT 1395.930 1667.550 1409.835 1667.850 ;
        RECT 1395.930 1667.360 1399.930 1667.550 ;
        RECT 1409.505 1667.535 1409.835 1667.550 ;
      LAYER met3 ;
        RECT 305.055 1663.600 1395.930 1666.960 ;
        RECT 305.055 1662.200 1395.530 1663.600 ;
      LAYER met3 ;
        RECT 1395.930 1663.090 1399.930 1663.200 ;
        RECT 1411.805 1663.090 1412.135 1663.105 ;
        RECT 1395.930 1662.790 1412.135 1663.090 ;
        RECT 1395.930 1662.600 1399.930 1662.790 ;
        RECT 1411.805 1662.775 1412.135 1662.790 ;
      LAYER met3 ;
        RECT 305.055 1658.160 1395.930 1662.200 ;
        RECT 305.055 1656.760 1395.530 1658.160 ;
      LAYER met3 ;
        RECT 1395.930 1657.650 1399.930 1657.760 ;
        RECT 1410.630 1657.650 1411.010 1657.660 ;
        RECT 1395.930 1657.350 1411.010 1657.650 ;
        RECT 1395.930 1657.160 1399.930 1657.350 ;
        RECT 1410.630 1657.340 1411.010 1657.350 ;
      LAYER met3 ;
        RECT 305.055 1653.400 1395.930 1656.760 ;
        RECT 305.055 1652.000 1395.530 1653.400 ;
      LAYER met3 ;
        RECT 1395.930 1652.890 1399.930 1653.000 ;
        RECT 1414.105 1652.890 1414.435 1652.905 ;
        RECT 1395.930 1652.590 1414.435 1652.890 ;
        RECT 1395.930 1652.400 1399.930 1652.590 ;
        RECT 1414.105 1652.575 1414.435 1652.590 ;
      LAYER met3 ;
        RECT 305.055 1647.960 1395.930 1652.000 ;
        RECT 305.055 1646.560 1395.530 1647.960 ;
      LAYER met3 ;
        RECT 1395.930 1647.450 1399.930 1647.560 ;
        RECT 1409.505 1647.450 1409.835 1647.465 ;
        RECT 1395.930 1647.150 1409.835 1647.450 ;
        RECT 1395.930 1646.960 1399.930 1647.150 ;
        RECT 1409.505 1647.135 1409.835 1647.150 ;
      LAYER met3 ;
        RECT 305.055 1643.200 1395.930 1646.560 ;
        RECT 305.055 1641.800 1395.530 1643.200 ;
      LAYER met3 ;
        RECT 1395.930 1642.690 1399.930 1642.800 ;
        RECT 1410.425 1642.690 1410.755 1642.705 ;
        RECT 1395.930 1642.390 1410.755 1642.690 ;
        RECT 1395.930 1642.200 1399.930 1642.390 ;
        RECT 1410.425 1642.375 1410.755 1642.390 ;
      LAYER met3 ;
        RECT 305.055 1637.760 1395.930 1641.800 ;
        RECT 305.055 1636.360 1395.530 1637.760 ;
      LAYER met3 ;
        RECT 1395.930 1637.250 1399.930 1637.360 ;
        RECT 1411.345 1637.250 1411.675 1637.265 ;
        RECT 1395.930 1636.950 1411.675 1637.250 ;
        RECT 1395.930 1636.760 1399.930 1636.950 ;
        RECT 1411.345 1636.935 1411.675 1636.950 ;
      LAYER met3 ;
        RECT 305.055 1633.000 1395.930 1636.360 ;
        RECT 305.055 1631.600 1395.530 1633.000 ;
      LAYER met3 ;
        RECT 1395.930 1632.490 1399.930 1632.600 ;
        RECT 1410.425 1632.490 1410.755 1632.505 ;
        RECT 1395.930 1632.190 1410.755 1632.490 ;
        RECT 1395.930 1632.000 1399.930 1632.190 ;
        RECT 1410.425 1632.175 1410.755 1632.190 ;
      LAYER met3 ;
        RECT 305.055 1628.240 1395.930 1631.600 ;
        RECT 305.055 1626.840 1395.530 1628.240 ;
      LAYER met3 ;
        RECT 1395.930 1627.730 1399.930 1627.840 ;
        RECT 1417.070 1627.730 1417.450 1627.740 ;
        RECT 1395.930 1627.430 1417.450 1627.730 ;
        RECT 1395.930 1627.240 1399.930 1627.430 ;
        RECT 1417.070 1627.420 1417.450 1627.430 ;
      LAYER met3 ;
        RECT 305.055 1622.800 1395.930 1626.840 ;
        RECT 305.055 1621.400 1395.530 1622.800 ;
      LAYER met3 ;
        RECT 1395.930 1622.290 1399.930 1622.400 ;
        RECT 1412.265 1622.290 1412.595 1622.305 ;
        RECT 1395.930 1621.990 1412.595 1622.290 ;
        RECT 1395.930 1621.800 1399.930 1621.990 ;
        RECT 1412.265 1621.975 1412.595 1621.990 ;
      LAYER met3 ;
        RECT 305.055 1618.040 1395.930 1621.400 ;
        RECT 305.055 1616.640 1395.530 1618.040 ;
      LAYER met3 ;
        RECT 1395.930 1617.530 1399.930 1617.640 ;
        RECT 1410.885 1617.530 1411.215 1617.545 ;
        RECT 1395.930 1617.230 1411.215 1617.530 ;
        RECT 1395.930 1617.040 1399.930 1617.230 ;
        RECT 1410.885 1617.215 1411.215 1617.230 ;
      LAYER met3 ;
        RECT 305.055 1612.600 1395.930 1616.640 ;
        RECT 305.055 1611.200 1395.530 1612.600 ;
      LAYER met3 ;
        RECT 1395.930 1612.090 1399.930 1612.200 ;
        RECT 1408.125 1612.090 1408.455 1612.105 ;
        RECT 1395.930 1611.790 1408.455 1612.090 ;
        RECT 1395.930 1611.600 1399.930 1611.790 ;
        RECT 1408.125 1611.775 1408.455 1611.790 ;
      LAYER met3 ;
        RECT 305.055 1607.840 1395.930 1611.200 ;
        RECT 305.055 1606.440 1395.530 1607.840 ;
      LAYER met3 ;
        RECT 1550.000 1607.670 1554.600 1607.970 ;
        RECT 1395.930 1607.330 1399.930 1607.440 ;
        RECT 1407.665 1607.330 1407.995 1607.345 ;
        RECT 1395.930 1607.030 1407.995 1607.330 ;
        RECT 1395.930 1606.840 1399.930 1607.030 ;
        RECT 1407.665 1607.015 1407.995 1607.030 ;
      LAYER met3 ;
        RECT 305.055 1603.080 1395.930 1606.440 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
      LAYER met3 ;
        RECT 2200.000 2032.785 2204.600 2033.085 ;
        RECT 2200.000 2027.145 2204.600 2027.445 ;
        RECT 2200.000 2018.645 2204.600 2018.945 ;
        RECT 2200.000 2013.005 2204.600 2013.305 ;
        RECT 2200.000 2004.505 2204.600 2004.805 ;
        RECT 2200.000 1998.865 2204.600 1999.165 ;
        RECT 2200.000 1990.365 2204.600 1990.665 ;
        RECT 1931.880 1963.310 1936.480 1963.610 ;
        RECT 1931.880 1954.810 1936.480 1955.110 ;
        RECT 2200.000 1701.125 2204.600 1701.425 ;
        RECT 2200.000 1692.625 2204.600 1692.925 ;
        RECT 1931.880 1665.570 1936.480 1665.870 ;
        RECT 1931.880 1657.070 1936.480 1657.370 ;
        RECT 1931.880 1651.430 1936.480 1651.730 ;
        RECT 1931.880 1642.930 1936.480 1643.230 ;
        RECT 1931.880 1637.290 1936.480 1637.590 ;
        RECT 1931.880 1628.790 1936.480 1629.090 ;
        RECT 1931.880 1623.150 1936.480 1623.450 ;
      LAYER met3 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
      LAYER met3 ;
        RECT 2581.880 2048.265 2586.480 2048.565 ;
        RECT 2581.880 1746.910 2586.480 1747.210 ;
        RECT 2581.880 1738.410 2586.480 1738.710 ;
        RECT 2581.880 1732.770 2586.480 1733.070 ;
        RECT 2581.880 1724.270 2586.480 1724.570 ;
        RECT 2581.880 1718.630 2586.480 1718.930 ;
        RECT 2581.880 1710.130 2586.480 1710.430 ;
        RECT 2581.880 1704.490 2586.480 1704.790 ;
        RECT 1575.460 1604.095 1577.200 1605.000 ;
        RECT 1397.545 1603.930 1397.875 1603.945 ;
        RECT 1397.545 1603.615 1398.090 1603.930 ;
      LAYER met3 ;
        RECT 305.055 1602.215 1395.530 1603.080 ;
      LAYER met3 ;
        RECT 1397.790 1602.680 1398.090 1603.615 ;
        RECT 1395.930 1602.080 1399.930 1602.680 ;
      LAYER met3 ;
        RECT 1555.055 1496.480 2645.530 1497.345 ;
      LAYER met3 ;
        RECT 2645.930 1496.880 2649.930 1497.480 ;
      LAYER met3 ;
        RECT 1555.055 1493.120 2645.930 1496.480 ;
        RECT 1555.055 1491.720 2645.530 1493.120 ;
      LAYER met3 ;
        RECT 2645.930 1492.120 2649.930 1492.720 ;
      LAYER met3 ;
        RECT 1555.055 1487.680 2645.930 1491.720 ;
        RECT 1555.055 1486.280 2645.530 1487.680 ;
      LAYER met3 ;
        RECT 2645.930 1486.680 2649.930 1487.280 ;
      LAYER met3 ;
        RECT 1555.055 1482.920 2645.930 1486.280 ;
        RECT 1555.055 1481.520 2645.530 1482.920 ;
      LAYER met3 ;
        RECT 2645.930 1481.920 2649.930 1482.520 ;
      LAYER met3 ;
        RECT 1555.055 1477.480 2645.930 1481.520 ;
        RECT 1555.055 1476.080 2645.530 1477.480 ;
      LAYER met3 ;
        RECT 2645.930 1476.480 2649.930 1477.080 ;
      LAYER met3 ;
        RECT 1555.055 1472.720 2645.930 1476.080 ;
        RECT 1555.055 1471.320 2645.530 1472.720 ;
      LAYER met3 ;
        RECT 2645.930 1471.720 2649.930 1472.320 ;
      LAYER met3 ;
        RECT 1555.055 1467.960 2645.930 1471.320 ;
        RECT 1555.055 1466.560 2645.530 1467.960 ;
      LAYER met3 ;
        RECT 2645.930 1466.960 2649.930 1467.560 ;
      LAYER met3 ;
        RECT 1555.055 1462.520 2645.930 1466.560 ;
        RECT 1555.055 1461.120 2645.530 1462.520 ;
      LAYER met3 ;
        RECT 2645.930 1461.520 2649.930 1462.120 ;
      LAYER met3 ;
        RECT 1555.055 1457.760 2645.930 1461.120 ;
        RECT 1555.055 1456.360 2645.530 1457.760 ;
      LAYER met3 ;
        RECT 2645.930 1456.760 2649.930 1457.360 ;
      LAYER met3 ;
        RECT 1555.055 1452.320 2645.930 1456.360 ;
        RECT 1555.055 1450.920 2645.530 1452.320 ;
      LAYER met3 ;
        RECT 2645.930 1451.320 2649.930 1451.920 ;
      LAYER met3 ;
        RECT 1555.055 1447.560 2645.930 1450.920 ;
        RECT 1555.055 1446.160 2645.530 1447.560 ;
      LAYER met3 ;
        RECT 2645.930 1446.560 2649.930 1447.160 ;
      LAYER met3 ;
        RECT 1555.055 1442.120 2645.930 1446.160 ;
        RECT 1555.055 1440.720 2645.530 1442.120 ;
      LAYER met3 ;
        RECT 2645.930 1441.120 2649.930 1441.720 ;
      LAYER met3 ;
        RECT 1555.055 1437.360 2645.930 1440.720 ;
        RECT 1555.055 1435.960 2645.530 1437.360 ;
      LAYER met3 ;
        RECT 2645.930 1436.360 2649.930 1436.960 ;
      LAYER met3 ;
        RECT 1555.055 1432.600 2645.930 1435.960 ;
        RECT 1555.055 1431.200 2645.530 1432.600 ;
      LAYER met3 ;
        RECT 2645.930 1431.600 2649.930 1432.200 ;
      LAYER met3 ;
        RECT 1555.055 1427.160 2645.930 1431.200 ;
        RECT 1555.055 1425.760 2645.530 1427.160 ;
      LAYER met3 ;
        RECT 2645.930 1426.160 2649.930 1426.760 ;
      LAYER met3 ;
        RECT 1555.055 1422.400 2645.930 1425.760 ;
        RECT 1555.055 1421.000 2645.530 1422.400 ;
      LAYER met3 ;
        RECT 2645.930 1421.400 2649.930 1422.000 ;
      LAYER met3 ;
        RECT 1555.055 1416.960 2645.930 1421.000 ;
        RECT 1555.055 1415.560 2645.530 1416.960 ;
      LAYER met3 ;
        RECT 2645.930 1415.960 2649.930 1416.560 ;
      LAYER met3 ;
        RECT 1555.055 1412.200 2645.930 1415.560 ;
        RECT 1555.055 1410.800 2645.530 1412.200 ;
      LAYER met3 ;
        RECT 2645.930 1411.200 2649.930 1411.800 ;
      LAYER met3 ;
        RECT 1555.055 1406.760 2645.930 1410.800 ;
        RECT 1555.055 1405.360 2645.530 1406.760 ;
      LAYER met3 ;
        RECT 2645.930 1405.760 2649.930 1406.360 ;
      LAYER met3 ;
        RECT 1555.055 1402.000 2645.930 1405.360 ;
        RECT 1555.055 1400.600 2645.530 1402.000 ;
      LAYER met3 ;
        RECT 2645.930 1401.000 2649.930 1401.600 ;
      LAYER met3 ;
        RECT 1555.055 1397.240 2645.930 1400.600 ;
        RECT 1555.055 1395.840 2645.530 1397.240 ;
      LAYER met3 ;
        RECT 2645.930 1396.240 2649.930 1396.840 ;
      LAYER met3 ;
        RECT 1555.055 1391.800 2645.930 1395.840 ;
        RECT 1555.055 1390.400 2645.530 1391.800 ;
      LAYER met3 ;
        RECT 2645.930 1390.800 2649.930 1391.400 ;
      LAYER met3 ;
        RECT 1555.055 1387.040 2645.930 1390.400 ;
        RECT 1555.055 1385.640 2645.530 1387.040 ;
      LAYER met3 ;
        RECT 2645.930 1386.040 2649.930 1386.640 ;
      LAYER met3 ;
        RECT 1555.055 1381.600 2645.930 1385.640 ;
        RECT 1555.055 1380.200 2645.530 1381.600 ;
      LAYER met3 ;
        RECT 2645.930 1380.600 2649.930 1381.200 ;
      LAYER met3 ;
        RECT 1555.055 1376.840 2645.930 1380.200 ;
        RECT 1555.055 1375.440 2645.530 1376.840 ;
      LAYER met3 ;
        RECT 2645.930 1375.840 2649.930 1376.440 ;
      LAYER met3 ;
        RECT 1555.055 1372.080 2645.930 1375.440 ;
        RECT 1555.055 1370.680 2645.530 1372.080 ;
      LAYER met3 ;
        RECT 2645.930 1371.080 2649.930 1371.680 ;
      LAYER met3 ;
        RECT 1555.055 1366.640 2645.930 1370.680 ;
        RECT 1555.055 1365.240 2645.530 1366.640 ;
      LAYER met3 ;
        RECT 2645.930 1365.640 2649.930 1366.240 ;
      LAYER met3 ;
        RECT 1555.055 1361.880 2645.930 1365.240 ;
        RECT 1555.055 1360.480 2645.530 1361.880 ;
      LAYER met3 ;
        RECT 2645.930 1360.880 2649.930 1361.480 ;
      LAYER met3 ;
        RECT 1555.055 1356.440 2645.930 1360.480 ;
        RECT 1555.055 1355.040 2645.530 1356.440 ;
      LAYER met3 ;
        RECT 2645.930 1355.440 2649.930 1356.040 ;
      LAYER met3 ;
        RECT 1555.055 1351.680 2645.930 1355.040 ;
        RECT 1555.055 1350.280 2645.530 1351.680 ;
      LAYER met3 ;
        RECT 2645.930 1350.680 2649.930 1351.280 ;
      LAYER met3 ;
        RECT 1555.055 1346.240 2645.930 1350.280 ;
        RECT 1555.055 1344.840 2645.530 1346.240 ;
      LAYER met3 ;
        RECT 2645.930 1345.240 2649.930 1345.840 ;
      LAYER met3 ;
        RECT 1555.055 1341.480 2645.930 1344.840 ;
        RECT 1555.055 1340.080 2645.530 1341.480 ;
      LAYER met3 ;
        RECT 2645.930 1340.480 2649.930 1341.080 ;
      LAYER met3 ;
        RECT 1555.055 1336.720 2645.930 1340.080 ;
        RECT 1555.055 1335.320 2645.530 1336.720 ;
      LAYER met3 ;
        RECT 2645.930 1335.720 2649.930 1336.320 ;
      LAYER met3 ;
        RECT 1555.055 1331.280 2645.930 1335.320 ;
        RECT 1555.055 1329.880 2645.530 1331.280 ;
      LAYER met3 ;
        RECT 2645.930 1330.280 2649.930 1330.880 ;
      LAYER met3 ;
        RECT 1555.055 1326.520 2645.930 1329.880 ;
        RECT 1555.055 1325.120 2645.530 1326.520 ;
      LAYER met3 ;
        RECT 2645.930 1325.520 2649.930 1326.120 ;
      LAYER met3 ;
        RECT 1555.055 1321.080 2645.930 1325.120 ;
        RECT 1555.055 1319.680 2645.530 1321.080 ;
      LAYER met3 ;
        RECT 2645.930 1320.080 2649.930 1320.680 ;
      LAYER met3 ;
        RECT 1555.055 1316.320 2645.930 1319.680 ;
        RECT 1555.055 1314.920 2645.530 1316.320 ;
      LAYER met3 ;
        RECT 2645.930 1315.320 2649.930 1315.920 ;
      LAYER met3 ;
        RECT 1555.055 1310.880 2645.930 1314.920 ;
        RECT 1555.055 1309.480 2645.530 1310.880 ;
      LAYER met3 ;
        RECT 2645.930 1309.880 2649.930 1310.480 ;
      LAYER met3 ;
        RECT 1555.055 1306.120 2645.930 1309.480 ;
        RECT 1555.055 1304.720 2645.530 1306.120 ;
      LAYER met3 ;
        RECT 2645.930 1305.120 2649.930 1305.720 ;
      LAYER met3 ;
        RECT 1555.055 1301.360 2645.930 1304.720 ;
        RECT 1555.055 1299.960 2645.530 1301.360 ;
      LAYER met3 ;
        RECT 2645.930 1300.360 2649.930 1300.960 ;
      LAYER met3 ;
        RECT 1555.055 1295.920 2645.930 1299.960 ;
        RECT 1555.055 1294.520 2645.530 1295.920 ;
      LAYER met3 ;
        RECT 2645.930 1294.920 2649.930 1295.520 ;
      LAYER met3 ;
        RECT 1555.055 1291.160 2645.930 1294.520 ;
        RECT 1555.055 1289.760 2645.530 1291.160 ;
      LAYER met3 ;
        RECT 2645.930 1290.160 2649.930 1290.760 ;
      LAYER met3 ;
        RECT 1555.055 1285.720 2645.930 1289.760 ;
        RECT 1555.055 1284.320 2645.530 1285.720 ;
      LAYER met3 ;
        RECT 2645.930 1284.720 2649.930 1285.320 ;
      LAYER met3 ;
        RECT 1555.055 1280.960 2645.930 1284.320 ;
        RECT 1555.055 1279.560 2645.530 1280.960 ;
      LAYER met3 ;
        RECT 2645.930 1279.960 2649.930 1280.560 ;
      LAYER met3 ;
        RECT 1555.055 1276.200 2645.930 1279.560 ;
        RECT 1555.055 1274.800 2645.530 1276.200 ;
      LAYER met3 ;
        RECT 2645.930 1275.200 2649.930 1275.800 ;
      LAYER met3 ;
        RECT 1555.055 1270.760 2645.930 1274.800 ;
        RECT 1555.055 1269.360 2645.530 1270.760 ;
      LAYER met3 ;
        RECT 2645.930 1269.760 2649.930 1270.360 ;
      LAYER met3 ;
        RECT 1555.055 1266.000 2645.930 1269.360 ;
        RECT 1555.055 1264.600 2645.530 1266.000 ;
      LAYER met3 ;
        RECT 2645.930 1265.000 2649.930 1265.600 ;
      LAYER met3 ;
        RECT 1555.055 1260.560 2645.930 1264.600 ;
        RECT 1555.055 1259.160 2645.530 1260.560 ;
      LAYER met3 ;
        RECT 2645.930 1259.560 2649.930 1260.160 ;
      LAYER met3 ;
        RECT 1555.055 1255.800 2645.930 1259.160 ;
        RECT 1555.055 1254.400 2645.530 1255.800 ;
      LAYER met3 ;
        RECT 2645.930 1254.800 2649.930 1255.400 ;
      LAYER met3 ;
        RECT 1555.055 1250.360 2645.930 1254.400 ;
        RECT 1555.055 1248.960 2645.530 1250.360 ;
      LAYER met3 ;
        RECT 2645.930 1249.360 2649.930 1249.960 ;
      LAYER met3 ;
        RECT 1555.055 1245.600 2645.930 1248.960 ;
        RECT 1555.055 1244.200 2645.530 1245.600 ;
      LAYER met3 ;
        RECT 2645.930 1244.600 2649.930 1245.200 ;
      LAYER met3 ;
        RECT 1555.055 1240.840 2645.930 1244.200 ;
        RECT 1555.055 1239.440 2645.530 1240.840 ;
      LAYER met3 ;
        RECT 2645.930 1239.840 2649.930 1240.440 ;
      LAYER met3 ;
        RECT 1555.055 1235.400 2645.930 1239.440 ;
        RECT 1555.055 1234.000 2645.530 1235.400 ;
      LAYER met3 ;
        RECT 2645.930 1234.400 2649.930 1235.000 ;
      LAYER met3 ;
        RECT 1555.055 1230.640 2645.930 1234.000 ;
        RECT 1555.055 1229.240 2645.530 1230.640 ;
      LAYER met3 ;
        RECT 2645.930 1229.640 2649.930 1230.240 ;
      LAYER met3 ;
        RECT 1555.055 1225.200 2645.930 1229.240 ;
        RECT 1555.055 1223.800 2645.530 1225.200 ;
      LAYER met3 ;
        RECT 2645.930 1224.200 2649.930 1224.800 ;
      LAYER met3 ;
        RECT 1555.055 1220.440 2645.930 1223.800 ;
        RECT 1555.055 1219.040 2645.530 1220.440 ;
      LAYER met3 ;
        RECT 2645.930 1219.440 2649.930 1220.040 ;
      LAYER met3 ;
        RECT 1555.055 1215.000 2645.930 1219.040 ;
        RECT 1555.055 1213.600 2645.530 1215.000 ;
      LAYER met3 ;
        RECT 2645.930 1214.000 2649.930 1214.600 ;
      LAYER met3 ;
        RECT 1555.055 1210.240 2645.930 1213.600 ;
        RECT 1555.055 1208.840 2645.530 1210.240 ;
      LAYER met3 ;
        RECT 2645.930 1209.240 2649.930 1209.840 ;
      LAYER met3 ;
        RECT 1555.055 1205.480 2645.930 1208.840 ;
        RECT 1555.055 1204.080 2645.530 1205.480 ;
      LAYER met3 ;
        RECT 2645.930 1204.480 2649.930 1205.080 ;
      LAYER met3 ;
        RECT 1555.055 1200.040 2645.930 1204.080 ;
        RECT 1555.055 1198.640 2645.530 1200.040 ;
      LAYER met3 ;
        RECT 2645.930 1199.040 2649.930 1199.640 ;
      LAYER met3 ;
        RECT 1555.055 1195.280 2645.930 1198.640 ;
        RECT 1555.055 1193.880 2645.530 1195.280 ;
      LAYER met3 ;
        RECT 2645.930 1194.280 2649.930 1194.880 ;
      LAYER met3 ;
        RECT 1555.055 1189.840 2645.930 1193.880 ;
        RECT 1555.055 1188.440 2645.530 1189.840 ;
      LAYER met3 ;
        RECT 2645.930 1188.840 2649.930 1189.440 ;
      LAYER met3 ;
        RECT 1555.055 1185.080 2645.930 1188.440 ;
        RECT 1555.055 1183.680 2645.530 1185.080 ;
      LAYER met3 ;
        RECT 2645.930 1184.080 2649.930 1184.680 ;
      LAYER met3 ;
        RECT 1555.055 1179.640 2645.930 1183.680 ;
        RECT 1555.055 1178.240 2645.530 1179.640 ;
      LAYER met3 ;
        RECT 2645.930 1178.640 2649.930 1179.240 ;
      LAYER met3 ;
        RECT 1555.055 1174.880 2645.930 1178.240 ;
        RECT 1555.055 1173.480 2645.530 1174.880 ;
      LAYER met3 ;
        RECT 2645.930 1173.880 2649.930 1174.480 ;
      LAYER met3 ;
        RECT 1555.055 1170.120 2645.930 1173.480 ;
        RECT 1555.055 1168.720 2645.530 1170.120 ;
      LAYER met3 ;
        RECT 2645.930 1169.120 2649.930 1169.720 ;
      LAYER met3 ;
        RECT 1555.055 1164.680 2645.930 1168.720 ;
        RECT 1555.055 1163.280 2645.530 1164.680 ;
      LAYER met3 ;
        RECT 2645.930 1163.680 2649.930 1164.280 ;
      LAYER met3 ;
        RECT 1555.055 1159.920 2645.930 1163.280 ;
        RECT 1555.055 1158.520 2645.530 1159.920 ;
      LAYER met3 ;
        RECT 2645.930 1158.920 2649.930 1159.520 ;
      LAYER met3 ;
        RECT 1555.055 1154.480 2645.930 1158.520 ;
        RECT 1555.055 1153.080 2645.530 1154.480 ;
      LAYER met3 ;
        RECT 2645.930 1153.480 2649.930 1154.080 ;
      LAYER met3 ;
        RECT 1555.055 1149.720 2645.930 1153.080 ;
        RECT 1555.055 1148.320 2645.530 1149.720 ;
      LAYER met3 ;
        RECT 2645.930 1148.720 2649.930 1149.320 ;
      LAYER met3 ;
        RECT 1555.055 1144.960 2645.930 1148.320 ;
        RECT 1555.055 1143.560 2645.530 1144.960 ;
      LAYER met3 ;
        RECT 2645.930 1143.960 2649.930 1144.560 ;
      LAYER met3 ;
        RECT 1555.055 1139.520 2645.930 1143.560 ;
        RECT 1555.055 1138.120 2645.530 1139.520 ;
      LAYER met3 ;
        RECT 2645.930 1138.520 2649.930 1139.120 ;
      LAYER met3 ;
        RECT 1555.055 1134.760 2645.930 1138.120 ;
        RECT 1555.055 1133.360 2645.530 1134.760 ;
      LAYER met3 ;
        RECT 2645.930 1133.760 2649.930 1134.360 ;
      LAYER met3 ;
        RECT 1555.055 1129.320 2645.930 1133.360 ;
        RECT 1555.055 1127.920 2645.530 1129.320 ;
      LAYER met3 ;
        RECT 2645.930 1128.320 2649.930 1128.920 ;
      LAYER met3 ;
        RECT 1555.055 1124.560 2645.930 1127.920 ;
        RECT 1555.055 1123.160 2645.530 1124.560 ;
      LAYER met3 ;
        RECT 2645.930 1123.560 2649.930 1124.160 ;
      LAYER met3 ;
        RECT 1555.055 1119.120 2645.930 1123.160 ;
        RECT 1555.055 1117.720 2645.530 1119.120 ;
      LAYER met3 ;
        RECT 2645.930 1118.120 2649.930 1118.720 ;
      LAYER met3 ;
        RECT 1555.055 1114.360 2645.930 1117.720 ;
        RECT 1555.055 1112.960 2645.530 1114.360 ;
      LAYER met3 ;
        RECT 2645.930 1113.360 2649.930 1113.960 ;
      LAYER met3 ;
        RECT 1555.055 1109.600 2645.930 1112.960 ;
        RECT 1555.055 1108.200 2645.530 1109.600 ;
      LAYER met3 ;
        RECT 2645.930 1108.600 2649.930 1109.200 ;
      LAYER met3 ;
        RECT 1555.055 1104.160 2645.930 1108.200 ;
        RECT 1555.055 1102.760 2645.530 1104.160 ;
      LAYER met3 ;
        RECT 2645.930 1103.160 2649.930 1103.760 ;
      LAYER met3 ;
        RECT 1555.055 1099.400 2645.930 1102.760 ;
        RECT 1555.055 1098.000 2645.530 1099.400 ;
      LAYER met3 ;
        RECT 2645.930 1098.400 2649.930 1099.000 ;
      LAYER met3 ;
        RECT 1555.055 1093.960 2645.930 1098.000 ;
        RECT 1555.055 1092.560 2645.530 1093.960 ;
      LAYER met3 ;
        RECT 2645.930 1092.960 2649.930 1093.560 ;
      LAYER met3 ;
        RECT 1555.055 1089.200 2645.930 1092.560 ;
        RECT 1555.055 1087.800 2645.530 1089.200 ;
      LAYER met3 ;
        RECT 2645.930 1088.200 2649.930 1088.800 ;
      LAYER met3 ;
        RECT 1555.055 1083.760 2645.930 1087.800 ;
        RECT 1555.055 1082.360 2645.530 1083.760 ;
      LAYER met3 ;
        RECT 2645.930 1082.760 2649.930 1083.360 ;
      LAYER met3 ;
        RECT 1555.055 1079.000 2645.930 1082.360 ;
        RECT 1555.055 1077.600 2645.530 1079.000 ;
      LAYER met3 ;
        RECT 2645.930 1078.000 2649.930 1078.600 ;
      LAYER met3 ;
        RECT 1555.055 1074.240 2645.930 1077.600 ;
        RECT 1555.055 1072.840 2645.530 1074.240 ;
      LAYER met3 ;
        RECT 2645.930 1073.240 2649.930 1073.840 ;
      LAYER met3 ;
        RECT 1555.055 1068.800 2645.930 1072.840 ;
        RECT 1555.055 1067.400 2645.530 1068.800 ;
      LAYER met3 ;
        RECT 2645.930 1067.800 2649.930 1068.400 ;
      LAYER met3 ;
        RECT 1555.055 1064.040 2645.930 1067.400 ;
        RECT 1555.055 1062.640 2645.530 1064.040 ;
      LAYER met3 ;
        RECT 2645.930 1063.040 2649.930 1063.640 ;
      LAYER met3 ;
        RECT 1555.055 1058.600 2645.930 1062.640 ;
        RECT 1555.055 1057.200 2645.530 1058.600 ;
      LAYER met3 ;
        RECT 2645.930 1057.600 2649.930 1058.200 ;
      LAYER met3 ;
        RECT 1555.055 1053.840 2645.930 1057.200 ;
        RECT 1555.055 1052.440 2645.530 1053.840 ;
      LAYER met3 ;
        RECT 2645.930 1052.840 2649.930 1053.440 ;
      LAYER met3 ;
        RECT 1555.055 1049.080 2645.930 1052.440 ;
        RECT 1555.055 1047.680 2645.530 1049.080 ;
      LAYER met3 ;
        RECT 2645.930 1048.080 2649.930 1048.680 ;
      LAYER met3 ;
        RECT 1555.055 1043.640 2645.930 1047.680 ;
        RECT 1555.055 1042.240 2645.530 1043.640 ;
      LAYER met3 ;
        RECT 2645.930 1042.640 2649.930 1043.240 ;
      LAYER met3 ;
        RECT 1555.055 1038.880 2645.930 1042.240 ;
        RECT 1555.055 1037.480 2645.530 1038.880 ;
      LAYER met3 ;
        RECT 2645.930 1037.880 2649.930 1038.480 ;
      LAYER met3 ;
        RECT 1555.055 1033.440 2645.930 1037.480 ;
        RECT 1555.055 1032.040 2645.530 1033.440 ;
      LAYER met3 ;
        RECT 2645.930 1032.440 2649.930 1033.040 ;
      LAYER met3 ;
        RECT 1555.055 1028.680 2645.930 1032.040 ;
        RECT 1555.055 1027.280 2645.530 1028.680 ;
      LAYER met3 ;
        RECT 2645.930 1027.680 2649.930 1028.280 ;
      LAYER met3 ;
        RECT 1555.055 1023.240 2645.930 1027.280 ;
        RECT 1555.055 1021.840 2645.530 1023.240 ;
      LAYER met3 ;
        RECT 2645.930 1022.240 2649.930 1022.840 ;
      LAYER met3 ;
        RECT 1555.055 1018.480 2645.930 1021.840 ;
        RECT 1555.055 1017.080 2645.530 1018.480 ;
      LAYER met3 ;
        RECT 2645.930 1017.480 2649.930 1018.080 ;
      LAYER met3 ;
        RECT 1555.055 1013.720 2645.930 1017.080 ;
        RECT 1555.055 1012.320 2645.530 1013.720 ;
      LAYER met3 ;
        RECT 2645.930 1012.720 2649.930 1013.320 ;
      LAYER met3 ;
        RECT 1555.055 1008.280 2645.930 1012.320 ;
        RECT 1555.055 1006.880 2645.530 1008.280 ;
      LAYER met3 ;
        RECT 2645.930 1007.280 2649.930 1007.880 ;
      LAYER met3 ;
        RECT 1555.055 1003.520 2645.930 1006.880 ;
        RECT 1555.055 1002.120 2645.530 1003.520 ;
      LAYER met3 ;
        RECT 2645.930 1002.520 2649.930 1003.120 ;
      LAYER met3 ;
        RECT 1555.055 998.080 2645.930 1002.120 ;
        RECT 1555.055 996.680 2645.530 998.080 ;
      LAYER met3 ;
        RECT 2645.930 997.080 2649.930 997.680 ;
      LAYER met3 ;
        RECT 1555.055 993.320 2645.930 996.680 ;
        RECT 1555.055 991.920 2645.530 993.320 ;
      LAYER met3 ;
        RECT 2645.930 992.320 2649.930 992.920 ;
      LAYER met3 ;
        RECT 1555.055 987.880 2645.930 991.920 ;
        RECT 1555.055 986.480 2645.530 987.880 ;
      LAYER met3 ;
        RECT 2645.930 986.880 2649.930 987.480 ;
      LAYER met3 ;
        RECT 1555.055 983.120 2645.930 986.480 ;
        RECT 1555.055 981.720 2645.530 983.120 ;
      LAYER met3 ;
        RECT 2645.930 982.120 2649.930 982.720 ;
      LAYER met3 ;
        RECT 1555.055 978.360 2645.930 981.720 ;
        RECT 1555.055 976.960 2645.530 978.360 ;
      LAYER met3 ;
        RECT 2645.930 977.360 2649.930 977.960 ;
      LAYER met3 ;
        RECT 1555.055 972.920 2645.930 976.960 ;
        RECT 1555.055 971.520 2645.530 972.920 ;
      LAYER met3 ;
        RECT 2645.930 971.920 2649.930 972.520 ;
      LAYER met3 ;
        RECT 1555.055 968.160 2645.930 971.520 ;
        RECT 1555.055 966.760 2645.530 968.160 ;
      LAYER met3 ;
        RECT 2645.930 967.160 2649.930 967.760 ;
      LAYER met3 ;
        RECT 1555.055 962.720 2645.930 966.760 ;
        RECT 1555.055 961.320 2645.530 962.720 ;
      LAYER met3 ;
        RECT 2645.930 961.720 2649.930 962.320 ;
      LAYER met3 ;
        RECT 1555.055 957.960 2645.930 961.320 ;
        RECT 1555.055 956.560 2645.530 957.960 ;
      LAYER met3 ;
        RECT 2645.930 956.960 2649.930 957.560 ;
      LAYER met3 ;
        RECT 1555.055 953.200 2645.930 956.560 ;
        RECT 1555.055 951.800 2645.530 953.200 ;
      LAYER met3 ;
        RECT 2645.930 952.200 2649.930 952.800 ;
      LAYER met3 ;
        RECT 1555.055 947.760 2645.930 951.800 ;
        RECT 1555.055 946.360 2645.530 947.760 ;
      LAYER met3 ;
        RECT 2645.930 946.760 2649.930 947.360 ;
      LAYER met3 ;
        RECT 1555.055 943.000 2645.930 946.360 ;
        RECT 1555.055 941.600 2645.530 943.000 ;
      LAYER met3 ;
        RECT 2645.930 942.000 2649.930 942.600 ;
      LAYER met3 ;
        RECT 1555.055 937.560 2645.930 941.600 ;
        RECT 1555.055 936.160 2645.530 937.560 ;
      LAYER met3 ;
        RECT 2645.930 936.560 2649.930 937.160 ;
      LAYER met3 ;
        RECT 1555.055 932.800 2645.930 936.160 ;
        RECT 1555.055 931.400 2645.530 932.800 ;
      LAYER met3 ;
        RECT 2645.930 931.800 2649.930 932.400 ;
      LAYER met3 ;
        RECT 1555.055 927.360 2645.930 931.400 ;
        RECT 1555.055 925.960 2645.530 927.360 ;
      LAYER met3 ;
        RECT 2645.930 926.360 2649.930 926.960 ;
      LAYER met3 ;
        RECT 1555.055 922.600 2645.930 925.960 ;
        RECT 1555.055 921.200 2645.530 922.600 ;
      LAYER met3 ;
        RECT 2645.930 921.600 2649.930 922.200 ;
      LAYER met3 ;
        RECT 1555.055 917.840 2645.930 921.200 ;
        RECT 1555.055 916.440 2645.530 917.840 ;
      LAYER met3 ;
        RECT 2645.930 916.840 2649.930 917.440 ;
      LAYER met3 ;
        RECT 1555.055 912.400 2645.930 916.440 ;
        RECT 1555.055 911.000 2645.530 912.400 ;
      LAYER met3 ;
        RECT 2645.930 911.400 2649.930 912.000 ;
      LAYER met3 ;
        RECT 1555.055 907.640 2645.930 911.000 ;
        RECT 1555.055 906.240 2645.530 907.640 ;
      LAYER met3 ;
        RECT 2645.930 906.640 2649.930 907.240 ;
      LAYER met3 ;
        RECT 1555.055 902.200 2645.930 906.240 ;
        RECT 1555.055 900.800 2645.530 902.200 ;
      LAYER met3 ;
        RECT 2645.930 901.200 2649.930 901.800 ;
      LAYER met3 ;
        RECT 1555.055 897.440 2645.930 900.800 ;
        RECT 1555.055 896.040 2645.530 897.440 ;
      LAYER met3 ;
        RECT 2645.930 896.440 2649.930 897.040 ;
      LAYER met3 ;
        RECT 1555.055 892.000 2645.930 896.040 ;
        RECT 1555.055 890.600 2645.530 892.000 ;
      LAYER met3 ;
        RECT 2645.930 891.000 2649.930 891.600 ;
      LAYER met3 ;
        RECT 1555.055 887.240 2645.930 890.600 ;
        RECT 1555.055 885.840 2645.530 887.240 ;
      LAYER met3 ;
        RECT 2645.930 886.240 2649.930 886.840 ;
      LAYER met3 ;
        RECT 1555.055 882.480 2645.930 885.840 ;
        RECT 1555.055 881.080 2645.530 882.480 ;
      LAYER met3 ;
        RECT 2645.930 881.480 2649.930 882.080 ;
      LAYER met3 ;
        RECT 1555.055 877.040 2645.930 881.080 ;
        RECT 1555.055 875.640 2645.530 877.040 ;
      LAYER met3 ;
        RECT 2645.930 876.040 2649.930 876.640 ;
      LAYER met3 ;
        RECT 1555.055 872.280 2645.930 875.640 ;
        RECT 1555.055 870.880 2645.530 872.280 ;
      LAYER met3 ;
        RECT 2645.930 871.280 2649.930 871.880 ;
      LAYER met3 ;
        RECT 1555.055 866.840 2645.930 870.880 ;
        RECT 1555.055 865.440 2645.530 866.840 ;
      LAYER met3 ;
        RECT 2645.930 865.840 2649.930 866.440 ;
      LAYER met3 ;
        RECT 1555.055 862.080 2645.930 865.440 ;
        RECT 1555.055 860.680 2645.530 862.080 ;
      LAYER met3 ;
        RECT 2645.930 861.080 2649.930 861.680 ;
      LAYER met3 ;
        RECT 1555.055 856.640 2645.930 860.680 ;
        RECT 1555.055 855.240 2645.530 856.640 ;
      LAYER met3 ;
        RECT 2645.930 855.640 2649.930 856.240 ;
      LAYER met3 ;
        RECT 1555.055 851.880 2645.930 855.240 ;
        RECT 1555.055 850.480 2645.530 851.880 ;
      LAYER met3 ;
        RECT 2645.930 850.880 2649.930 851.480 ;
      LAYER met3 ;
        RECT 1555.055 847.120 2645.930 850.480 ;
        RECT 1555.055 845.720 2645.530 847.120 ;
      LAYER met3 ;
        RECT 2645.930 846.120 2649.930 846.720 ;
      LAYER met3 ;
        RECT 1555.055 841.680 2645.930 845.720 ;
        RECT 1555.055 840.280 2645.530 841.680 ;
      LAYER met3 ;
        RECT 2645.930 840.680 2649.930 841.280 ;
      LAYER met3 ;
        RECT 1555.055 836.920 2645.930 840.280 ;
        RECT 1555.055 835.520 2645.530 836.920 ;
      LAYER met3 ;
        RECT 2645.930 835.920 2649.930 836.520 ;
      LAYER met3 ;
        RECT 1555.055 831.480 2645.930 835.520 ;
        RECT 1555.055 830.080 2645.530 831.480 ;
      LAYER met3 ;
        RECT 2645.930 830.480 2649.930 831.080 ;
      LAYER met3 ;
        RECT 1555.055 826.720 2645.930 830.080 ;
        RECT 1555.055 825.320 2645.530 826.720 ;
      LAYER met3 ;
        RECT 2645.930 825.720 2649.930 826.320 ;
      LAYER met3 ;
        RECT 1555.055 821.960 2645.930 825.320 ;
        RECT 1555.055 820.560 2645.530 821.960 ;
      LAYER met3 ;
        RECT 2645.930 820.960 2649.930 821.560 ;
      LAYER met3 ;
        RECT 1555.055 816.520 2645.930 820.560 ;
        RECT 1555.055 815.120 2645.530 816.520 ;
      LAYER met3 ;
        RECT 2645.930 815.520 2649.930 816.120 ;
      LAYER met3 ;
        RECT 1555.055 811.760 2645.930 815.120 ;
        RECT 1555.055 810.360 2645.530 811.760 ;
      LAYER met3 ;
        RECT 2645.930 810.760 2649.930 811.360 ;
      LAYER met3 ;
        RECT 1555.055 806.320 2645.930 810.360 ;
        RECT 1555.055 804.920 2645.530 806.320 ;
      LAYER met3 ;
        RECT 2645.930 805.320 2649.930 805.920 ;
      LAYER met3 ;
        RECT 1555.055 801.560 2645.930 804.920 ;
        RECT 1555.055 800.160 2645.530 801.560 ;
      LAYER met3 ;
        RECT 2645.930 800.560 2649.930 801.160 ;
      LAYER met3 ;
        RECT 1555.055 796.120 2645.930 800.160 ;
        RECT 1555.055 794.720 2645.530 796.120 ;
      LAYER met3 ;
        RECT 2645.930 795.120 2649.930 795.720 ;
      LAYER met3 ;
        RECT 1555.055 791.360 2645.930 794.720 ;
        RECT 1555.055 789.960 2645.530 791.360 ;
      LAYER met3 ;
        RECT 2645.930 790.360 2649.930 790.960 ;
      LAYER met3 ;
        RECT 1555.055 786.600 2645.930 789.960 ;
        RECT 1555.055 785.200 2645.530 786.600 ;
      LAYER met3 ;
        RECT 2645.930 785.600 2649.930 786.200 ;
      LAYER met3 ;
        RECT 1555.055 781.160 2645.930 785.200 ;
        RECT 1555.055 779.760 2645.530 781.160 ;
      LAYER met3 ;
        RECT 2645.930 780.160 2649.930 780.760 ;
      LAYER met3 ;
        RECT 1555.055 776.400 2645.930 779.760 ;
        RECT 1555.055 775.000 2645.530 776.400 ;
      LAYER met3 ;
        RECT 2645.930 775.400 2649.930 776.000 ;
      LAYER met3 ;
        RECT 1555.055 770.960 2645.930 775.000 ;
        RECT 1555.055 769.560 2645.530 770.960 ;
      LAYER met3 ;
        RECT 2645.930 769.960 2649.930 770.560 ;
      LAYER met3 ;
        RECT 1555.055 766.200 2645.930 769.560 ;
        RECT 1555.055 764.800 2645.530 766.200 ;
      LAYER met3 ;
        RECT 2645.930 765.200 2649.930 765.800 ;
      LAYER met3 ;
        RECT 1555.055 760.760 2645.930 764.800 ;
        RECT 1555.055 759.360 2645.530 760.760 ;
      LAYER met3 ;
        RECT 2645.930 759.760 2649.930 760.360 ;
      LAYER met3 ;
        RECT 1555.055 756.000 2645.930 759.360 ;
        RECT 1555.055 754.600 2645.530 756.000 ;
      LAYER met3 ;
        RECT 2645.930 755.000 2649.930 755.600 ;
      LAYER met3 ;
        RECT 1555.055 751.240 2645.930 754.600 ;
        RECT 1555.055 749.840 2645.530 751.240 ;
      LAYER met3 ;
        RECT 2645.930 750.240 2649.930 750.840 ;
      LAYER met3 ;
        RECT 1555.055 745.800 2645.930 749.840 ;
        RECT 1555.055 744.400 2645.530 745.800 ;
      LAYER met3 ;
        RECT 2645.930 744.800 2649.930 745.400 ;
      LAYER met3 ;
        RECT 1555.055 741.040 2645.930 744.400 ;
        RECT 1555.055 739.640 2645.530 741.040 ;
      LAYER met3 ;
        RECT 2645.930 740.040 2649.930 740.640 ;
      LAYER met3 ;
        RECT 1555.055 735.600 2645.930 739.640 ;
        RECT 1555.055 734.200 2645.530 735.600 ;
      LAYER met3 ;
        RECT 2645.930 734.600 2649.930 735.200 ;
      LAYER met3 ;
        RECT 1555.055 730.840 2645.930 734.200 ;
        RECT 1555.055 729.440 2645.530 730.840 ;
      LAYER met3 ;
        RECT 2645.930 729.840 2649.930 730.440 ;
      LAYER met3 ;
        RECT 1555.055 726.080 2645.930 729.440 ;
        RECT 1555.055 724.680 2645.530 726.080 ;
      LAYER met3 ;
        RECT 2645.930 725.080 2649.930 725.680 ;
      LAYER met3 ;
        RECT 1555.055 720.640 2645.930 724.680 ;
        RECT 1555.055 719.240 2645.530 720.640 ;
      LAYER met3 ;
        RECT 2645.930 719.640 2649.930 720.240 ;
      LAYER met3 ;
        RECT 1555.055 715.880 2645.930 719.240 ;
        RECT 1555.055 714.480 2645.530 715.880 ;
      LAYER met3 ;
        RECT 2645.930 714.880 2649.930 715.480 ;
      LAYER met3 ;
        RECT 1555.055 710.440 2645.930 714.480 ;
        RECT 1555.055 709.040 2645.530 710.440 ;
      LAYER met3 ;
        RECT 2645.930 709.440 2649.930 710.040 ;
      LAYER met3 ;
        RECT 1555.055 705.680 2645.930 709.040 ;
        RECT 1555.055 704.280 2645.530 705.680 ;
      LAYER met3 ;
        RECT 2645.930 704.680 2649.930 705.280 ;
      LAYER met3 ;
        RECT 1555.055 700.240 2645.930 704.280 ;
        RECT 1555.055 698.840 2645.530 700.240 ;
      LAYER met3 ;
        RECT 2645.930 699.240 2649.930 699.840 ;
      LAYER met3 ;
        RECT 1555.055 695.480 2645.930 698.840 ;
        RECT 1555.055 694.080 2645.530 695.480 ;
      LAYER met3 ;
        RECT 2645.930 694.480 2649.930 695.080 ;
      LAYER met3 ;
        RECT 1555.055 690.720 2645.930 694.080 ;
        RECT 1555.055 689.320 2645.530 690.720 ;
      LAYER met3 ;
        RECT 2645.930 689.720 2649.930 690.320 ;
      LAYER met3 ;
        RECT 1555.055 685.280 2645.930 689.320 ;
        RECT 1555.055 683.880 2645.530 685.280 ;
      LAYER met3 ;
        RECT 2645.930 684.280 2649.930 684.880 ;
      LAYER met3 ;
        RECT 1555.055 680.520 2645.930 683.880 ;
        RECT 1555.055 679.120 2645.530 680.520 ;
      LAYER met3 ;
        RECT 2645.930 679.520 2649.930 680.120 ;
      LAYER met3 ;
        RECT 1555.055 675.080 2645.930 679.120 ;
        RECT 1555.055 673.680 2645.530 675.080 ;
      LAYER met3 ;
        RECT 2645.930 674.080 2649.930 674.680 ;
      LAYER met3 ;
        RECT 1555.055 670.320 2645.930 673.680 ;
        RECT 1555.055 668.920 2645.530 670.320 ;
      LAYER met3 ;
        RECT 2645.930 669.320 2649.930 669.920 ;
      LAYER met3 ;
        RECT 1555.055 664.880 2645.930 668.920 ;
        RECT 1555.055 663.480 2645.530 664.880 ;
      LAYER met3 ;
        RECT 2645.930 663.880 2649.930 664.480 ;
      LAYER met3 ;
        RECT 1555.055 660.120 2645.930 663.480 ;
        RECT 1555.055 658.720 2645.530 660.120 ;
      LAYER met3 ;
        RECT 2645.930 659.120 2649.930 659.720 ;
      LAYER met3 ;
        RECT 1555.055 655.360 2645.930 658.720 ;
        RECT 1555.055 653.960 2645.530 655.360 ;
      LAYER met3 ;
        RECT 2645.930 654.360 2649.930 654.960 ;
      LAYER met3 ;
        RECT 1555.055 649.920 2645.930 653.960 ;
        RECT 1555.055 648.520 2645.530 649.920 ;
      LAYER met3 ;
        RECT 2645.930 648.920 2649.930 649.520 ;
      LAYER met3 ;
        RECT 1555.055 645.160 2645.930 648.520 ;
        RECT 1555.055 643.760 2645.530 645.160 ;
      LAYER met3 ;
        RECT 2645.930 644.160 2649.930 644.760 ;
      LAYER met3 ;
        RECT 1555.055 639.720 2645.930 643.760 ;
        RECT 1555.055 638.320 2645.530 639.720 ;
      LAYER met3 ;
        RECT 2645.930 638.720 2649.930 639.320 ;
      LAYER met3 ;
        RECT 1555.055 634.960 2645.930 638.320 ;
        RECT 1555.055 633.560 2645.530 634.960 ;
      LAYER met3 ;
        RECT 2645.930 633.960 2649.930 634.560 ;
      LAYER met3 ;
        RECT 1555.055 629.520 2645.930 633.560 ;
        RECT 1555.055 628.120 2645.530 629.520 ;
      LAYER met3 ;
        RECT 2645.930 628.520 2649.930 629.120 ;
      LAYER met3 ;
        RECT 1555.055 624.760 2645.930 628.120 ;
        RECT 1555.055 623.360 2645.530 624.760 ;
      LAYER met3 ;
        RECT 2645.930 623.760 2649.930 624.360 ;
      LAYER met3 ;
        RECT 1555.055 620.000 2645.930 623.360 ;
        RECT 1555.055 618.600 2645.530 620.000 ;
      LAYER met3 ;
        RECT 2645.930 619.000 2649.930 619.600 ;
      LAYER met3 ;
        RECT 1555.055 614.560 2645.930 618.600 ;
        RECT 1555.055 613.160 2645.530 614.560 ;
      LAYER met3 ;
        RECT 2645.930 613.560 2649.930 614.160 ;
      LAYER met3 ;
        RECT 1555.055 609.800 2645.930 613.160 ;
        RECT 1555.055 608.400 2645.530 609.800 ;
      LAYER met3 ;
        RECT 2645.930 608.800 2649.930 609.400 ;
      LAYER met3 ;
        RECT 1555.055 604.360 2645.930 608.400 ;
        RECT 1555.055 602.960 2645.530 604.360 ;
      LAYER met3 ;
        RECT 2645.930 603.360 2649.930 603.960 ;
      LAYER met3 ;
        RECT 1555.055 599.600 2645.930 602.960 ;
        RECT 1555.055 598.200 2645.530 599.600 ;
      LAYER met3 ;
        RECT 2645.930 598.600 2649.930 599.200 ;
      LAYER met3 ;
        RECT 1555.055 594.840 2645.930 598.200 ;
        RECT 1555.055 593.440 2645.530 594.840 ;
      LAYER met3 ;
        RECT 2645.930 593.840 2649.930 594.440 ;
      LAYER met3 ;
        RECT 1555.055 589.400 2645.930 593.440 ;
        RECT 1555.055 588.000 2645.530 589.400 ;
      LAYER met3 ;
        RECT 2645.930 588.400 2649.930 589.000 ;
      LAYER met3 ;
        RECT 1555.055 584.640 2645.930 588.000 ;
        RECT 1555.055 583.240 2645.530 584.640 ;
      LAYER met3 ;
        RECT 2645.930 583.640 2649.930 584.240 ;
      LAYER met3 ;
        RECT 1555.055 579.200 2645.930 583.240 ;
        RECT 1555.055 577.800 2645.530 579.200 ;
      LAYER met3 ;
        RECT 2645.930 578.200 2649.930 578.800 ;
      LAYER met3 ;
        RECT 1555.055 574.440 2645.930 577.800 ;
        RECT 1555.055 573.040 2645.530 574.440 ;
      LAYER met3 ;
        RECT 2645.930 573.440 2649.930 574.040 ;
      LAYER met3 ;
        RECT 1555.055 569.000 2645.930 573.040 ;
        RECT 1555.055 567.600 2645.530 569.000 ;
      LAYER met3 ;
        RECT 2645.930 568.000 2649.930 568.600 ;
      LAYER met3 ;
        RECT 1555.055 564.240 2645.930 567.600 ;
        RECT 1555.055 562.840 2645.530 564.240 ;
      LAYER met3 ;
        RECT 2645.930 563.240 2649.930 563.840 ;
      LAYER met3 ;
        RECT 1555.055 559.480 2645.930 562.840 ;
        RECT 1555.055 558.080 2645.530 559.480 ;
      LAYER met3 ;
        RECT 2645.930 558.480 2649.930 559.080 ;
      LAYER met3 ;
        RECT 1555.055 554.040 2645.930 558.080 ;
        RECT 1555.055 552.640 2645.530 554.040 ;
      LAYER met3 ;
        RECT 2645.930 553.040 2649.930 553.640 ;
      LAYER met3 ;
        RECT 1555.055 549.280 2645.930 552.640 ;
        RECT 1555.055 547.880 2645.530 549.280 ;
      LAYER met3 ;
        RECT 2645.930 548.280 2649.930 548.880 ;
      LAYER met3 ;
        RECT 1555.055 543.840 2645.930 547.880 ;
        RECT 1555.055 542.440 2645.530 543.840 ;
      LAYER met3 ;
        RECT 2645.930 542.840 2649.930 543.440 ;
      LAYER met3 ;
        RECT 1555.055 539.080 2645.930 542.440 ;
        RECT 1555.055 537.680 2645.530 539.080 ;
      LAYER met3 ;
        RECT 2645.930 538.080 2649.930 538.680 ;
      LAYER met3 ;
        RECT 1555.055 533.640 2645.930 537.680 ;
        RECT 1555.055 532.240 2645.530 533.640 ;
      LAYER met3 ;
        RECT 2645.930 532.640 2649.930 533.240 ;
      LAYER met3 ;
        RECT 1555.055 528.880 2645.930 532.240 ;
        RECT 1555.055 527.480 2645.530 528.880 ;
      LAYER met3 ;
        RECT 2645.930 527.880 2649.930 528.480 ;
      LAYER met3 ;
        RECT 1555.055 524.120 2645.930 527.480 ;
        RECT 1555.055 522.720 2645.530 524.120 ;
      LAYER met3 ;
        RECT 2645.930 523.120 2649.930 523.720 ;
      LAYER met3 ;
        RECT 1555.055 518.680 2645.930 522.720 ;
        RECT 1555.055 517.280 2645.530 518.680 ;
      LAYER met3 ;
        RECT 2645.930 517.680 2649.930 518.280 ;
      LAYER met3 ;
        RECT 1555.055 513.920 2645.930 517.280 ;
        RECT 1555.055 512.520 2645.530 513.920 ;
      LAYER met3 ;
        RECT 2645.930 512.920 2649.930 513.520 ;
      LAYER met3 ;
        RECT 1555.055 508.480 2645.930 512.520 ;
        RECT 1555.055 507.080 2645.530 508.480 ;
      LAYER met3 ;
        RECT 2645.930 507.480 2649.930 508.080 ;
      LAYER met3 ;
        RECT 1555.055 503.720 2645.930 507.080 ;
        RECT 1555.055 502.320 2645.530 503.720 ;
      LAYER met3 ;
        RECT 2645.930 502.720 2649.930 503.320 ;
      LAYER met3 ;
        RECT 1555.055 498.960 2645.930 502.320 ;
        RECT 1555.055 497.560 2645.530 498.960 ;
      LAYER met3 ;
        RECT 2645.930 497.960 2649.930 498.560 ;
      LAYER met3 ;
        RECT 1555.055 493.520 2645.930 497.560 ;
        RECT 1555.055 492.120 2645.530 493.520 ;
      LAYER met3 ;
        RECT 2645.930 492.520 2649.930 493.120 ;
      LAYER met3 ;
        RECT 1555.055 488.760 2645.930 492.120 ;
        RECT 1555.055 487.360 2645.530 488.760 ;
      LAYER met3 ;
        RECT 2645.930 487.760 2649.930 488.360 ;
      LAYER met3 ;
        RECT 1555.055 483.320 2645.930 487.360 ;
        RECT 1555.055 481.920 2645.530 483.320 ;
      LAYER met3 ;
        RECT 2645.930 482.320 2649.930 482.920 ;
      LAYER met3 ;
        RECT 1555.055 478.560 2645.930 481.920 ;
        RECT 1555.055 477.160 2645.530 478.560 ;
      LAYER met3 ;
        RECT 2645.930 477.560 2649.930 478.160 ;
      LAYER met3 ;
        RECT 1555.055 473.120 2645.930 477.160 ;
        RECT 1555.055 471.720 2645.530 473.120 ;
      LAYER met3 ;
        RECT 2645.930 472.120 2649.930 472.720 ;
      LAYER met3 ;
        RECT 1555.055 468.360 2645.930 471.720 ;
        RECT 1555.055 466.960 2645.530 468.360 ;
      LAYER met3 ;
        RECT 2645.930 467.360 2649.930 467.960 ;
      LAYER met3 ;
        RECT 1555.055 463.600 2645.930 466.960 ;
        RECT 1555.055 462.200 2645.530 463.600 ;
      LAYER met3 ;
        RECT 2645.930 462.600 2649.930 463.200 ;
      LAYER met3 ;
        RECT 1555.055 458.160 2645.930 462.200 ;
        RECT 1555.055 456.760 2645.530 458.160 ;
      LAYER met3 ;
        RECT 2645.930 457.160 2649.930 457.760 ;
      LAYER met3 ;
        RECT 1555.055 453.400 2645.930 456.760 ;
        RECT 1555.055 452.000 2645.530 453.400 ;
      LAYER met3 ;
        RECT 2645.930 452.400 2649.930 453.000 ;
      LAYER met3 ;
        RECT 1555.055 447.960 2645.930 452.000 ;
        RECT 1555.055 446.560 2645.530 447.960 ;
      LAYER met3 ;
        RECT 2645.930 446.960 2649.930 447.560 ;
      LAYER met3 ;
        RECT 1555.055 443.200 2645.930 446.560 ;
        RECT 1555.055 441.800 2645.530 443.200 ;
      LAYER met3 ;
        RECT 2645.930 442.200 2649.930 442.800 ;
      LAYER met3 ;
        RECT 1555.055 437.760 2645.930 441.800 ;
        RECT 1555.055 436.360 2645.530 437.760 ;
      LAYER met3 ;
        RECT 2645.930 436.760 2649.930 437.360 ;
      LAYER met3 ;
        RECT 1555.055 433.000 2645.930 436.360 ;
        RECT 1555.055 431.600 2645.530 433.000 ;
      LAYER met3 ;
        RECT 2645.930 432.000 2649.930 432.600 ;
      LAYER met3 ;
        RECT 1555.055 428.240 2645.930 431.600 ;
        RECT 1555.055 426.840 2645.530 428.240 ;
      LAYER met3 ;
        RECT 2645.930 427.240 2649.930 427.840 ;
      LAYER met3 ;
        RECT 1555.055 422.800 2645.930 426.840 ;
        RECT 1555.055 421.400 2645.530 422.800 ;
      LAYER met3 ;
        RECT 2645.930 421.800 2649.930 422.400 ;
      LAYER met3 ;
        RECT 1555.055 418.040 2645.930 421.400 ;
        RECT 1555.055 416.640 2645.530 418.040 ;
      LAYER met3 ;
        RECT 2645.930 417.040 2649.930 417.640 ;
      LAYER met3 ;
        RECT 1555.055 412.600 2645.930 416.640 ;
        RECT 1555.055 411.200 2645.530 412.600 ;
      LAYER met3 ;
        RECT 2645.930 411.600 2649.930 412.200 ;
      LAYER met3 ;
        RECT 1555.055 407.840 2645.930 411.200 ;
        RECT 1555.055 406.440 2645.530 407.840 ;
      LAYER met3 ;
        RECT 2645.930 406.840 2649.930 407.440 ;
      LAYER met3 ;
        RECT 1555.055 403.080 2645.930 406.440 ;
        RECT 1555.055 402.215 2645.530 403.080 ;
      LAYER met3 ;
        RECT 2645.930 402.080 2649.930 402.680 ;
      LAYER via3 ;
        RECT 646.140 3264.180 646.460 3264.500 ;
        RECT 668.220 3264.180 668.540 3264.500 ;
        RECT 1292.900 3264.180 1293.220 3264.500 ;
        RECT 1890.900 3264.180 1891.220 3264.500 ;
        RECT 1917.580 3264.180 1917.900 3264.500 ;
        RECT 2542.260 3264.180 2542.580 3264.500 ;
        RECT 2567.100 3264.180 2567.420 3264.500 ;
        RECT 1317.855 3258.060 1318.175 3258.380 ;
        RECT 302.980 2894.940 303.300 2895.260 ;
        RECT 944.220 2894.940 944.540 2895.260 ;
        RECT 1351.780 2935.740 1352.100 2936.060 ;
        RECT 1412.500 2894.940 1412.820 2895.260 ;
        RECT 1551.420 2894.940 1551.740 2895.260 ;
        RECT 1946.100 2935.740 1946.420 2936.060 ;
        RECT 2187.140 2894.940 2187.460 2895.260 ;
        RECT 2587.340 2935.740 2587.660 2936.060 ;
        RECT 1055.540 2799.740 1055.860 2800.060 ;
        RECT 1794.860 2799.060 1795.180 2799.380 ;
        RECT 1795.220 2797.700 1795.540 2798.020 ;
        RECT 1052.780 2795.660 1053.100 2795.980 ;
        RECT 1732.660 2795.660 1732.980 2795.980 ;
        RECT 337.020 2794.300 337.340 2794.620 ;
        RECT 342.540 2794.300 342.860 2794.620 ;
        RECT 350.820 2794.300 351.140 2794.620 ;
        RECT 358.180 2794.300 358.500 2794.620 ;
        RECT 361.860 2794.300 362.180 2794.620 ;
        RECT 364.620 2794.300 364.940 2794.620 ;
        RECT 368.300 2794.300 368.620 2794.620 ;
        RECT 371.060 2794.300 371.380 2794.620 ;
        RECT 374.740 2794.300 375.060 2794.620 ;
        RECT 378.420 2794.300 378.740 2794.620 ;
        RECT 379.340 2794.300 379.660 2794.620 ;
        RECT 383.940 2794.300 384.260 2794.620 ;
        RECT 386.700 2794.300 387.020 2794.620 ;
        RECT 390.380 2794.300 390.700 2794.620 ;
        RECT 392.220 2794.300 392.540 2794.620 ;
        RECT 395.900 2794.300 396.220 2794.620 ;
        RECT 399.580 2794.300 399.900 2794.620 ;
        RECT 403.260 2794.300 403.580 2794.620 ;
        RECT 406.020 2794.300 406.340 2794.620 ;
        RECT 409.700 2794.300 410.020 2794.620 ;
        RECT 413.380 2794.300 413.700 2794.620 ;
        RECT 414.300 2794.300 414.620 2794.620 ;
        RECT 417.980 2794.300 418.300 2794.620 ;
        RECT 420.740 2794.300 421.060 2794.620 ;
        RECT 425.340 2794.300 425.660 2794.620 ;
        RECT 431.780 2794.300 432.100 2794.620 ;
        RECT 433.620 2794.300 433.940 2794.620 ;
        RECT 439.140 2794.300 439.460 2794.620 ;
        RECT 440.980 2794.300 441.300 2794.620 ;
        RECT 444.660 2794.300 444.980 2794.620 ;
        RECT 445.580 2794.300 445.900 2794.620 ;
        RECT 450.180 2794.300 450.500 2794.620 ;
        RECT 454.780 2794.300 455.100 2794.620 ;
        RECT 460.300 2794.300 460.620 2794.620 ;
        RECT 466.740 2794.300 467.060 2794.620 ;
        RECT 468.580 2794.300 468.900 2794.620 ;
        RECT 475.020 2794.300 475.340 2794.620 ;
        RECT 478.700 2794.300 479.020 2794.620 ;
        RECT 482.380 2794.300 482.700 2794.620 ;
        RECT 485.140 2794.300 485.460 2794.620 ;
        RECT 488.820 2794.300 489.140 2794.620 ;
        RECT 491.580 2794.300 491.900 2794.620 ;
        RECT 495.260 2794.300 495.580 2794.620 ;
        RECT 500.780 2794.300 501.100 2794.620 ;
        RECT 507.220 2794.300 507.540 2794.620 ;
        RECT 513.660 2794.300 513.980 2794.620 ;
        RECT 516.420 2794.300 516.740 2794.620 ;
        RECT 523.780 2794.300 524.100 2794.620 ;
        RECT 526.540 2794.300 526.860 2794.620 ;
        RECT 530.220 2794.300 530.540 2794.620 ;
        RECT 535.740 2794.300 536.060 2794.620 ;
        RECT 538.500 2794.300 538.820 2794.620 ;
        RECT 542.180 2794.300 542.500 2794.620 ;
        RECT 547.700 2794.300 548.020 2794.620 ;
        RECT 981.020 2794.300 981.340 2794.620 ;
        RECT 1013.220 2794.300 1013.540 2794.620 ;
        RECT 1018.740 2794.300 1019.060 2794.620 ;
        RECT 1019.660 2794.300 1019.980 2794.620 ;
        RECT 1027.020 2794.300 1027.340 2794.620 ;
        RECT 1030.700 2794.300 1031.020 2794.620 ;
        RECT 1041.740 2794.300 1042.060 2794.620 ;
        RECT 1059.220 2794.300 1059.540 2794.620 ;
        RECT 1065.660 2794.300 1065.980 2794.620 ;
        RECT 1070.260 2794.300 1070.580 2794.620 ;
        RECT 1081.300 2794.300 1081.620 2794.620 ;
        RECT 1087.740 2794.300 1088.060 2794.620 ;
        RECT 1089.580 2794.300 1089.900 2794.620 ;
        RECT 1094.180 2794.300 1094.500 2794.620 ;
        RECT 1096.020 2794.300 1096.340 2794.620 ;
        RECT 1100.620 2794.300 1100.940 2794.620 ;
        RECT 1103.380 2794.300 1103.700 2794.620 ;
        RECT 1105.220 2794.300 1105.540 2794.620 ;
        RECT 1109.820 2794.300 1110.140 2794.620 ;
        RECT 1111.660 2794.300 1111.980 2794.620 ;
        RECT 1118.100 2794.300 1118.420 2794.620 ;
        RECT 1121.780 2794.300 1122.100 2794.620 ;
        RECT 1129.140 2794.300 1129.460 2794.620 ;
        RECT 1130.980 2794.300 1131.300 2794.620 ;
        RECT 1135.580 2794.300 1135.900 2794.620 ;
        RECT 1137.420 2794.300 1137.740 2794.620 ;
        RECT 1140.180 2794.300 1140.500 2794.620 ;
        RECT 1143.860 2794.300 1144.180 2794.620 ;
        RECT 1146.620 2794.300 1146.940 2794.620 ;
        RECT 1151.220 2794.300 1151.540 2794.620 ;
        RECT 1153.980 2794.300 1154.300 2794.620 ;
        RECT 1165.020 2794.300 1165.340 2794.620 ;
        RECT 1172.380 2794.300 1172.700 2794.620 ;
        RECT 1178.820 2794.300 1179.140 2794.620 ;
        RECT 1186.180 2794.300 1186.500 2794.620 ;
        RECT 1198.140 2794.300 1198.460 2794.620 ;
        RECT 1613.060 2794.300 1613.380 2794.620 ;
        RECT 1642.500 2794.300 1642.820 2794.620 ;
        RECT 1652.620 2794.300 1652.940 2794.620 ;
        RECT 1659.060 2794.300 1659.380 2794.620 ;
        RECT 1665.500 2794.300 1665.820 2794.620 ;
        RECT 1670.100 2794.300 1670.420 2794.620 ;
        RECT 1677.460 2794.300 1677.780 2794.620 ;
        RECT 1694.940 2794.300 1695.260 2794.620 ;
        RECT 1699.540 2794.300 1699.860 2794.620 ;
        RECT 1705.980 2794.300 1706.300 2794.620 ;
        RECT 1712.420 2794.300 1712.740 2794.620 ;
        RECT 1717.940 2794.300 1718.260 2794.620 ;
        RECT 1723.460 2794.300 1723.780 2794.620 ;
        RECT 1728.980 2794.300 1729.300 2794.620 ;
        RECT 1740.940 2794.300 1741.260 2794.620 ;
        RECT 1747.380 2794.300 1747.700 2794.620 ;
        RECT 1762.100 2794.300 1762.420 2794.620 ;
        RECT 2243.260 2794.300 2243.580 2794.620 ;
        RECT 2257.060 2794.300 2257.380 2794.620 ;
        RECT 2264.420 2794.300 2264.740 2794.620 ;
        RECT 2268.100 2794.300 2268.420 2794.620 ;
        RECT 2276.380 2794.300 2276.700 2794.620 ;
        RECT 2282.820 2794.300 2283.140 2794.620 ;
        RECT 2287.420 2794.300 2287.740 2794.620 ;
        RECT 2293.860 2794.300 2294.180 2794.620 ;
        RECT 2300.300 2794.300 2300.620 2794.620 ;
        RECT 2304.900 2794.300 2305.220 2794.620 ;
        RECT 2308.580 2794.300 2308.900 2794.620 ;
        RECT 2316.860 2794.300 2317.180 2794.620 ;
        RECT 2322.380 2794.300 2322.700 2794.620 ;
        RECT 2328.820 2794.300 2329.140 2794.620 ;
        RECT 2334.340 2794.300 2334.660 2794.620 ;
        RECT 2339.860 2794.300 2340.180 2794.620 ;
        RECT 2343.540 2794.300 2343.860 2794.620 ;
        RECT 2351.820 2794.300 2352.140 2794.620 ;
        RECT 2357.340 2794.300 2357.660 2794.620 ;
        RECT 2363.780 2794.300 2364.100 2794.620 ;
        RECT 2370.220 2794.300 2370.540 2794.620 ;
        RECT 2373.900 2794.300 2374.220 2794.620 ;
        RECT 2385.860 2794.300 2386.180 2794.620 ;
        RECT 2391.380 2794.300 2391.700 2794.620 ;
        RECT 2395.060 2794.300 2395.380 2794.620 ;
        RECT 2420.820 2794.300 2421.140 2794.620 ;
        RECT 2430.020 2794.300 2430.340 2794.620 ;
        RECT 396.820 2793.620 397.140 2793.940 ;
        RECT 427.180 2793.620 427.500 2793.940 ;
        RECT 430.860 2793.620 431.180 2793.940 ;
        RECT 455.700 2793.620 456.020 2793.940 ;
        RECT 462.140 2793.620 462.460 2793.940 ;
        RECT 465.820 2793.620 466.140 2793.940 ;
        RECT 474.100 2793.620 474.420 2793.940 ;
        RECT 498.020 2793.620 498.340 2793.940 ;
        RECT 509.060 2793.620 509.380 2793.940 ;
        RECT 509.980 2793.620 510.300 2793.940 ;
        RECT 531.140 2793.620 531.460 2793.940 ;
        RECT 987.460 2793.620 987.780 2793.940 ;
        RECT 1001.260 2793.620 1001.580 2793.940 ;
        RECT 1076.700 2793.620 1077.020 2793.940 ;
        RECT 1083.140 2793.620 1083.460 2793.940 ;
        RECT 1086.820 2793.620 1087.140 2793.940 ;
        RECT 1122.700 2793.620 1123.020 2793.940 ;
        RECT 1128.220 2793.620 1128.540 2793.940 ;
        RECT 1163.180 2793.620 1163.500 2793.940 ;
        RECT 1173.300 2793.620 1173.620 2793.940 ;
        RECT 1180.660 2793.620 1180.980 2793.940 ;
        RECT 1187.100 2793.620 1187.420 2793.940 ;
        RECT 1688.500 2793.620 1688.820 2793.940 ;
        RECT 1767.620 2793.620 1767.940 2793.940 ;
        RECT 1780.500 2793.620 1780.820 2793.940 ;
        RECT 2269.020 2793.620 2269.340 2793.940 ;
        RECT 2273.620 2793.620 2273.940 2793.940 ;
        RECT 2280.060 2793.620 2280.380 2793.940 ;
        RECT 2284.660 2793.620 2284.980 2793.940 ;
        RECT 2297.540 2793.620 2297.860 2793.940 ;
        RECT 2303.980 2793.620 2304.300 2793.940 ;
        RECT 2310.420 2793.620 2310.740 2793.940 ;
        RECT 2315.020 2793.620 2315.340 2793.940 ;
        RECT 2321.460 2793.620 2321.780 2793.940 ;
        RECT 2326.060 2793.620 2326.380 2793.940 ;
        RECT 2332.500 2793.620 2332.820 2793.940 ;
        RECT 2345.380 2793.620 2345.700 2793.940 ;
        RECT 2348.140 2793.620 2348.460 2793.940 ;
        RECT 2356.420 2793.620 2356.740 2793.940 ;
        RECT 2361.020 2793.620 2361.340 2793.940 ;
        RECT 2367.460 2793.620 2367.780 2793.940 ;
        RECT 2377.580 2793.620 2377.900 2793.940 ;
        RECT 2403.340 2793.620 2403.660 2793.940 ;
        RECT 2423.580 2793.620 2423.900 2793.940 ;
        RECT 2436.460 2793.620 2436.780 2793.940 ;
        RECT 501.700 2792.940 502.020 2793.260 ;
        RECT 520.100 2792.940 520.420 2793.260 ;
        RECT 543.100 2792.940 543.420 2793.260 ;
        RECT 1012.300 2792.940 1012.620 2793.260 ;
        RECT 1024.260 2792.940 1024.580 2793.260 ;
        RECT 1048.180 2792.940 1048.500 2793.260 ;
        RECT 1167.780 2792.940 1168.100 2793.260 ;
        RECT 1636.980 2792.940 1637.300 2793.260 ;
        RECT 1681.140 2792.940 1681.460 2793.260 ;
        RECT 1787.860 2792.940 1788.180 2793.260 ;
        RECT 2263.500 2792.940 2263.820 2793.260 ;
        RECT 2292.020 2792.940 2292.340 2793.260 ;
        RECT 2338.940 2792.940 2339.260 2793.260 ;
        RECT 2374.820 2792.940 2375.140 2793.260 ;
        RECT 2404.260 2792.940 2404.580 2793.260 ;
        RECT 2407.940 2792.940 2408.260 2793.260 ;
        RECT 2415.300 2792.940 2415.620 2793.260 ;
        RECT 2442.900 2792.940 2443.220 2793.260 ;
        RECT 348.980 2792.260 349.300 2792.580 ;
        RECT 1116.260 2792.260 1116.580 2792.580 ;
        RECT 1153.060 2792.260 1153.380 2792.580 ;
        RECT 1637.900 2792.260 1638.220 2792.580 ;
        RECT 1752.900 2792.260 1753.220 2792.580 ;
        RECT 2418.060 2792.260 2418.380 2792.580 ;
        RECT 1159.500 2791.580 1159.820 2791.900 ;
        RECT 1193.540 2791.580 1193.860 2791.900 ;
        RECT 1587.300 2791.580 1587.620 2791.900 ;
        RECT 1602.940 2791.580 1603.260 2791.900 ;
        RECT 1759.340 2791.580 1759.660 2791.900 ;
        RECT 1774.060 2791.580 1774.380 2791.900 ;
        RECT 1794.300 2791.580 1794.620 2791.900 ;
        RECT 2392.300 2791.580 2392.620 2791.900 ;
        RECT 2433.700 2791.580 2434.020 2791.900 ;
        RECT 2439.220 2791.580 2439.540 2791.900 ;
        RECT 993.900 2790.900 994.220 2791.220 ;
        RECT 1164.100 2790.900 1164.420 2791.220 ;
        RECT 1417.100 2790.900 1417.420 2791.220 ;
        RECT 2249.700 2790.900 2250.020 2791.220 ;
        RECT 1191.700 2790.220 1192.020 2790.540 ;
        RECT 1644.340 2790.220 1644.660 2790.540 ;
        RECT 2386.780 2790.220 2387.100 2790.540 ;
        RECT 2398.740 2790.220 2399.060 2790.540 ;
        RECT 2410.700 2790.900 2411.020 2791.220 ;
        RECT 2445.660 2790.220 2445.980 2790.540 ;
        RECT 1648.020 2789.540 1648.340 2789.860 ;
        RECT 2381.260 2789.540 2381.580 2789.860 ;
        RECT 2236.820 2788.860 2237.140 2789.180 ;
        RECT 2417.140 2788.860 2417.460 2789.180 ;
        RECT 1007.700 2788.180 1008.020 2788.500 ;
        RECT 1035.300 2788.180 1035.620 2788.500 ;
        RECT 1051.860 2788.180 1052.180 2788.500 ;
        RECT 1618.580 2788.180 1618.900 2788.500 ;
        RECT 1624.100 2788.180 1624.420 2788.500 ;
        RECT 1631.460 2788.180 1631.780 2788.500 ;
        RECT 1655.380 2788.180 1655.700 2788.500 ;
        RECT 1689.420 2788.180 1689.740 2788.500 ;
        RECT 1724.380 2788.180 1724.700 2788.500 ;
        RECT 1765.780 2788.180 1766.100 2788.500 ;
        RECT 2428.180 2788.180 2428.500 2788.500 ;
        RECT 1034.380 2787.500 1034.700 2787.820 ;
        RECT 1039.900 2787.500 1040.220 2787.820 ;
        RECT 1046.340 2787.500 1046.660 2787.820 ;
        RECT 1061.980 2787.500 1062.300 2787.820 ;
        RECT 1067.500 2787.500 1067.820 2787.820 ;
        RECT 1073.940 2787.500 1074.260 2787.820 ;
        RECT 1580.860 2787.500 1581.180 2787.820 ;
        RECT 1594.660 2787.500 1594.980 2787.820 ;
        RECT 1604.780 2787.500 1605.100 2787.820 ;
        RECT 1613.980 2787.500 1614.300 2787.820 ;
        RECT 1620.420 2787.500 1620.740 2787.820 ;
        RECT 1626.860 2787.500 1627.180 2787.820 ;
        RECT 1630.540 2787.500 1630.860 2787.820 ;
        RECT 1648.940 2787.500 1649.260 2787.820 ;
        RECT 1660.900 2787.500 1661.220 2787.820 ;
        RECT 1666.420 2787.500 1666.740 2787.820 ;
        RECT 1672.860 2787.500 1673.180 2787.820 ;
        RECT 1678.380 2787.500 1678.700 2787.820 ;
        RECT 1683.900 2787.500 1684.220 2787.820 ;
        RECT 1695.860 2787.500 1696.180 2787.820 ;
        RECT 1702.300 2787.500 1702.620 2787.820 ;
        RECT 1708.740 2787.500 1709.060 2787.820 ;
        RECT 1713.340 2787.500 1713.660 2787.820 ;
        RECT 1719.780 2787.500 1720.100 2787.820 ;
        RECT 1730.820 2787.500 1731.140 2787.820 ;
        RECT 1737.260 2787.500 1737.580 2787.820 ;
        RECT 1743.700 2787.500 1744.020 2787.820 ;
        RECT 1748.300 2787.500 1748.620 2787.820 ;
        RECT 1754.740 2787.500 1755.060 2787.820 ;
        RECT 1760.260 2787.500 1760.580 2787.820 ;
        RECT 1772.220 2787.500 1772.540 2787.820 ;
        RECT 1777.740 2787.500 1778.060 2787.820 ;
        RECT 1783.260 2787.500 1783.580 2787.820 ;
        RECT 1789.700 2787.500 1790.020 2787.820 ;
        RECT 1795.220 2787.500 1795.540 2787.820 ;
        RECT 2231.300 2787.500 2231.620 2787.820 ;
        RECT 1410.660 2087.100 1410.980 2087.420 ;
        RECT 1410.660 1657.340 1410.980 1657.660 ;
        RECT 1417.100 1627.420 1417.420 1627.740 ;
      LAYER met4 ;
        RECT 646.135 3264.175 646.465 3264.505 ;
        RECT 668.215 3264.175 668.545 3264.505 ;
        RECT 1292.895 3264.175 1293.225 3264.505 ;
        RECT 1890.895 3264.175 1891.225 3264.505 ;
        RECT 1917.575 3264.175 1917.905 3264.505 ;
        RECT 2542.255 3264.175 2542.585 3264.505 ;
        RECT 2567.095 3264.175 2567.425 3264.505 ;
        RECT 394.025 3251.635 394.325 3256.235 ;
        RECT 400.265 3251.635 400.565 3256.235 ;
        RECT 406.505 3251.635 406.805 3256.235 ;
        RECT 412.745 3251.635 413.045 3256.235 ;
        RECT 418.985 3251.635 419.285 3256.235 ;
        RECT 425.225 3251.635 425.525 3256.235 ;
        RECT 431.465 3251.635 431.765 3256.235 ;
        RECT 437.705 3251.635 438.005 3256.235 ;
        RECT 443.945 3251.635 444.245 3256.235 ;
        RECT 450.185 3251.635 450.485 3256.235 ;
        RECT 456.425 3251.635 456.725 3256.235 ;
        RECT 462.665 3251.635 462.965 3256.235 ;
        RECT 468.905 3251.635 469.205 3256.235 ;
        RECT 475.145 3251.635 475.445 3256.235 ;
        RECT 481.385 3251.635 481.685 3256.235 ;
        RECT 487.625 3251.635 487.925 3256.235 ;
        RECT 493.865 3251.635 494.165 3256.235 ;
        RECT 500.105 3251.635 500.405 3256.235 ;
        RECT 506.345 3251.635 506.645 3256.235 ;
        RECT 512.585 3251.635 512.885 3256.235 ;
        RECT 518.825 3251.635 519.125 3256.235 ;
        RECT 525.065 3251.635 525.365 3256.235 ;
        RECT 531.305 3251.635 531.605 3256.235 ;
        RECT 537.545 3251.635 537.845 3256.235 ;
        RECT 543.785 3251.635 544.085 3256.235 ;
        RECT 550.025 3251.635 550.325 3256.235 ;
        RECT 556.265 3251.635 556.565 3256.235 ;
        RECT 562.505 3251.635 562.805 3256.235 ;
        RECT 568.745 3251.635 569.045 3256.235 ;
        RECT 574.985 3251.635 575.285 3256.235 ;
        RECT 581.225 3251.635 581.525 3256.235 ;
        RECT 587.465 3251.635 587.765 3256.235 ;
        RECT 642.890 3255.650 643.190 3256.235 ;
        RECT 646.150 3255.650 646.450 3264.175 ;
        RECT 668.230 3259.050 668.530 3264.175 ;
        RECT 642.890 3255.350 646.450 3255.650 ;
        RECT 667.865 3258.750 668.530 3259.050 ;
        RECT 642.890 3251.635 643.190 3255.350 ;
        RECT 667.865 3251.635 668.165 3258.750 ;
        RECT 1292.910 3256.235 1293.210 3264.175 ;
        RECT 1317.850 3258.055 1318.180 3258.385 ;
        RECT 1044.025 3251.635 1044.325 3256.235 ;
        RECT 1050.265 3251.635 1050.565 3256.235 ;
        RECT 1056.505 3251.635 1056.805 3256.235 ;
        RECT 1062.745 3251.635 1063.045 3256.235 ;
        RECT 1068.985 3251.635 1069.285 3256.235 ;
        RECT 1075.225 3251.635 1075.525 3256.235 ;
        RECT 1081.465 3251.635 1081.765 3256.235 ;
        RECT 1087.705 3251.635 1088.005 3256.235 ;
        RECT 1093.945 3251.635 1094.245 3256.235 ;
        RECT 1100.185 3251.635 1100.485 3256.235 ;
        RECT 1106.425 3251.635 1106.725 3256.235 ;
        RECT 1112.665 3251.635 1112.965 3256.235 ;
        RECT 1118.905 3251.635 1119.205 3256.235 ;
        RECT 1125.145 3251.635 1125.445 3256.235 ;
        RECT 1131.385 3251.635 1131.685 3256.235 ;
        RECT 1137.625 3251.635 1137.925 3256.235 ;
        RECT 1143.865 3251.635 1144.165 3256.235 ;
        RECT 1150.105 3251.635 1150.405 3256.235 ;
        RECT 1156.345 3251.635 1156.645 3256.235 ;
        RECT 1162.585 3251.635 1162.885 3256.235 ;
        RECT 1168.825 3251.635 1169.125 3256.235 ;
        RECT 1175.065 3251.635 1175.365 3256.235 ;
        RECT 1181.305 3251.635 1181.605 3256.235 ;
        RECT 1187.545 3251.635 1187.845 3256.235 ;
        RECT 1193.785 3251.635 1194.085 3256.235 ;
        RECT 1200.025 3251.635 1200.325 3256.235 ;
        RECT 1206.265 3251.635 1206.565 3256.235 ;
        RECT 1212.505 3251.635 1212.805 3256.235 ;
        RECT 1218.745 3251.635 1219.045 3256.235 ;
        RECT 1224.985 3251.635 1225.285 3256.235 ;
        RECT 1231.225 3251.635 1231.525 3256.235 ;
        RECT 1237.465 3251.635 1237.765 3256.235 ;
        RECT 1292.890 3255.350 1293.210 3256.235 ;
        RECT 1292.890 3251.635 1293.190 3255.350 ;
        RECT 1317.865 3251.635 1318.165 3258.055 ;
        RECT 1644.025 3251.635 1644.325 3256.235 ;
        RECT 1650.265 3251.635 1650.565 3256.235 ;
        RECT 1656.505 3251.635 1656.805 3256.235 ;
        RECT 1662.745 3251.635 1663.045 3256.235 ;
        RECT 1668.985 3251.635 1669.285 3256.235 ;
        RECT 1675.225 3251.635 1675.525 3256.235 ;
        RECT 1681.465 3251.635 1681.765 3256.235 ;
        RECT 1687.705 3251.635 1688.005 3256.235 ;
        RECT 1693.945 3251.635 1694.245 3256.235 ;
        RECT 1700.185 3251.635 1700.485 3256.235 ;
        RECT 1706.425 3251.635 1706.725 3256.235 ;
        RECT 1712.665 3251.635 1712.965 3256.235 ;
        RECT 1718.905 3251.635 1719.205 3256.235 ;
        RECT 1725.145 3251.635 1725.445 3256.235 ;
        RECT 1731.385 3251.635 1731.685 3256.235 ;
        RECT 1737.625 3251.635 1737.925 3256.235 ;
        RECT 1743.865 3251.635 1744.165 3256.235 ;
        RECT 1750.105 3251.635 1750.405 3256.235 ;
        RECT 1756.345 3251.635 1756.645 3256.235 ;
        RECT 1762.585 3251.635 1762.885 3256.235 ;
        RECT 1768.825 3251.635 1769.125 3256.235 ;
        RECT 1775.065 3251.635 1775.365 3256.235 ;
        RECT 1781.305 3251.635 1781.605 3256.235 ;
        RECT 1787.545 3251.635 1787.845 3256.235 ;
        RECT 1793.785 3251.635 1794.085 3256.235 ;
        RECT 1800.025 3251.635 1800.325 3256.235 ;
        RECT 1806.265 3251.635 1806.565 3256.235 ;
        RECT 1812.505 3251.635 1812.805 3256.235 ;
        RECT 1818.745 3251.635 1819.045 3256.235 ;
        RECT 1824.985 3251.635 1825.285 3256.235 ;
        RECT 1831.225 3251.635 1831.525 3256.235 ;
        RECT 1837.465 3251.635 1837.765 3256.235 ;
        RECT 1890.910 3255.650 1891.210 3264.175 ;
        RECT 1917.590 3256.235 1917.890 3264.175 ;
        RECT 1892.890 3255.650 1893.190 3256.235 ;
        RECT 1890.910 3255.350 1893.190 3255.650 ;
        RECT 1917.590 3255.350 1918.165 3256.235 ;
        RECT 1892.890 3251.635 1893.190 3255.350 ;
        RECT 1917.865 3251.635 1918.165 3255.350 ;
        RECT 2294.025 3251.635 2294.325 3256.235 ;
        RECT 2300.265 3251.635 2300.565 3256.235 ;
        RECT 2306.505 3251.635 2306.805 3256.235 ;
        RECT 2312.745 3251.635 2313.045 3256.235 ;
        RECT 2318.985 3251.635 2319.285 3256.235 ;
        RECT 2325.225 3251.635 2325.525 3256.235 ;
        RECT 2331.465 3251.635 2331.765 3256.235 ;
        RECT 2337.705 3251.635 2338.005 3256.235 ;
        RECT 2343.945 3251.635 2344.245 3256.235 ;
        RECT 2350.185 3251.635 2350.485 3256.235 ;
        RECT 2356.425 3251.635 2356.725 3256.235 ;
        RECT 2362.665 3251.635 2362.965 3256.235 ;
        RECT 2368.905 3251.635 2369.205 3256.235 ;
        RECT 2375.145 3251.635 2375.445 3256.235 ;
        RECT 2381.385 3251.635 2381.685 3256.235 ;
        RECT 2387.625 3251.635 2387.925 3256.235 ;
        RECT 2393.865 3251.635 2394.165 3256.235 ;
        RECT 2400.105 3251.635 2400.405 3256.235 ;
        RECT 2406.345 3251.635 2406.645 3256.235 ;
        RECT 2412.585 3251.635 2412.885 3256.235 ;
        RECT 2418.825 3251.635 2419.125 3256.235 ;
        RECT 2425.065 3251.635 2425.365 3256.235 ;
        RECT 2431.305 3251.635 2431.605 3256.235 ;
        RECT 2437.545 3251.635 2437.845 3256.235 ;
        RECT 2443.785 3251.635 2444.085 3256.235 ;
        RECT 2450.025 3251.635 2450.325 3256.235 ;
        RECT 2456.265 3251.635 2456.565 3256.235 ;
        RECT 2462.505 3251.635 2462.805 3256.235 ;
        RECT 2468.745 3251.635 2469.045 3256.235 ;
        RECT 2474.985 3251.635 2475.285 3256.235 ;
        RECT 2481.225 3251.635 2481.525 3256.235 ;
        RECT 2487.465 3251.635 2487.765 3256.235 ;
        RECT 2542.270 3255.650 2542.570 3264.175 ;
        RECT 2542.890 3255.650 2543.190 3256.235 ;
        RECT 2542.270 3255.350 2543.190 3255.650 ;
        RECT 2567.110 3255.650 2567.410 3264.175 ;
        RECT 2567.865 3255.650 2568.165 3256.235 ;
        RECT 2567.110 3255.350 2568.165 3255.650 ;
        RECT 2542.890 3251.635 2543.190 3255.350 ;
        RECT 2567.865 3251.635 2568.165 3255.350 ;
        RECT 302.550 2894.510 303.730 2895.690 ;
      LAYER met4 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met4 ;
        RECT 943.790 2894.510 944.970 2895.690 ;
      LAYER met4 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met4 ;
        RECT 1351.350 2935.310 1352.530 2936.490 ;
        RECT 1412.070 2894.510 1413.250 2895.690 ;
        RECT 1550.990 2894.510 1552.170 2895.690 ;
      LAYER met4 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met4 ;
        RECT 1945.670 2935.310 1946.850 2936.490 ;
        RECT 2186.710 2894.510 2187.890 2895.690 ;
      LAYER met4 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met4 ;
        RECT 2586.910 2935.310 2588.090 2936.490 ;
        RECT 334.010 2801.750 334.310 2804.600 ;
        RECT 339.850 2801.750 340.150 2804.600 ;
        RECT 345.690 2801.750 345.990 2804.600 ;
        RECT 351.530 2801.750 351.830 2804.600 ;
        RECT 334.010 2801.450 337.330 2801.750 ;
        RECT 334.010 2800.000 334.310 2801.450 ;
        RECT 337.030 2794.625 337.330 2801.450 ;
        RECT 339.850 2801.450 342.850 2801.750 ;
        RECT 339.850 2800.000 340.150 2801.450 ;
        RECT 342.550 2794.625 342.850 2801.450 ;
        RECT 345.690 2801.450 349.290 2801.750 ;
        RECT 345.690 2800.000 345.990 2801.450 ;
        RECT 337.015 2794.295 337.345 2794.625 ;
        RECT 342.535 2794.295 342.865 2794.625 ;
        RECT 348.990 2792.585 349.290 2801.450 ;
        RECT 350.830 2801.450 351.830 2801.750 ;
        RECT 350.830 2794.625 351.130 2801.450 ;
        RECT 351.530 2800.000 351.830 2801.450 ;
        RECT 357.370 2801.750 357.670 2804.600 ;
        RECT 363.210 2802.450 363.510 2804.600 ;
        RECT 361.870 2802.150 363.510 2802.450 ;
        RECT 357.370 2801.450 358.490 2801.750 ;
        RECT 357.370 2800.000 357.670 2801.450 ;
        RECT 358.190 2794.625 358.490 2801.450 ;
        RECT 361.870 2794.625 362.170 2802.150 ;
        RECT 363.210 2800.000 363.510 2802.150 ;
        RECT 363.830 2801.750 364.130 2804.600 ;
        RECT 369.050 2801.750 369.350 2804.600 ;
        RECT 363.830 2801.450 364.930 2801.750 ;
        RECT 363.830 2800.000 364.130 2801.450 ;
        RECT 364.630 2794.625 364.930 2801.450 ;
        RECT 368.310 2801.450 369.350 2801.750 ;
        RECT 368.310 2794.625 368.610 2801.450 ;
        RECT 369.050 2800.000 369.350 2801.450 ;
        RECT 369.670 2801.750 369.970 2804.600 ;
        RECT 374.890 2801.750 375.190 2804.600 ;
        RECT 369.670 2801.450 371.370 2801.750 ;
        RECT 369.670 2800.000 369.970 2801.450 ;
        RECT 371.070 2794.625 371.370 2801.450 ;
        RECT 374.750 2800.000 375.190 2801.750 ;
        RECT 375.510 2801.750 375.810 2804.600 ;
        RECT 380.730 2802.450 381.030 2804.600 ;
        RECT 379.350 2802.150 381.030 2802.450 ;
        RECT 375.510 2801.450 378.730 2801.750 ;
        RECT 375.510 2800.000 375.810 2801.450 ;
        RECT 374.750 2794.625 375.050 2800.000 ;
        RECT 378.430 2794.625 378.730 2801.450 ;
        RECT 379.350 2794.625 379.650 2802.150 ;
        RECT 380.730 2800.000 381.030 2802.150 ;
        RECT 381.350 2801.750 381.650 2804.600 ;
        RECT 381.350 2801.450 384.250 2801.750 ;
        RECT 381.350 2800.000 381.650 2801.450 ;
        RECT 383.950 2794.625 384.250 2801.450 ;
        RECT 386.570 2796.650 386.870 2804.600 ;
        RECT 387.190 2801.750 387.490 2804.600 ;
        RECT 392.410 2801.750 392.710 2804.600 ;
        RECT 387.190 2801.450 390.690 2801.750 ;
        RECT 387.190 2800.000 387.490 2801.450 ;
        RECT 386.570 2796.350 387.010 2796.650 ;
        RECT 386.710 2794.625 387.010 2796.350 ;
        RECT 390.390 2794.625 390.690 2801.450 ;
        RECT 392.230 2800.000 392.710 2801.750 ;
        RECT 393.030 2801.750 393.330 2804.600 ;
        RECT 398.250 2802.450 398.550 2804.600 ;
        RECT 396.830 2802.150 398.550 2802.450 ;
        RECT 393.030 2801.450 396.210 2801.750 ;
        RECT 393.030 2800.000 393.330 2801.450 ;
        RECT 392.230 2794.625 392.530 2800.000 ;
        RECT 395.910 2794.625 396.210 2801.450 ;
        RECT 350.815 2794.295 351.145 2794.625 ;
        RECT 358.175 2794.295 358.505 2794.625 ;
        RECT 361.855 2794.295 362.185 2794.625 ;
        RECT 364.615 2794.295 364.945 2794.625 ;
        RECT 368.295 2794.295 368.625 2794.625 ;
        RECT 371.055 2794.295 371.385 2794.625 ;
        RECT 374.735 2794.295 375.065 2794.625 ;
        RECT 378.415 2794.295 378.745 2794.625 ;
        RECT 379.335 2794.295 379.665 2794.625 ;
        RECT 383.935 2794.295 384.265 2794.625 ;
        RECT 386.695 2794.295 387.025 2794.625 ;
        RECT 390.375 2794.295 390.705 2794.625 ;
        RECT 392.215 2794.295 392.545 2794.625 ;
        RECT 395.895 2794.295 396.225 2794.625 ;
        RECT 396.830 2793.945 397.130 2802.150 ;
        RECT 398.250 2800.000 398.550 2802.150 ;
        RECT 398.870 2801.750 399.170 2804.600 ;
        RECT 404.090 2801.750 404.390 2804.600 ;
        RECT 398.870 2801.450 399.890 2801.750 ;
        RECT 398.870 2800.000 399.170 2801.450 ;
        RECT 399.590 2794.625 399.890 2801.450 ;
        RECT 403.270 2801.450 404.390 2801.750 ;
        RECT 403.270 2794.625 403.570 2801.450 ;
        RECT 404.090 2800.000 404.390 2801.450 ;
        RECT 404.710 2801.750 405.010 2804.600 ;
        RECT 409.930 2801.750 410.230 2804.600 ;
        RECT 404.710 2801.450 406.330 2801.750 ;
        RECT 404.710 2800.000 405.010 2801.450 ;
        RECT 406.030 2794.625 406.330 2801.450 ;
        RECT 409.710 2800.000 410.230 2801.750 ;
        RECT 410.550 2801.750 410.850 2804.600 ;
        RECT 415.770 2802.450 416.070 2804.600 ;
        RECT 414.310 2802.150 416.070 2802.450 ;
        RECT 410.550 2801.450 413.690 2801.750 ;
        RECT 410.550 2800.000 410.850 2801.450 ;
        RECT 409.710 2794.625 410.010 2800.000 ;
        RECT 413.390 2794.625 413.690 2801.450 ;
        RECT 414.310 2794.625 414.610 2802.150 ;
        RECT 415.770 2800.000 416.070 2802.150 ;
        RECT 416.390 2801.750 416.690 2804.600 ;
        RECT 421.610 2801.750 421.910 2804.600 ;
        RECT 416.390 2801.450 418.290 2801.750 ;
        RECT 416.390 2800.000 416.690 2801.450 ;
        RECT 417.990 2794.625 418.290 2801.450 ;
        RECT 420.750 2801.450 421.910 2801.750 ;
        RECT 420.750 2794.625 421.050 2801.450 ;
        RECT 421.610 2800.000 421.910 2801.450 ;
        RECT 422.230 2801.750 422.530 2804.600 ;
        RECT 427.450 2801.750 427.750 2804.600 ;
        RECT 422.230 2801.450 425.650 2801.750 ;
        RECT 422.230 2800.000 422.530 2801.450 ;
        RECT 425.350 2794.625 425.650 2801.450 ;
        RECT 427.190 2800.000 427.750 2801.750 ;
        RECT 428.070 2801.750 428.370 2804.600 ;
        RECT 433.290 2802.450 433.590 2804.600 ;
        RECT 431.790 2802.150 433.590 2802.450 ;
        RECT 428.070 2801.450 431.170 2801.750 ;
        RECT 428.070 2800.000 428.370 2801.450 ;
        RECT 399.575 2794.295 399.905 2794.625 ;
        RECT 403.255 2794.295 403.585 2794.625 ;
        RECT 406.015 2794.295 406.345 2794.625 ;
        RECT 409.695 2794.295 410.025 2794.625 ;
        RECT 413.375 2794.295 413.705 2794.625 ;
        RECT 414.295 2794.295 414.625 2794.625 ;
        RECT 417.975 2794.295 418.305 2794.625 ;
        RECT 420.735 2794.295 421.065 2794.625 ;
        RECT 425.335 2794.295 425.665 2794.625 ;
        RECT 427.190 2793.945 427.490 2800.000 ;
        RECT 430.870 2793.945 431.170 2801.450 ;
        RECT 431.790 2794.625 432.090 2802.150 ;
        RECT 433.290 2800.000 433.590 2802.150 ;
        RECT 433.910 2796.650 434.210 2804.600 ;
        RECT 439.130 2800.050 439.430 2804.600 ;
        RECT 439.750 2801.750 440.050 2804.600 ;
        RECT 444.970 2801.750 445.270 2804.600 ;
        RECT 439.750 2801.450 441.290 2801.750 ;
        RECT 439.130 2799.750 439.450 2800.050 ;
        RECT 439.750 2800.000 440.050 2801.450 ;
        RECT 433.630 2796.350 434.210 2796.650 ;
        RECT 433.630 2794.625 433.930 2796.350 ;
        RECT 439.150 2794.625 439.450 2799.750 ;
        RECT 440.990 2794.625 441.290 2801.450 ;
        RECT 444.670 2800.000 445.270 2801.750 ;
        RECT 444.670 2794.625 444.970 2800.000 ;
        RECT 445.590 2794.625 445.890 2804.600 ;
        RECT 450.810 2801.750 451.110 2804.600 ;
        RECT 450.190 2801.450 451.110 2801.750 ;
        RECT 450.190 2794.625 450.490 2801.450 ;
        RECT 450.810 2800.000 451.110 2801.450 ;
        RECT 451.430 2801.750 451.730 2804.600 ;
        RECT 456.650 2801.750 456.950 2804.600 ;
        RECT 451.430 2801.450 455.090 2801.750 ;
        RECT 451.430 2800.000 451.730 2801.450 ;
        RECT 454.790 2794.625 455.090 2801.450 ;
        RECT 455.710 2801.450 456.950 2801.750 ;
        RECT 431.775 2794.295 432.105 2794.625 ;
        RECT 433.615 2794.295 433.945 2794.625 ;
        RECT 439.135 2794.295 439.465 2794.625 ;
        RECT 440.975 2794.295 441.305 2794.625 ;
        RECT 444.655 2794.295 444.985 2794.625 ;
        RECT 445.575 2794.295 445.905 2794.625 ;
        RECT 450.175 2794.295 450.505 2794.625 ;
        RECT 454.775 2794.295 455.105 2794.625 ;
        RECT 455.710 2793.945 456.010 2801.450 ;
        RECT 456.650 2800.000 456.950 2801.450 ;
        RECT 457.270 2801.750 457.570 2804.600 ;
        RECT 457.270 2801.450 460.610 2801.750 ;
        RECT 457.270 2800.000 457.570 2801.450 ;
        RECT 460.310 2794.625 460.610 2801.450 ;
        RECT 462.490 2800.050 462.790 2804.600 ;
        RECT 462.150 2799.750 462.790 2800.050 ;
        RECT 463.110 2801.750 463.410 2804.600 ;
        RECT 468.330 2801.750 468.630 2804.600 ;
        RECT 463.110 2801.450 466.130 2801.750 ;
        RECT 463.110 2800.000 463.410 2801.450 ;
        RECT 460.295 2794.295 460.625 2794.625 ;
        RECT 462.150 2793.945 462.450 2799.750 ;
        RECT 465.830 2793.945 466.130 2801.450 ;
        RECT 466.750 2801.450 468.630 2801.750 ;
        RECT 466.750 2794.625 467.050 2801.450 ;
        RECT 468.330 2800.000 468.630 2801.450 ;
        RECT 468.950 2796.650 469.250 2804.600 ;
        RECT 474.170 2801.750 474.470 2804.600 ;
        RECT 468.590 2796.350 469.250 2796.650 ;
        RECT 474.110 2800.000 474.470 2801.750 ;
        RECT 474.790 2801.750 475.090 2804.600 ;
        RECT 480.010 2801.750 480.310 2804.600 ;
        RECT 474.790 2800.000 475.330 2801.750 ;
        RECT 468.590 2794.625 468.890 2796.350 ;
        RECT 466.735 2794.295 467.065 2794.625 ;
        RECT 468.575 2794.295 468.905 2794.625 ;
        RECT 474.110 2793.945 474.410 2800.000 ;
        RECT 475.030 2794.625 475.330 2800.000 ;
        RECT 478.710 2801.450 480.310 2801.750 ;
        RECT 478.710 2794.625 479.010 2801.450 ;
        RECT 480.010 2800.000 480.310 2801.450 ;
        RECT 480.630 2801.750 480.930 2804.600 ;
        RECT 485.850 2801.750 486.150 2804.600 ;
        RECT 480.630 2801.450 482.690 2801.750 ;
        RECT 480.630 2800.000 480.930 2801.450 ;
        RECT 482.390 2794.625 482.690 2801.450 ;
        RECT 485.150 2801.450 486.150 2801.750 ;
        RECT 485.150 2794.625 485.450 2801.450 ;
        RECT 485.850 2800.000 486.150 2801.450 ;
        RECT 486.470 2801.750 486.770 2804.600 ;
        RECT 491.690 2801.750 491.990 2804.600 ;
        RECT 486.470 2801.450 489.130 2801.750 ;
        RECT 486.470 2800.000 486.770 2801.450 ;
        RECT 488.830 2794.625 489.130 2801.450 ;
        RECT 491.590 2800.000 491.990 2801.750 ;
        RECT 492.310 2801.750 492.610 2804.600 ;
        RECT 492.310 2801.450 495.570 2801.750 ;
        RECT 492.310 2800.000 492.610 2801.450 ;
        RECT 491.590 2794.625 491.890 2800.000 ;
        RECT 495.270 2794.625 495.570 2801.450 ;
        RECT 497.530 2796.650 497.830 2804.600 ;
        RECT 498.150 2801.750 498.450 2804.600 ;
        RECT 503.370 2801.750 503.670 2804.600 ;
        RECT 498.150 2801.450 501.090 2801.750 ;
        RECT 498.150 2800.000 498.450 2801.450 ;
        RECT 497.530 2796.350 498.330 2796.650 ;
        RECT 475.015 2794.295 475.345 2794.625 ;
        RECT 478.695 2794.295 479.025 2794.625 ;
        RECT 482.375 2794.295 482.705 2794.625 ;
        RECT 485.135 2794.295 485.465 2794.625 ;
        RECT 488.815 2794.295 489.145 2794.625 ;
        RECT 491.575 2794.295 491.905 2794.625 ;
        RECT 495.255 2794.295 495.585 2794.625 ;
        RECT 498.030 2793.945 498.330 2796.350 ;
        RECT 500.790 2794.625 501.090 2801.450 ;
        RECT 501.710 2801.450 503.670 2801.750 ;
        RECT 500.775 2794.295 501.105 2794.625 ;
        RECT 396.815 2793.615 397.145 2793.945 ;
        RECT 427.175 2793.615 427.505 2793.945 ;
        RECT 430.855 2793.615 431.185 2793.945 ;
        RECT 455.695 2793.615 456.025 2793.945 ;
        RECT 462.135 2793.615 462.465 2793.945 ;
        RECT 465.815 2793.615 466.145 2793.945 ;
        RECT 474.095 2793.615 474.425 2793.945 ;
        RECT 498.015 2793.615 498.345 2793.945 ;
        RECT 501.710 2793.265 502.010 2801.450 ;
        RECT 503.370 2800.000 503.670 2801.450 ;
        RECT 503.990 2801.750 504.290 2804.600 ;
        RECT 509.210 2801.750 509.510 2804.600 ;
        RECT 503.990 2801.450 507.530 2801.750 ;
        RECT 503.990 2800.000 504.290 2801.450 ;
        RECT 507.230 2794.625 507.530 2801.450 ;
        RECT 509.070 2800.000 509.510 2801.750 ;
        RECT 509.830 2801.750 510.130 2804.600 ;
        RECT 515.050 2801.750 515.350 2804.600 ;
        RECT 509.830 2800.000 510.290 2801.750 ;
        RECT 507.215 2794.295 507.545 2794.625 ;
        RECT 509.070 2793.945 509.370 2800.000 ;
        RECT 509.990 2793.945 510.290 2800.000 ;
        RECT 513.670 2801.450 515.350 2801.750 ;
        RECT 513.670 2794.625 513.970 2801.450 ;
        RECT 515.050 2800.000 515.350 2801.450 ;
        RECT 515.670 2801.750 515.970 2804.600 ;
        RECT 520.890 2801.750 521.190 2804.600 ;
        RECT 515.670 2801.450 516.730 2801.750 ;
        RECT 515.670 2800.000 515.970 2801.450 ;
        RECT 516.430 2794.625 516.730 2801.450 ;
        RECT 520.110 2801.450 521.190 2801.750 ;
        RECT 513.655 2794.295 513.985 2794.625 ;
        RECT 516.415 2794.295 516.745 2794.625 ;
        RECT 509.055 2793.615 509.385 2793.945 ;
        RECT 509.975 2793.615 510.305 2793.945 ;
        RECT 520.110 2793.265 520.410 2801.450 ;
        RECT 520.890 2800.000 521.190 2801.450 ;
        RECT 521.510 2801.750 521.810 2804.600 ;
        RECT 526.730 2801.750 527.030 2804.600 ;
        RECT 521.510 2801.450 524.090 2801.750 ;
        RECT 521.510 2800.000 521.810 2801.450 ;
        RECT 523.790 2794.625 524.090 2801.450 ;
        RECT 526.550 2800.000 527.030 2801.750 ;
        RECT 527.350 2801.750 527.650 2804.600 ;
        RECT 532.570 2802.450 532.870 2804.600 ;
        RECT 531.150 2802.150 532.870 2802.450 ;
        RECT 527.350 2801.450 530.530 2801.750 ;
        RECT 527.350 2800.000 527.650 2801.450 ;
        RECT 526.550 2794.625 526.850 2800.000 ;
        RECT 530.230 2794.625 530.530 2801.450 ;
        RECT 523.775 2794.295 524.105 2794.625 ;
        RECT 526.535 2794.295 526.865 2794.625 ;
        RECT 530.215 2794.295 530.545 2794.625 ;
        RECT 531.150 2793.945 531.450 2802.150 ;
        RECT 532.570 2800.000 532.870 2802.150 ;
        RECT 533.190 2801.750 533.490 2804.600 ;
        RECT 533.190 2801.450 536.050 2801.750 ;
        RECT 533.190 2800.000 533.490 2801.450 ;
        RECT 535.750 2794.625 536.050 2801.450 ;
        RECT 538.410 2796.650 538.710 2804.600 ;
        RECT 539.030 2801.750 539.330 2804.600 ;
        RECT 544.250 2801.750 544.550 2804.600 ;
        RECT 539.030 2801.450 542.490 2801.750 ;
        RECT 539.030 2800.000 539.330 2801.450 ;
        RECT 538.410 2796.350 538.810 2796.650 ;
        RECT 538.510 2794.625 538.810 2796.350 ;
        RECT 542.190 2794.625 542.490 2801.450 ;
        RECT 543.110 2801.450 544.550 2801.750 ;
        RECT 535.735 2794.295 536.065 2794.625 ;
        RECT 538.495 2794.295 538.825 2794.625 ;
        RECT 542.175 2794.295 542.505 2794.625 ;
        RECT 531.135 2793.615 531.465 2793.945 ;
        RECT 543.110 2793.265 543.410 2801.450 ;
        RECT 544.250 2800.000 544.550 2801.450 ;
        RECT 544.870 2801.750 545.170 2804.600 ;
        RECT 984.010 2801.750 984.310 2804.600 ;
        RECT 989.850 2801.750 990.150 2804.600 ;
        RECT 995.690 2801.750 995.990 2804.600 ;
        RECT 1001.530 2801.750 1001.830 2804.600 ;
        RECT 544.870 2801.450 548.010 2801.750 ;
        RECT 544.870 2800.000 545.170 2801.450 ;
        RECT 547.710 2794.625 548.010 2801.450 ;
        RECT 981.030 2801.450 984.310 2801.750 ;
        RECT 981.030 2794.625 981.330 2801.450 ;
        RECT 984.010 2800.000 984.310 2801.450 ;
        RECT 987.470 2801.450 990.150 2801.750 ;
        RECT 547.695 2794.295 548.025 2794.625 ;
        RECT 981.015 2794.295 981.345 2794.625 ;
        RECT 987.470 2793.945 987.770 2801.450 ;
        RECT 989.850 2800.000 990.150 2801.450 ;
        RECT 993.910 2801.450 995.990 2801.750 ;
        RECT 987.455 2793.615 987.785 2793.945 ;
        RECT 501.695 2792.935 502.025 2793.265 ;
        RECT 520.095 2792.935 520.425 2793.265 ;
        RECT 543.095 2792.935 543.425 2793.265 ;
        RECT 348.975 2792.255 349.305 2792.585 ;
        RECT 993.910 2791.225 994.210 2801.450 ;
        RECT 995.690 2800.000 995.990 2801.450 ;
        RECT 1001.270 2800.000 1001.830 2801.750 ;
        RECT 1007.370 2800.050 1007.670 2804.600 ;
        RECT 1013.210 2801.750 1013.510 2804.600 ;
        RECT 1012.310 2801.450 1013.510 2801.750 ;
        RECT 1001.270 2793.945 1001.570 2800.000 ;
        RECT 1007.370 2799.750 1008.010 2800.050 ;
        RECT 1001.255 2793.615 1001.585 2793.945 ;
        RECT 993.895 2790.895 994.225 2791.225 ;
        RECT 1007.710 2788.505 1008.010 2799.750 ;
        RECT 1012.310 2793.265 1012.610 2801.450 ;
        RECT 1013.210 2800.000 1013.510 2801.450 ;
        RECT 1013.830 2796.650 1014.130 2804.600 ;
        RECT 1019.050 2801.750 1019.350 2804.600 ;
        RECT 1013.230 2796.350 1014.130 2796.650 ;
        RECT 1018.750 2800.000 1019.350 2801.750 ;
        RECT 1013.230 2794.625 1013.530 2796.350 ;
        RECT 1018.750 2794.625 1019.050 2800.000 ;
        RECT 1019.670 2794.625 1019.970 2804.600 ;
        RECT 1024.890 2801.750 1025.190 2804.600 ;
        RECT 1024.270 2801.450 1025.190 2801.750 ;
        RECT 1013.215 2794.295 1013.545 2794.625 ;
        RECT 1018.735 2794.295 1019.065 2794.625 ;
        RECT 1019.655 2794.295 1019.985 2794.625 ;
        RECT 1024.270 2793.265 1024.570 2801.450 ;
        RECT 1024.890 2800.000 1025.190 2801.450 ;
        RECT 1025.510 2801.750 1025.810 2804.600 ;
        RECT 1030.730 2801.750 1031.030 2804.600 ;
        RECT 1025.510 2801.450 1027.330 2801.750 ;
        RECT 1025.510 2800.000 1025.810 2801.450 ;
        RECT 1027.030 2794.625 1027.330 2801.450 ;
        RECT 1030.710 2800.000 1031.030 2801.750 ;
        RECT 1031.350 2801.750 1031.650 2804.600 ;
        RECT 1036.570 2802.450 1036.870 2804.600 ;
        RECT 1035.310 2802.150 1036.870 2802.450 ;
        RECT 1031.350 2801.450 1034.690 2801.750 ;
        RECT 1031.350 2800.000 1031.650 2801.450 ;
        RECT 1030.710 2794.625 1031.010 2800.000 ;
        RECT 1027.015 2794.295 1027.345 2794.625 ;
        RECT 1030.695 2794.295 1031.025 2794.625 ;
        RECT 1012.295 2792.935 1012.625 2793.265 ;
        RECT 1024.255 2792.935 1024.585 2793.265 ;
        RECT 1007.695 2788.175 1008.025 2788.505 ;
        RECT 1034.390 2787.825 1034.690 2801.450 ;
        RECT 1035.310 2788.505 1035.610 2802.150 ;
        RECT 1036.570 2800.000 1036.870 2802.150 ;
        RECT 1037.190 2801.750 1037.490 2804.600 ;
        RECT 1042.410 2801.750 1042.710 2804.600 ;
        RECT 1037.190 2801.450 1040.210 2801.750 ;
        RECT 1037.190 2800.000 1037.490 2801.450 ;
        RECT 1035.295 2788.175 1035.625 2788.505 ;
        RECT 1039.910 2787.825 1040.210 2801.450 ;
        RECT 1041.750 2801.450 1042.710 2801.750 ;
        RECT 1041.750 2794.625 1042.050 2801.450 ;
        RECT 1042.410 2800.000 1042.710 2801.450 ;
        RECT 1043.030 2801.750 1043.330 2804.600 ;
        RECT 1048.250 2801.750 1048.550 2804.600 ;
        RECT 1043.030 2801.450 1046.650 2801.750 ;
        RECT 1043.030 2800.000 1043.330 2801.450 ;
        RECT 1041.735 2794.295 1042.065 2794.625 ;
        RECT 1046.350 2787.825 1046.650 2801.450 ;
        RECT 1048.190 2800.000 1048.550 2801.750 ;
        RECT 1048.870 2801.750 1049.170 2804.600 ;
        RECT 1054.090 2802.450 1054.390 2804.600 ;
        RECT 1052.790 2802.150 1054.390 2802.450 ;
        RECT 1048.870 2801.450 1052.170 2801.750 ;
        RECT 1048.870 2800.000 1049.170 2801.450 ;
        RECT 1048.190 2793.265 1048.490 2800.000 ;
        RECT 1048.175 2792.935 1048.505 2793.265 ;
        RECT 1051.870 2788.505 1052.170 2801.450 ;
        RECT 1052.790 2795.985 1053.090 2802.150 ;
        RECT 1054.090 2800.000 1054.390 2802.150 ;
        RECT 1054.710 2800.050 1055.010 2804.600 ;
        RECT 1059.930 2801.750 1060.230 2804.600 ;
        RECT 1059.230 2801.450 1060.230 2801.750 ;
        RECT 1055.535 2800.050 1055.865 2800.065 ;
        RECT 1054.710 2799.750 1055.865 2800.050 ;
        RECT 1055.535 2799.735 1055.865 2799.750 ;
        RECT 1052.775 2795.655 1053.105 2795.985 ;
        RECT 1059.230 2794.625 1059.530 2801.450 ;
        RECT 1059.930 2800.000 1060.230 2801.450 ;
        RECT 1060.550 2801.750 1060.850 2804.600 ;
        RECT 1065.770 2801.750 1066.070 2804.600 ;
        RECT 1060.550 2801.450 1062.290 2801.750 ;
        RECT 1060.550 2800.000 1060.850 2801.450 ;
        RECT 1059.215 2794.295 1059.545 2794.625 ;
        RECT 1051.855 2788.175 1052.185 2788.505 ;
        RECT 1061.990 2787.825 1062.290 2801.450 ;
        RECT 1065.670 2800.000 1066.070 2801.750 ;
        RECT 1066.390 2801.750 1066.690 2804.600 ;
        RECT 1071.610 2801.750 1071.910 2804.600 ;
        RECT 1066.390 2801.450 1067.810 2801.750 ;
        RECT 1066.390 2800.000 1066.690 2801.450 ;
        RECT 1065.670 2794.625 1065.970 2800.000 ;
        RECT 1065.655 2794.295 1065.985 2794.625 ;
        RECT 1067.510 2787.825 1067.810 2801.450 ;
        RECT 1070.270 2801.450 1071.910 2801.750 ;
        RECT 1070.270 2794.625 1070.570 2801.450 ;
        RECT 1071.610 2800.000 1071.910 2801.450 ;
        RECT 1072.230 2801.750 1072.530 2804.600 ;
        RECT 1077.450 2801.750 1077.750 2804.600 ;
        RECT 1072.230 2801.450 1074.250 2801.750 ;
        RECT 1072.230 2800.000 1072.530 2801.450 ;
        RECT 1070.255 2794.295 1070.585 2794.625 ;
        RECT 1073.950 2787.825 1074.250 2801.450 ;
        RECT 1076.710 2801.450 1077.750 2801.750 ;
        RECT 1076.710 2793.945 1077.010 2801.450 ;
        RECT 1077.450 2800.000 1077.750 2801.450 ;
        RECT 1078.070 2801.750 1078.370 2804.600 ;
        RECT 1083.290 2801.750 1083.590 2804.600 ;
        RECT 1078.070 2801.450 1081.610 2801.750 ;
        RECT 1078.070 2800.000 1078.370 2801.450 ;
        RECT 1081.310 2794.625 1081.610 2801.450 ;
        RECT 1083.150 2800.000 1083.590 2801.750 ;
        RECT 1083.910 2801.750 1084.210 2804.600 ;
        RECT 1089.130 2801.750 1089.430 2804.600 ;
        RECT 1083.910 2801.450 1087.130 2801.750 ;
        RECT 1083.910 2800.000 1084.210 2801.450 ;
        RECT 1081.295 2794.295 1081.625 2794.625 ;
        RECT 1083.150 2793.945 1083.450 2800.000 ;
        RECT 1086.830 2793.945 1087.130 2801.450 ;
        RECT 1087.750 2801.450 1089.430 2801.750 ;
        RECT 1087.750 2794.625 1088.050 2801.450 ;
        RECT 1089.130 2800.000 1089.430 2801.450 ;
        RECT 1089.750 2796.650 1090.050 2804.600 ;
        RECT 1094.970 2801.750 1095.270 2804.600 ;
        RECT 1089.590 2796.350 1090.050 2796.650 ;
        RECT 1094.190 2801.450 1095.270 2801.750 ;
        RECT 1089.590 2794.625 1089.890 2796.350 ;
        RECT 1094.190 2794.625 1094.490 2801.450 ;
        RECT 1094.970 2800.000 1095.270 2801.450 ;
        RECT 1095.590 2800.050 1095.890 2804.600 ;
        RECT 1100.810 2801.750 1101.110 2804.600 ;
        RECT 1095.590 2799.750 1096.330 2800.050 ;
        RECT 1096.030 2794.625 1096.330 2799.750 ;
        RECT 1100.630 2800.000 1101.110 2801.750 ;
        RECT 1101.430 2801.750 1101.730 2804.600 ;
        RECT 1106.650 2802.450 1106.950 2804.600 ;
        RECT 1105.230 2802.150 1106.950 2802.450 ;
        RECT 1101.430 2801.450 1103.690 2801.750 ;
        RECT 1101.430 2800.000 1101.730 2801.450 ;
        RECT 1100.630 2794.625 1100.930 2800.000 ;
        RECT 1103.390 2794.625 1103.690 2801.450 ;
        RECT 1105.230 2794.625 1105.530 2802.150 ;
        RECT 1106.650 2800.000 1106.950 2802.150 ;
        RECT 1107.270 2801.750 1107.570 2804.600 ;
        RECT 1112.490 2801.750 1112.790 2804.600 ;
        RECT 1107.270 2801.450 1110.130 2801.750 ;
        RECT 1107.270 2800.000 1107.570 2801.450 ;
        RECT 1109.830 2794.625 1110.130 2801.450 ;
        RECT 1111.670 2801.450 1112.790 2801.750 ;
        RECT 1111.670 2794.625 1111.970 2801.450 ;
        RECT 1112.490 2800.000 1112.790 2801.450 ;
        RECT 1113.110 2801.750 1113.410 2804.600 ;
        RECT 1118.330 2801.750 1118.630 2804.600 ;
        RECT 1113.110 2801.450 1116.570 2801.750 ;
        RECT 1113.110 2800.000 1113.410 2801.450 ;
        RECT 1087.735 2794.295 1088.065 2794.625 ;
        RECT 1089.575 2794.295 1089.905 2794.625 ;
        RECT 1094.175 2794.295 1094.505 2794.625 ;
        RECT 1096.015 2794.295 1096.345 2794.625 ;
        RECT 1100.615 2794.295 1100.945 2794.625 ;
        RECT 1103.375 2794.295 1103.705 2794.625 ;
        RECT 1105.215 2794.295 1105.545 2794.625 ;
        RECT 1109.815 2794.295 1110.145 2794.625 ;
        RECT 1111.655 2794.295 1111.985 2794.625 ;
        RECT 1076.695 2793.615 1077.025 2793.945 ;
        RECT 1083.135 2793.615 1083.465 2793.945 ;
        RECT 1086.815 2793.615 1087.145 2793.945 ;
        RECT 1116.270 2792.585 1116.570 2801.450 ;
        RECT 1118.110 2800.000 1118.630 2801.750 ;
        RECT 1118.950 2801.750 1119.250 2804.600 ;
        RECT 1124.170 2801.750 1124.470 2804.600 ;
        RECT 1118.950 2801.450 1122.090 2801.750 ;
        RECT 1118.950 2800.000 1119.250 2801.450 ;
        RECT 1118.110 2794.625 1118.410 2800.000 ;
        RECT 1121.790 2794.625 1122.090 2801.450 ;
        RECT 1122.710 2801.450 1124.470 2801.750 ;
        RECT 1118.095 2794.295 1118.425 2794.625 ;
        RECT 1121.775 2794.295 1122.105 2794.625 ;
        RECT 1122.710 2793.945 1123.010 2801.450 ;
        RECT 1124.170 2800.000 1124.470 2801.450 ;
        RECT 1124.790 2801.750 1125.090 2804.600 ;
        RECT 1130.010 2801.750 1130.310 2804.600 ;
        RECT 1124.790 2801.450 1128.530 2801.750 ;
        RECT 1124.790 2800.000 1125.090 2801.450 ;
        RECT 1128.230 2793.945 1128.530 2801.450 ;
        RECT 1129.150 2801.450 1130.310 2801.750 ;
        RECT 1129.150 2794.625 1129.450 2801.450 ;
        RECT 1130.010 2800.000 1130.310 2801.450 ;
        RECT 1130.630 2800.050 1130.930 2804.600 ;
        RECT 1135.850 2801.750 1136.150 2804.600 ;
        RECT 1130.630 2799.750 1131.290 2800.050 ;
        RECT 1130.990 2794.625 1131.290 2799.750 ;
        RECT 1135.590 2800.000 1136.150 2801.750 ;
        RECT 1136.470 2801.750 1136.770 2804.600 ;
        RECT 1141.690 2802.450 1141.990 2804.600 ;
        RECT 1140.190 2802.150 1141.990 2802.450 ;
        RECT 1136.470 2801.450 1137.730 2801.750 ;
        RECT 1136.470 2800.000 1136.770 2801.450 ;
        RECT 1135.590 2794.625 1135.890 2800.000 ;
        RECT 1137.430 2794.625 1137.730 2801.450 ;
        RECT 1140.190 2794.625 1140.490 2802.150 ;
        RECT 1141.690 2800.000 1141.990 2802.150 ;
        RECT 1142.310 2801.750 1142.610 2804.600 ;
        RECT 1147.530 2801.750 1147.830 2804.600 ;
        RECT 1142.310 2801.450 1144.170 2801.750 ;
        RECT 1142.310 2800.000 1142.610 2801.450 ;
        RECT 1143.870 2794.625 1144.170 2801.450 ;
        RECT 1146.630 2801.450 1147.830 2801.750 ;
        RECT 1146.630 2794.625 1146.930 2801.450 ;
        RECT 1147.530 2800.000 1147.830 2801.450 ;
        RECT 1148.150 2801.750 1148.450 2804.600 ;
        RECT 1153.370 2801.750 1153.670 2804.600 ;
        RECT 1148.150 2801.450 1151.530 2801.750 ;
        RECT 1148.150 2800.000 1148.450 2801.450 ;
        RECT 1151.230 2794.625 1151.530 2801.450 ;
        RECT 1153.070 2800.000 1153.670 2801.750 ;
        RECT 1129.135 2794.295 1129.465 2794.625 ;
        RECT 1130.975 2794.295 1131.305 2794.625 ;
        RECT 1135.575 2794.295 1135.905 2794.625 ;
        RECT 1137.415 2794.295 1137.745 2794.625 ;
        RECT 1140.175 2794.295 1140.505 2794.625 ;
        RECT 1143.855 2794.295 1144.185 2794.625 ;
        RECT 1146.615 2794.295 1146.945 2794.625 ;
        RECT 1151.215 2794.295 1151.545 2794.625 ;
        RECT 1122.695 2793.615 1123.025 2793.945 ;
        RECT 1128.215 2793.615 1128.545 2793.945 ;
        RECT 1153.070 2792.585 1153.370 2800.000 ;
        RECT 1153.990 2794.625 1154.290 2804.600 ;
        RECT 1159.210 2796.650 1159.510 2804.600 ;
        RECT 1159.830 2801.750 1160.130 2804.600 ;
        RECT 1165.050 2801.750 1165.350 2804.600 ;
        RECT 1159.830 2801.450 1163.490 2801.750 ;
        RECT 1159.830 2800.000 1160.130 2801.450 ;
        RECT 1159.210 2796.350 1159.810 2796.650 ;
        RECT 1153.975 2794.295 1154.305 2794.625 ;
        RECT 1116.255 2792.255 1116.585 2792.585 ;
        RECT 1153.055 2792.255 1153.385 2792.585 ;
        RECT 1159.510 2791.905 1159.810 2796.350 ;
        RECT 1163.190 2793.945 1163.490 2801.450 ;
        RECT 1164.110 2801.450 1165.350 2801.750 ;
        RECT 1163.175 2793.615 1163.505 2793.945 ;
        RECT 1159.495 2791.575 1159.825 2791.905 ;
        RECT 1164.110 2791.225 1164.410 2801.450 ;
        RECT 1165.050 2800.000 1165.350 2801.450 ;
        RECT 1165.670 2796.650 1165.970 2804.600 ;
        RECT 1170.890 2801.750 1171.190 2804.600 ;
        RECT 1165.030 2796.350 1165.970 2796.650 ;
        RECT 1167.790 2801.450 1171.190 2801.750 ;
        RECT 1165.030 2794.625 1165.330 2796.350 ;
        RECT 1165.015 2794.295 1165.345 2794.625 ;
        RECT 1167.790 2793.265 1168.090 2801.450 ;
        RECT 1170.890 2800.000 1171.190 2801.450 ;
        RECT 1171.510 2801.750 1171.810 2804.600 ;
        RECT 1176.730 2801.750 1177.030 2804.600 ;
        RECT 1171.510 2801.450 1172.690 2801.750 ;
        RECT 1171.510 2800.000 1171.810 2801.450 ;
        RECT 1172.390 2794.625 1172.690 2801.450 ;
        RECT 1173.310 2801.450 1177.030 2801.750 ;
        RECT 1172.375 2794.295 1172.705 2794.625 ;
        RECT 1173.310 2793.945 1173.610 2801.450 ;
        RECT 1176.730 2800.000 1177.030 2801.450 ;
        RECT 1177.350 2801.750 1177.650 2804.600 ;
        RECT 1182.570 2801.750 1182.870 2804.600 ;
        RECT 1177.350 2801.450 1179.130 2801.750 ;
        RECT 1177.350 2800.000 1177.650 2801.450 ;
        RECT 1178.830 2794.625 1179.130 2801.450 ;
        RECT 1180.670 2801.450 1182.870 2801.750 ;
        RECT 1178.815 2794.295 1179.145 2794.625 ;
        RECT 1180.670 2793.945 1180.970 2801.450 ;
        RECT 1182.570 2800.000 1182.870 2801.450 ;
        RECT 1183.190 2801.750 1183.490 2804.600 ;
        RECT 1188.410 2801.750 1188.710 2804.600 ;
        RECT 1183.190 2801.450 1186.490 2801.750 ;
        RECT 1183.190 2800.000 1183.490 2801.450 ;
        RECT 1186.190 2794.625 1186.490 2801.450 ;
        RECT 1187.110 2801.450 1188.710 2801.750 ;
        RECT 1186.175 2794.295 1186.505 2794.625 ;
        RECT 1187.110 2793.945 1187.410 2801.450 ;
        RECT 1188.410 2800.000 1188.710 2801.450 ;
        RECT 1189.030 2801.750 1189.330 2804.600 ;
        RECT 1194.250 2801.750 1194.550 2804.600 ;
        RECT 1189.030 2801.450 1192.010 2801.750 ;
        RECT 1189.030 2800.000 1189.330 2801.450 ;
        RECT 1173.295 2793.615 1173.625 2793.945 ;
        RECT 1180.655 2793.615 1180.985 2793.945 ;
        RECT 1187.095 2793.615 1187.425 2793.945 ;
        RECT 1167.775 2792.935 1168.105 2793.265 ;
        RECT 1164.095 2790.895 1164.425 2791.225 ;
        RECT 1191.710 2790.545 1192.010 2801.450 ;
        RECT 1193.550 2801.450 1194.550 2801.750 ;
        RECT 1193.550 2791.905 1193.850 2801.450 ;
        RECT 1194.250 2800.000 1194.550 2801.450 ;
        RECT 1194.870 2801.750 1195.170 2804.600 ;
        RECT 1584.010 2801.750 1584.310 2804.600 ;
        RECT 1589.850 2801.750 1590.150 2804.600 ;
        RECT 1595.690 2801.750 1595.990 2804.600 ;
        RECT 1194.870 2801.450 1198.450 2801.750 ;
        RECT 1194.870 2800.000 1195.170 2801.450 ;
        RECT 1198.150 2794.625 1198.450 2801.450 ;
        RECT 1580.870 2801.450 1584.310 2801.750 ;
        RECT 1198.135 2794.295 1198.465 2794.625 ;
        RECT 1193.535 2791.575 1193.865 2791.905 ;
        RECT 1417.095 2790.895 1417.425 2791.225 ;
        RECT 1191.695 2790.215 1192.025 2790.545 ;
        RECT 1034.375 2787.495 1034.705 2787.825 ;
        RECT 1039.895 2787.495 1040.225 2787.825 ;
        RECT 1046.335 2787.495 1046.665 2787.825 ;
        RECT 1061.975 2787.495 1062.305 2787.825 ;
        RECT 1067.495 2787.495 1067.825 2787.825 ;
        RECT 1073.935 2787.495 1074.265 2787.825 ;
        RECT 292.020 2715.000 295.020 2785.000 ;
        RECT 310.020 2715.000 313.020 2785.000 ;
        RECT 328.020 2715.000 331.020 2785.000 ;
        RECT 364.020 2715.000 367.020 2785.000 ;
        RECT 454.020 2715.000 457.020 2785.000 ;
        RECT 472.020 2715.000 475.020 2785.000 ;
        RECT 490.020 2715.000 493.020 2785.000 ;
        RECT 508.020 2715.000 511.020 2785.000 ;
        RECT 544.020 2715.000 547.020 2785.000 ;
        RECT 634.020 2715.000 637.020 2785.000 ;
        RECT 652.020 2715.000 655.020 2785.000 ;
        RECT 670.020 2715.000 673.020 2785.000 ;
        RECT 688.020 2715.000 691.020 2785.000 ;
        RECT 994.020 2715.000 997.020 2785.000 ;
        RECT 1012.020 2715.000 1015.020 2785.000 ;
        RECT 1030.020 2715.000 1033.020 2785.000 ;
        RECT 1048.020 2715.000 1051.020 2785.000 ;
        RECT 1084.020 2715.000 1087.020 2785.000 ;
        RECT 1174.020 2715.000 1177.020 2785.000 ;
        RECT 1192.020 2715.000 1195.020 2785.000 ;
        RECT 1210.020 2715.000 1213.020 2785.000 ;
        RECT 1228.020 2715.000 1231.020 2785.000 ;
        RECT 1264.020 2715.000 1267.020 2785.000 ;
      LAYER met4 ;
        RECT 325.065 1610.640 397.370 2688.240 ;
        RECT 399.770 1610.640 1388.915 2688.240 ;
      LAYER met4 ;
        RECT 1410.655 2087.095 1410.985 2087.425 ;
        RECT 1410.670 1657.665 1410.970 2087.095 ;
        RECT 1410.655 1657.335 1410.985 1657.665 ;
        RECT 1417.110 1627.745 1417.410 2790.895 ;
        RECT 1580.870 2787.825 1581.170 2801.450 ;
        RECT 1584.010 2800.000 1584.310 2801.450 ;
        RECT 1587.310 2801.450 1590.150 2801.750 ;
        RECT 1587.310 2791.905 1587.610 2801.450 ;
        RECT 1589.850 2800.000 1590.150 2801.450 ;
        RECT 1594.670 2801.450 1595.990 2801.750 ;
        RECT 1587.295 2791.575 1587.625 2791.905 ;
        RECT 1594.670 2787.825 1594.970 2801.450 ;
        RECT 1595.690 2800.000 1595.990 2801.450 ;
        RECT 1601.530 2802.450 1601.830 2804.600 ;
        RECT 1601.530 2802.150 1603.250 2802.450 ;
        RECT 1601.530 2800.000 1601.830 2802.150 ;
        RECT 1602.950 2791.905 1603.250 2802.150 ;
        RECT 1607.370 2801.750 1607.670 2804.600 ;
        RECT 1613.210 2801.750 1613.510 2804.600 ;
        RECT 1604.790 2801.450 1607.670 2801.750 ;
        RECT 1602.935 2791.575 1603.265 2791.905 ;
        RECT 1604.790 2787.825 1605.090 2801.450 ;
        RECT 1607.370 2800.000 1607.670 2801.450 ;
        RECT 1613.070 2800.000 1613.510 2801.750 ;
        RECT 1613.830 2801.750 1614.130 2804.600 ;
        RECT 1613.830 2800.000 1614.290 2801.750 ;
        RECT 1619.050 2800.050 1619.350 2804.600 ;
        RECT 1613.070 2794.625 1613.370 2800.000 ;
        RECT 1613.055 2794.295 1613.385 2794.625 ;
        RECT 1613.990 2787.825 1614.290 2800.000 ;
        RECT 1618.590 2799.750 1619.350 2800.050 ;
        RECT 1619.670 2801.750 1619.970 2804.600 ;
        RECT 1624.890 2801.750 1625.190 2804.600 ;
        RECT 1619.670 2801.450 1620.730 2801.750 ;
        RECT 1619.670 2800.000 1619.970 2801.450 ;
        RECT 1618.590 2788.505 1618.890 2799.750 ;
        RECT 1618.575 2788.175 1618.905 2788.505 ;
        RECT 1620.430 2787.825 1620.730 2801.450 ;
        RECT 1624.110 2801.450 1625.190 2801.750 ;
        RECT 1624.110 2788.505 1624.410 2801.450 ;
        RECT 1624.890 2800.000 1625.190 2801.450 ;
        RECT 1625.510 2802.450 1625.810 2804.600 ;
        RECT 1625.510 2802.150 1627.170 2802.450 ;
        RECT 1625.510 2800.000 1625.810 2802.150 ;
        RECT 1624.095 2788.175 1624.425 2788.505 ;
        RECT 1626.870 2787.825 1627.170 2802.150 ;
        RECT 1630.730 2801.750 1631.030 2804.600 ;
        RECT 1630.550 2800.000 1631.030 2801.750 ;
        RECT 1631.350 2801.750 1631.650 2804.600 ;
        RECT 1631.350 2800.000 1631.770 2801.750 ;
        RECT 1636.570 2800.050 1636.870 2804.600 ;
        RECT 1630.550 2787.825 1630.850 2800.000 ;
        RECT 1631.470 2788.505 1631.770 2800.000 ;
        RECT 1636.070 2799.750 1636.870 2800.050 ;
        RECT 1637.190 2801.750 1637.490 2804.600 ;
        RECT 1637.190 2801.450 1638.210 2801.750 ;
        RECT 1637.190 2800.000 1637.490 2801.450 ;
        RECT 1636.070 2796.650 1636.370 2799.750 ;
        RECT 1636.070 2796.350 1637.290 2796.650 ;
        RECT 1636.990 2793.265 1637.290 2796.350 ;
        RECT 1636.975 2792.935 1637.305 2793.265 ;
        RECT 1637.910 2792.585 1638.210 2801.450 ;
        RECT 1642.410 2796.650 1642.710 2804.600 ;
        RECT 1643.030 2802.450 1643.330 2804.600 ;
        RECT 1643.030 2802.150 1644.650 2802.450 ;
        RECT 1643.030 2800.000 1643.330 2802.150 ;
        RECT 1642.410 2796.350 1642.810 2796.650 ;
        RECT 1642.510 2794.625 1642.810 2796.350 ;
        RECT 1642.495 2794.295 1642.825 2794.625 ;
        RECT 1637.895 2792.255 1638.225 2792.585 ;
        RECT 1644.350 2790.545 1644.650 2802.150 ;
        RECT 1648.250 2801.750 1648.550 2804.600 ;
        RECT 1648.030 2800.000 1648.550 2801.750 ;
        RECT 1648.870 2801.750 1649.170 2804.600 ;
        RECT 1654.090 2802.450 1654.390 2804.600 ;
        RECT 1652.630 2802.150 1654.390 2802.450 ;
        RECT 1648.870 2800.000 1649.250 2801.750 ;
        RECT 1644.335 2790.215 1644.665 2790.545 ;
        RECT 1648.030 2789.865 1648.330 2800.000 ;
        RECT 1648.015 2789.535 1648.345 2789.865 ;
        RECT 1631.455 2788.175 1631.785 2788.505 ;
        RECT 1648.950 2787.825 1649.250 2800.000 ;
        RECT 1652.630 2794.625 1652.930 2802.150 ;
        RECT 1654.090 2800.000 1654.390 2802.150 ;
        RECT 1654.710 2801.750 1655.010 2804.600 ;
        RECT 1659.930 2801.750 1660.230 2804.600 ;
        RECT 1654.710 2801.450 1655.690 2801.750 ;
        RECT 1654.710 2800.000 1655.010 2801.450 ;
        RECT 1652.615 2794.295 1652.945 2794.625 ;
        RECT 1655.390 2788.505 1655.690 2801.450 ;
        RECT 1659.070 2801.450 1660.230 2801.750 ;
        RECT 1659.070 2794.625 1659.370 2801.450 ;
        RECT 1659.930 2800.000 1660.230 2801.450 ;
        RECT 1660.550 2800.050 1660.850 2804.600 ;
        RECT 1665.770 2801.750 1666.070 2804.600 ;
        RECT 1660.550 2799.750 1661.210 2800.050 ;
        RECT 1659.055 2794.295 1659.385 2794.625 ;
        RECT 1655.375 2788.175 1655.705 2788.505 ;
        RECT 1660.910 2787.825 1661.210 2799.750 ;
        RECT 1665.510 2800.000 1666.070 2801.750 ;
        RECT 1666.390 2801.750 1666.690 2804.600 ;
        RECT 1671.610 2802.450 1671.910 2804.600 ;
        RECT 1670.110 2802.150 1671.910 2802.450 ;
        RECT 1666.390 2800.000 1666.730 2801.750 ;
        RECT 1665.510 2794.625 1665.810 2800.000 ;
        RECT 1665.495 2794.295 1665.825 2794.625 ;
        RECT 1666.430 2787.825 1666.730 2800.000 ;
        RECT 1670.110 2794.625 1670.410 2802.150 ;
        RECT 1671.610 2800.000 1671.910 2802.150 ;
        RECT 1672.230 2801.750 1672.530 2804.600 ;
        RECT 1672.230 2801.450 1673.170 2801.750 ;
        RECT 1672.230 2800.000 1672.530 2801.450 ;
        RECT 1670.095 2794.295 1670.425 2794.625 ;
        RECT 1672.870 2787.825 1673.170 2801.450 ;
        RECT 1677.450 2800.050 1677.750 2804.600 ;
        RECT 1678.070 2800.050 1678.370 2804.600 ;
        RECT 1683.290 2801.750 1683.590 2804.600 ;
        RECT 1681.150 2801.450 1683.590 2801.750 ;
        RECT 1677.450 2799.750 1677.770 2800.050 ;
        RECT 1678.070 2799.750 1678.690 2800.050 ;
        RECT 1677.470 2794.625 1677.770 2799.750 ;
        RECT 1677.455 2794.295 1677.785 2794.625 ;
        RECT 1678.390 2787.825 1678.690 2799.750 ;
        RECT 1681.150 2793.265 1681.450 2801.450 ;
        RECT 1683.290 2800.000 1683.590 2801.450 ;
        RECT 1681.135 2792.935 1681.465 2793.265 ;
        RECT 1683.910 2787.825 1684.210 2804.600 ;
        RECT 1689.130 2801.750 1689.430 2804.600 ;
        RECT 1688.510 2801.450 1689.430 2801.750 ;
        RECT 1688.510 2793.945 1688.810 2801.450 ;
        RECT 1689.130 2800.000 1689.430 2801.450 ;
        RECT 1689.750 2796.650 1690.050 2804.600 ;
        RECT 1694.970 2801.750 1695.270 2804.600 ;
        RECT 1689.430 2796.350 1690.050 2796.650 ;
        RECT 1694.950 2800.000 1695.270 2801.750 ;
        RECT 1695.590 2801.750 1695.890 2804.600 ;
        RECT 1700.810 2802.450 1701.110 2804.600 ;
        RECT 1699.550 2802.150 1701.110 2802.450 ;
        RECT 1695.590 2800.000 1696.170 2801.750 ;
        RECT 1688.495 2793.615 1688.825 2793.945 ;
        RECT 1689.430 2788.505 1689.730 2796.350 ;
        RECT 1694.950 2794.625 1695.250 2800.000 ;
        RECT 1694.935 2794.295 1695.265 2794.625 ;
        RECT 1689.415 2788.175 1689.745 2788.505 ;
        RECT 1695.870 2787.825 1696.170 2800.000 ;
        RECT 1699.550 2794.625 1699.850 2802.150 ;
        RECT 1700.810 2800.000 1701.110 2802.150 ;
        RECT 1701.430 2801.750 1701.730 2804.600 ;
        RECT 1706.650 2801.750 1706.950 2804.600 ;
        RECT 1701.430 2801.450 1702.610 2801.750 ;
        RECT 1701.430 2800.000 1701.730 2801.450 ;
        RECT 1699.535 2794.295 1699.865 2794.625 ;
        RECT 1702.310 2787.825 1702.610 2801.450 ;
        RECT 1705.990 2801.450 1706.950 2801.750 ;
        RECT 1705.990 2794.625 1706.290 2801.450 ;
        RECT 1706.650 2800.000 1706.950 2801.450 ;
        RECT 1707.270 2802.450 1707.570 2804.600 ;
        RECT 1707.270 2802.150 1709.050 2802.450 ;
        RECT 1707.270 2800.000 1707.570 2802.150 ;
        RECT 1705.975 2794.295 1706.305 2794.625 ;
        RECT 1708.750 2787.825 1709.050 2802.150 ;
        RECT 1712.490 2801.750 1712.790 2804.600 ;
        RECT 1712.430 2800.000 1712.790 2801.750 ;
        RECT 1713.110 2801.750 1713.410 2804.600 ;
        RECT 1713.110 2800.000 1713.650 2801.750 ;
        RECT 1718.330 2800.050 1718.630 2804.600 ;
        RECT 1712.430 2794.625 1712.730 2800.000 ;
        RECT 1712.415 2794.295 1712.745 2794.625 ;
        RECT 1713.350 2787.825 1713.650 2800.000 ;
        RECT 1717.950 2799.750 1718.630 2800.050 ;
        RECT 1718.950 2801.750 1719.250 2804.600 ;
        RECT 1724.170 2801.750 1724.470 2804.600 ;
        RECT 1718.950 2801.450 1720.090 2801.750 ;
        RECT 1718.950 2800.000 1719.250 2801.450 ;
        RECT 1717.950 2794.625 1718.250 2799.750 ;
        RECT 1717.935 2794.295 1718.265 2794.625 ;
        RECT 1719.790 2787.825 1720.090 2801.450 ;
        RECT 1723.470 2801.450 1724.470 2801.750 ;
        RECT 1723.470 2794.625 1723.770 2801.450 ;
        RECT 1724.170 2800.000 1724.470 2801.450 ;
        RECT 1724.790 2796.650 1725.090 2804.600 ;
        RECT 1730.010 2801.750 1730.310 2804.600 ;
        RECT 1724.390 2796.350 1725.090 2796.650 ;
        RECT 1728.990 2801.450 1730.310 2801.750 ;
        RECT 1723.455 2794.295 1723.785 2794.625 ;
        RECT 1724.390 2788.505 1724.690 2796.350 ;
        RECT 1728.990 2794.625 1729.290 2801.450 ;
        RECT 1730.010 2800.000 1730.310 2801.450 ;
        RECT 1730.630 2801.750 1730.930 2804.600 ;
        RECT 1735.850 2801.750 1736.150 2804.600 ;
        RECT 1730.630 2800.000 1731.130 2801.750 ;
        RECT 1728.975 2794.295 1729.305 2794.625 ;
        RECT 1724.375 2788.175 1724.705 2788.505 ;
        RECT 1730.830 2787.825 1731.130 2800.000 ;
        RECT 1732.670 2801.450 1736.150 2801.750 ;
        RECT 1732.670 2795.985 1732.970 2801.450 ;
        RECT 1735.850 2800.000 1736.150 2801.450 ;
        RECT 1736.470 2801.750 1736.770 2804.600 ;
        RECT 1741.690 2801.750 1741.990 2804.600 ;
        RECT 1736.470 2801.450 1737.570 2801.750 ;
        RECT 1736.470 2800.000 1736.770 2801.450 ;
        RECT 1732.655 2795.655 1732.985 2795.985 ;
        RECT 1737.270 2787.825 1737.570 2801.450 ;
        RECT 1740.950 2801.450 1741.990 2801.750 ;
        RECT 1740.950 2794.625 1741.250 2801.450 ;
        RECT 1741.690 2800.000 1741.990 2801.450 ;
        RECT 1742.310 2802.450 1742.610 2804.600 ;
        RECT 1742.310 2802.150 1744.010 2802.450 ;
        RECT 1742.310 2800.000 1742.610 2802.150 ;
        RECT 1740.935 2794.295 1741.265 2794.625 ;
        RECT 1743.710 2787.825 1744.010 2802.150 ;
        RECT 1747.530 2801.750 1747.830 2804.600 ;
        RECT 1747.390 2800.000 1747.830 2801.750 ;
        RECT 1748.150 2801.750 1748.450 2804.600 ;
        RECT 1748.150 2800.000 1748.610 2801.750 ;
        RECT 1753.370 2800.050 1753.670 2804.600 ;
        RECT 1747.390 2794.625 1747.690 2800.000 ;
        RECT 1747.375 2794.295 1747.705 2794.625 ;
        RECT 1748.310 2787.825 1748.610 2800.000 ;
        RECT 1752.910 2799.750 1753.670 2800.050 ;
        RECT 1753.990 2801.750 1754.290 2804.600 ;
        RECT 1753.990 2801.450 1755.050 2801.750 ;
        RECT 1753.990 2800.000 1754.290 2801.450 ;
        RECT 1752.910 2792.585 1753.210 2799.750 ;
        RECT 1752.895 2792.255 1753.225 2792.585 ;
        RECT 1754.750 2787.825 1755.050 2801.450 ;
        RECT 1759.210 2795.970 1759.510 2804.600 ;
        RECT 1759.830 2796.650 1760.130 2804.600 ;
        RECT 1765.050 2801.750 1765.350 2804.600 ;
        RECT 1762.110 2801.450 1765.350 2801.750 ;
        RECT 1759.830 2796.350 1760.570 2796.650 ;
        RECT 1759.210 2795.670 1759.650 2795.970 ;
        RECT 1759.350 2791.905 1759.650 2795.670 ;
        RECT 1759.335 2791.575 1759.665 2791.905 ;
        RECT 1760.270 2787.825 1760.570 2796.350 ;
        RECT 1762.110 2794.625 1762.410 2801.450 ;
        RECT 1765.050 2800.000 1765.350 2801.450 ;
        RECT 1765.670 2801.750 1765.970 2804.600 ;
        RECT 1770.890 2801.750 1771.190 2804.600 ;
        RECT 1765.670 2800.000 1766.090 2801.750 ;
        RECT 1762.095 2794.295 1762.425 2794.625 ;
        RECT 1765.790 2788.505 1766.090 2800.000 ;
        RECT 1767.630 2801.450 1771.190 2801.750 ;
        RECT 1767.630 2793.945 1767.930 2801.450 ;
        RECT 1770.890 2800.000 1771.190 2801.450 ;
        RECT 1771.510 2801.750 1771.810 2804.600 ;
        RECT 1776.730 2801.750 1777.030 2804.600 ;
        RECT 1771.510 2801.450 1772.530 2801.750 ;
        RECT 1771.510 2800.000 1771.810 2801.450 ;
        RECT 1767.615 2793.615 1767.945 2793.945 ;
        RECT 1765.775 2788.175 1766.105 2788.505 ;
        RECT 1772.230 2787.825 1772.530 2801.450 ;
        RECT 1774.070 2801.450 1777.030 2801.750 ;
        RECT 1774.070 2791.905 1774.370 2801.450 ;
        RECT 1776.730 2800.000 1777.030 2801.450 ;
        RECT 1777.350 2800.050 1777.650 2804.600 ;
        RECT 1782.570 2801.750 1782.870 2804.600 ;
        RECT 1780.510 2801.450 1782.870 2801.750 ;
        RECT 1777.350 2799.750 1778.050 2800.050 ;
        RECT 1774.055 2791.575 1774.385 2791.905 ;
        RECT 1777.750 2787.825 1778.050 2799.750 ;
        RECT 1780.510 2793.945 1780.810 2801.450 ;
        RECT 1782.570 2800.000 1782.870 2801.450 ;
        RECT 1783.190 2801.750 1783.490 2804.600 ;
        RECT 1783.190 2800.000 1783.570 2801.750 ;
        RECT 1788.410 2800.050 1788.710 2804.600 ;
        RECT 1780.495 2793.615 1780.825 2793.945 ;
        RECT 1783.270 2787.825 1783.570 2800.000 ;
        RECT 1787.870 2799.750 1788.710 2800.050 ;
        RECT 1789.030 2801.750 1789.330 2804.600 ;
        RECT 1789.030 2801.450 1790.010 2801.750 ;
        RECT 1789.030 2800.000 1789.330 2801.450 ;
        RECT 1787.870 2793.265 1788.170 2799.750 ;
        RECT 1787.855 2792.935 1788.185 2793.265 ;
        RECT 1789.710 2787.825 1790.010 2801.450 ;
        RECT 1794.250 2796.650 1794.550 2804.600 ;
        RECT 1794.870 2799.385 1795.170 2804.600 ;
        RECT 2234.010 2801.750 2234.310 2804.600 ;
        RECT 2239.850 2801.750 2240.150 2804.600 ;
        RECT 2245.690 2801.750 2245.990 2804.600 ;
        RECT 2251.530 2801.750 2251.830 2804.600 ;
        RECT 2257.370 2801.750 2257.670 2804.600 ;
        RECT 2231.310 2801.450 2234.310 2801.750 ;
        RECT 1794.855 2799.055 1795.185 2799.385 ;
        RECT 1795.215 2797.695 1795.545 2798.025 ;
        RECT 1794.250 2796.350 1794.610 2796.650 ;
        RECT 1794.310 2791.905 1794.610 2796.350 ;
        RECT 1794.295 2791.575 1794.625 2791.905 ;
        RECT 1795.230 2787.825 1795.530 2797.695 ;
        RECT 2231.310 2787.825 2231.610 2801.450 ;
        RECT 2234.010 2800.000 2234.310 2801.450 ;
        RECT 2236.830 2801.450 2240.150 2801.750 ;
        RECT 2236.830 2789.185 2237.130 2801.450 ;
        RECT 2239.850 2800.000 2240.150 2801.450 ;
        RECT 2243.270 2801.450 2245.990 2801.750 ;
        RECT 2243.270 2794.625 2243.570 2801.450 ;
        RECT 2245.690 2800.000 2245.990 2801.450 ;
        RECT 2249.710 2801.450 2251.830 2801.750 ;
        RECT 2243.255 2794.295 2243.585 2794.625 ;
        RECT 2249.710 2791.225 2250.010 2801.450 ;
        RECT 2251.530 2800.000 2251.830 2801.450 ;
        RECT 2257.070 2800.000 2257.670 2801.750 ;
        RECT 2257.070 2794.625 2257.370 2800.000 ;
        RECT 2263.210 2796.650 2263.510 2804.600 ;
        RECT 2263.830 2801.750 2264.130 2804.600 ;
        RECT 2269.050 2801.750 2269.350 2804.600 ;
        RECT 2263.830 2801.450 2264.730 2801.750 ;
        RECT 2263.830 2800.000 2264.130 2801.450 ;
        RECT 2263.210 2796.350 2263.810 2796.650 ;
        RECT 2257.055 2794.295 2257.385 2794.625 ;
        RECT 2263.510 2793.265 2263.810 2796.350 ;
        RECT 2264.430 2794.625 2264.730 2801.450 ;
        RECT 2268.110 2801.450 2269.350 2801.750 ;
        RECT 2268.110 2794.625 2268.410 2801.450 ;
        RECT 2269.050 2800.000 2269.350 2801.450 ;
        RECT 2269.670 2796.650 2269.970 2804.600 ;
        RECT 2274.890 2802.450 2275.190 2804.600 ;
        RECT 2269.030 2796.350 2269.970 2796.650 ;
        RECT 2273.630 2802.150 2275.190 2802.450 ;
        RECT 2264.415 2794.295 2264.745 2794.625 ;
        RECT 2268.095 2794.295 2268.425 2794.625 ;
        RECT 2269.030 2793.945 2269.330 2796.350 ;
        RECT 2273.630 2793.945 2273.930 2802.150 ;
        RECT 2274.890 2800.000 2275.190 2802.150 ;
        RECT 2275.510 2801.750 2275.810 2804.600 ;
        RECT 2280.730 2801.750 2281.030 2804.600 ;
        RECT 2275.510 2801.450 2276.690 2801.750 ;
        RECT 2275.510 2800.000 2275.810 2801.450 ;
        RECT 2276.390 2794.625 2276.690 2801.450 ;
        RECT 2280.070 2801.450 2281.030 2801.750 ;
        RECT 2276.375 2794.295 2276.705 2794.625 ;
        RECT 2280.070 2793.945 2280.370 2801.450 ;
        RECT 2280.730 2800.000 2281.030 2801.450 ;
        RECT 2281.350 2802.450 2281.650 2804.600 ;
        RECT 2281.350 2802.150 2283.130 2802.450 ;
        RECT 2281.350 2800.000 2281.650 2802.150 ;
        RECT 2282.830 2794.625 2283.130 2802.150 ;
        RECT 2286.570 2801.750 2286.870 2804.600 ;
        RECT 2284.670 2801.450 2286.870 2801.750 ;
        RECT 2282.815 2794.295 2283.145 2794.625 ;
        RECT 2284.670 2793.945 2284.970 2801.450 ;
        RECT 2286.570 2800.000 2286.870 2801.450 ;
        RECT 2287.190 2801.750 2287.490 2804.600 ;
        RECT 2287.190 2800.000 2287.730 2801.750 ;
        RECT 2292.410 2800.050 2292.710 2804.600 ;
        RECT 2287.430 2794.625 2287.730 2800.000 ;
        RECT 2292.030 2799.750 2292.710 2800.050 ;
        RECT 2293.030 2801.750 2293.330 2804.600 ;
        RECT 2298.250 2801.750 2298.550 2804.600 ;
        RECT 2293.030 2801.450 2294.170 2801.750 ;
        RECT 2293.030 2800.000 2293.330 2801.450 ;
        RECT 2287.415 2794.295 2287.745 2794.625 ;
        RECT 2269.015 2793.615 2269.345 2793.945 ;
        RECT 2273.615 2793.615 2273.945 2793.945 ;
        RECT 2280.055 2793.615 2280.385 2793.945 ;
        RECT 2284.655 2793.615 2284.985 2793.945 ;
        RECT 2292.030 2793.265 2292.330 2799.750 ;
        RECT 2293.870 2794.625 2294.170 2801.450 ;
        RECT 2297.550 2801.450 2298.550 2801.750 ;
        RECT 2293.855 2794.295 2294.185 2794.625 ;
        RECT 2297.550 2793.945 2297.850 2801.450 ;
        RECT 2298.250 2800.000 2298.550 2801.450 ;
        RECT 2298.870 2802.450 2299.170 2804.600 ;
        RECT 2298.870 2802.150 2300.610 2802.450 ;
        RECT 2298.870 2800.000 2299.170 2802.150 ;
        RECT 2300.310 2794.625 2300.610 2802.150 ;
        RECT 2304.090 2801.750 2304.390 2804.600 ;
        RECT 2303.990 2800.000 2304.390 2801.750 ;
        RECT 2304.710 2801.750 2305.010 2804.600 ;
        RECT 2309.930 2802.450 2310.230 2804.600 ;
        RECT 2308.590 2802.150 2310.230 2802.450 ;
        RECT 2304.710 2800.000 2305.210 2801.750 ;
        RECT 2300.295 2794.295 2300.625 2794.625 ;
        RECT 2303.990 2793.945 2304.290 2800.000 ;
        RECT 2304.910 2794.625 2305.210 2800.000 ;
        RECT 2308.590 2794.625 2308.890 2802.150 ;
        RECT 2309.930 2800.000 2310.230 2802.150 ;
        RECT 2310.550 2796.650 2310.850 2804.600 ;
        RECT 2315.770 2801.750 2316.070 2804.600 ;
        RECT 2310.430 2796.350 2310.850 2796.650 ;
        RECT 2315.030 2801.450 2316.070 2801.750 ;
        RECT 2304.895 2794.295 2305.225 2794.625 ;
        RECT 2308.575 2794.295 2308.905 2794.625 ;
        RECT 2310.430 2793.945 2310.730 2796.350 ;
        RECT 2315.030 2793.945 2315.330 2801.450 ;
        RECT 2315.770 2800.000 2316.070 2801.450 ;
        RECT 2316.390 2800.050 2316.690 2804.600 ;
        RECT 2321.610 2801.750 2321.910 2804.600 ;
        RECT 2316.390 2799.750 2317.170 2800.050 ;
        RECT 2316.870 2794.625 2317.170 2799.750 ;
        RECT 2321.470 2800.000 2321.910 2801.750 ;
        RECT 2322.230 2801.750 2322.530 2804.600 ;
        RECT 2327.450 2802.450 2327.750 2804.600 ;
        RECT 2326.070 2802.150 2327.750 2802.450 ;
        RECT 2322.230 2800.000 2322.690 2801.750 ;
        RECT 2316.855 2794.295 2317.185 2794.625 ;
        RECT 2321.470 2793.945 2321.770 2800.000 ;
        RECT 2322.390 2794.625 2322.690 2800.000 ;
        RECT 2322.375 2794.295 2322.705 2794.625 ;
        RECT 2326.070 2793.945 2326.370 2802.150 ;
        RECT 2327.450 2800.000 2327.750 2802.150 ;
        RECT 2328.070 2801.750 2328.370 2804.600 ;
        RECT 2333.290 2801.750 2333.590 2804.600 ;
        RECT 2328.070 2801.450 2329.130 2801.750 ;
        RECT 2328.070 2800.000 2328.370 2801.450 ;
        RECT 2328.830 2794.625 2329.130 2801.450 ;
        RECT 2332.510 2801.450 2333.590 2801.750 ;
        RECT 2328.815 2794.295 2329.145 2794.625 ;
        RECT 2332.510 2793.945 2332.810 2801.450 ;
        RECT 2333.290 2800.000 2333.590 2801.450 ;
        RECT 2333.910 2800.050 2334.210 2804.600 ;
        RECT 2339.130 2801.750 2339.430 2804.600 ;
        RECT 2333.910 2799.750 2334.650 2800.050 ;
        RECT 2334.350 2794.625 2334.650 2799.750 ;
        RECT 2338.950 2800.000 2339.430 2801.750 ;
        RECT 2339.750 2801.750 2340.050 2804.600 ;
        RECT 2344.970 2802.450 2345.270 2804.600 ;
        RECT 2343.550 2802.150 2345.270 2802.450 ;
        RECT 2339.750 2800.000 2340.170 2801.750 ;
        RECT 2334.335 2794.295 2334.665 2794.625 ;
        RECT 2297.535 2793.615 2297.865 2793.945 ;
        RECT 2303.975 2793.615 2304.305 2793.945 ;
        RECT 2310.415 2793.615 2310.745 2793.945 ;
        RECT 2315.015 2793.615 2315.345 2793.945 ;
        RECT 2321.455 2793.615 2321.785 2793.945 ;
        RECT 2326.055 2793.615 2326.385 2793.945 ;
        RECT 2332.495 2793.615 2332.825 2793.945 ;
        RECT 2338.950 2793.265 2339.250 2800.000 ;
        RECT 2339.870 2794.625 2340.170 2800.000 ;
        RECT 2343.550 2794.625 2343.850 2802.150 ;
        RECT 2344.970 2800.000 2345.270 2802.150 ;
        RECT 2345.590 2796.650 2345.890 2804.600 ;
        RECT 2350.810 2801.750 2351.110 2804.600 ;
        RECT 2345.390 2796.350 2345.890 2796.650 ;
        RECT 2348.150 2801.450 2351.110 2801.750 ;
        RECT 2339.855 2794.295 2340.185 2794.625 ;
        RECT 2343.535 2794.295 2343.865 2794.625 ;
        RECT 2345.390 2793.945 2345.690 2796.350 ;
        RECT 2348.150 2793.945 2348.450 2801.450 ;
        RECT 2350.810 2800.000 2351.110 2801.450 ;
        RECT 2351.430 2800.050 2351.730 2804.600 ;
        RECT 2356.650 2801.750 2356.950 2804.600 ;
        RECT 2351.430 2799.750 2352.130 2800.050 ;
        RECT 2351.830 2794.625 2352.130 2799.750 ;
        RECT 2356.430 2800.000 2356.950 2801.750 ;
        RECT 2357.270 2801.750 2357.570 2804.600 ;
        RECT 2362.490 2802.450 2362.790 2804.600 ;
        RECT 2361.030 2802.150 2362.790 2802.450 ;
        RECT 2357.270 2800.000 2357.650 2801.750 ;
        RECT 2351.815 2794.295 2352.145 2794.625 ;
        RECT 2356.430 2793.945 2356.730 2800.000 ;
        RECT 2357.350 2794.625 2357.650 2800.000 ;
        RECT 2357.335 2794.295 2357.665 2794.625 ;
        RECT 2361.030 2793.945 2361.330 2802.150 ;
        RECT 2362.490 2800.000 2362.790 2802.150 ;
        RECT 2363.110 2801.750 2363.410 2804.600 ;
        RECT 2368.330 2801.750 2368.630 2804.600 ;
        RECT 2363.110 2801.450 2364.090 2801.750 ;
        RECT 2363.110 2800.000 2363.410 2801.450 ;
        RECT 2363.790 2794.625 2364.090 2801.450 ;
        RECT 2367.470 2801.450 2368.630 2801.750 ;
        RECT 2363.775 2794.295 2364.105 2794.625 ;
        RECT 2367.470 2793.945 2367.770 2801.450 ;
        RECT 2368.330 2800.000 2368.630 2801.450 ;
        RECT 2368.950 2802.450 2369.250 2804.600 ;
        RECT 2368.950 2802.150 2370.530 2802.450 ;
        RECT 2368.950 2800.000 2369.250 2802.150 ;
        RECT 2370.230 2794.625 2370.530 2802.150 ;
        RECT 2374.170 2801.750 2374.470 2804.600 ;
        RECT 2373.910 2800.000 2374.470 2801.750 ;
        RECT 2374.790 2801.750 2375.090 2804.600 ;
        RECT 2380.010 2801.750 2380.310 2804.600 ;
        RECT 2374.790 2800.000 2375.130 2801.750 ;
        RECT 2373.910 2794.625 2374.210 2800.000 ;
        RECT 2370.215 2794.295 2370.545 2794.625 ;
        RECT 2373.895 2794.295 2374.225 2794.625 ;
        RECT 2345.375 2793.615 2345.705 2793.945 ;
        RECT 2348.135 2793.615 2348.465 2793.945 ;
        RECT 2356.415 2793.615 2356.745 2793.945 ;
        RECT 2361.015 2793.615 2361.345 2793.945 ;
        RECT 2367.455 2793.615 2367.785 2793.945 ;
        RECT 2374.830 2793.265 2375.130 2800.000 ;
        RECT 2377.590 2801.450 2380.310 2801.750 ;
        RECT 2377.590 2793.945 2377.890 2801.450 ;
        RECT 2380.010 2800.000 2380.310 2801.450 ;
        RECT 2380.630 2801.750 2380.930 2804.600 ;
        RECT 2380.630 2801.450 2381.570 2801.750 ;
        RECT 2380.630 2800.000 2380.930 2801.450 ;
        RECT 2377.575 2793.615 2377.905 2793.945 ;
        RECT 2263.495 2792.935 2263.825 2793.265 ;
        RECT 2292.015 2792.935 2292.345 2793.265 ;
        RECT 2338.935 2792.935 2339.265 2793.265 ;
        RECT 2374.815 2792.935 2375.145 2793.265 ;
        RECT 2249.695 2790.895 2250.025 2791.225 ;
        RECT 2381.270 2789.865 2381.570 2801.450 ;
        RECT 2385.850 2800.050 2386.150 2804.600 ;
        RECT 2386.470 2800.050 2386.770 2804.600 ;
        RECT 2391.690 2801.750 2391.990 2804.600 ;
        RECT 2385.850 2799.750 2386.170 2800.050 ;
        RECT 2386.470 2799.750 2387.090 2800.050 ;
        RECT 2385.870 2794.625 2386.170 2799.750 ;
        RECT 2385.855 2794.295 2386.185 2794.625 ;
        RECT 2386.790 2790.545 2387.090 2799.750 ;
        RECT 2391.390 2800.000 2391.990 2801.750 ;
        RECT 2391.390 2794.625 2391.690 2800.000 ;
        RECT 2391.375 2794.295 2391.705 2794.625 ;
        RECT 2392.310 2791.905 2392.610 2804.600 ;
        RECT 2397.530 2801.750 2397.830 2804.600 ;
        RECT 2395.070 2801.450 2397.830 2801.750 ;
        RECT 2395.070 2794.625 2395.370 2801.450 ;
        RECT 2397.530 2800.000 2397.830 2801.450 ;
        RECT 2398.150 2801.750 2398.450 2804.600 ;
        RECT 2403.370 2801.750 2403.670 2804.600 ;
        RECT 2398.150 2801.450 2399.050 2801.750 ;
        RECT 2398.150 2800.000 2398.450 2801.450 ;
        RECT 2395.055 2794.295 2395.385 2794.625 ;
        RECT 2392.295 2791.575 2392.625 2791.905 ;
        RECT 2398.750 2790.545 2399.050 2801.450 ;
        RECT 2403.350 2800.000 2403.670 2801.750 ;
        RECT 2403.990 2801.750 2404.290 2804.600 ;
        RECT 2409.210 2802.450 2409.510 2804.600 ;
        RECT 2407.950 2802.150 2409.510 2802.450 ;
        RECT 2403.990 2800.000 2404.570 2801.750 ;
        RECT 2403.350 2793.945 2403.650 2800.000 ;
        RECT 2403.335 2793.615 2403.665 2793.945 ;
        RECT 2404.270 2793.265 2404.570 2800.000 ;
        RECT 2407.950 2793.265 2408.250 2802.150 ;
        RECT 2409.210 2800.000 2409.510 2802.150 ;
        RECT 2409.830 2801.750 2410.130 2804.600 ;
        RECT 2409.830 2801.450 2411.010 2801.750 ;
        RECT 2409.830 2800.000 2410.130 2801.450 ;
        RECT 2404.255 2792.935 2404.585 2793.265 ;
        RECT 2407.935 2792.935 2408.265 2793.265 ;
        RECT 2410.710 2791.225 2411.010 2801.450 ;
        RECT 2415.050 2796.650 2415.350 2804.600 ;
        RECT 2415.670 2802.450 2415.970 2804.600 ;
        RECT 2415.670 2802.150 2417.450 2802.450 ;
        RECT 2415.670 2800.000 2415.970 2802.150 ;
        RECT 2415.050 2796.350 2415.610 2796.650 ;
        RECT 2415.310 2793.265 2415.610 2796.350 ;
        RECT 2415.295 2792.935 2415.625 2793.265 ;
        RECT 2410.695 2790.895 2411.025 2791.225 ;
        RECT 2386.775 2790.215 2387.105 2790.545 ;
        RECT 2398.735 2790.215 2399.065 2790.545 ;
        RECT 2381.255 2789.535 2381.585 2789.865 ;
        RECT 2417.150 2789.185 2417.450 2802.150 ;
        RECT 2420.890 2801.750 2421.190 2804.600 ;
        RECT 2418.070 2801.450 2421.190 2801.750 ;
        RECT 2418.070 2792.585 2418.370 2801.450 ;
        RECT 2420.890 2800.000 2421.190 2801.450 ;
        RECT 2421.510 2796.650 2421.810 2804.600 ;
        RECT 2426.730 2801.750 2427.030 2804.600 ;
        RECT 2420.830 2796.350 2421.810 2796.650 ;
        RECT 2423.590 2801.450 2427.030 2801.750 ;
        RECT 2420.830 2794.625 2421.130 2796.350 ;
        RECT 2420.815 2794.295 2421.145 2794.625 ;
        RECT 2423.590 2793.945 2423.890 2801.450 ;
        RECT 2426.730 2800.000 2427.030 2801.450 ;
        RECT 2427.350 2801.750 2427.650 2804.600 ;
        RECT 2432.570 2801.750 2432.870 2804.600 ;
        RECT 2427.350 2801.450 2428.490 2801.750 ;
        RECT 2427.350 2800.000 2427.650 2801.450 ;
        RECT 2423.575 2793.615 2423.905 2793.945 ;
        RECT 2418.055 2792.255 2418.385 2792.585 ;
        RECT 2236.815 2788.855 2237.145 2789.185 ;
        RECT 2417.135 2788.855 2417.465 2789.185 ;
        RECT 2428.190 2788.505 2428.490 2801.450 ;
        RECT 2430.030 2801.450 2432.870 2801.750 ;
        RECT 2430.030 2794.625 2430.330 2801.450 ;
        RECT 2432.570 2800.000 2432.870 2801.450 ;
        RECT 2433.190 2800.050 2433.490 2804.600 ;
        RECT 2438.410 2801.750 2438.710 2804.600 ;
        RECT 2436.470 2801.450 2438.710 2801.750 ;
        RECT 2433.190 2799.750 2434.010 2800.050 ;
        RECT 2430.015 2794.295 2430.345 2794.625 ;
        RECT 2433.710 2791.905 2434.010 2799.750 ;
        RECT 2436.470 2793.945 2436.770 2801.450 ;
        RECT 2438.410 2800.000 2438.710 2801.450 ;
        RECT 2439.030 2801.750 2439.330 2804.600 ;
        RECT 2444.250 2801.750 2444.550 2804.600 ;
        RECT 2439.030 2800.000 2439.530 2801.750 ;
        RECT 2436.455 2793.615 2436.785 2793.945 ;
        RECT 2439.230 2791.905 2439.530 2800.000 ;
        RECT 2442.910 2801.450 2444.550 2801.750 ;
        RECT 2442.910 2793.265 2443.210 2801.450 ;
        RECT 2444.250 2800.000 2444.550 2801.450 ;
        RECT 2444.870 2801.750 2445.170 2804.600 ;
        RECT 2444.870 2801.450 2445.970 2801.750 ;
        RECT 2444.870 2800.000 2445.170 2801.450 ;
        RECT 2442.895 2792.935 2443.225 2793.265 ;
        RECT 2433.695 2791.575 2434.025 2791.905 ;
        RECT 2439.215 2791.575 2439.545 2791.905 ;
        RECT 2445.670 2790.545 2445.970 2801.450 ;
        RECT 2445.655 2790.215 2445.985 2790.545 ;
        RECT 2428.175 2788.175 2428.505 2788.505 ;
        RECT 1580.855 2787.495 1581.185 2787.825 ;
        RECT 1594.655 2787.495 1594.985 2787.825 ;
        RECT 1604.775 2787.495 1605.105 2787.825 ;
        RECT 1613.975 2787.495 1614.305 2787.825 ;
        RECT 1620.415 2787.495 1620.745 2787.825 ;
        RECT 1626.855 2787.495 1627.185 2787.825 ;
        RECT 1630.535 2787.495 1630.865 2787.825 ;
        RECT 1648.935 2787.495 1649.265 2787.825 ;
        RECT 1660.895 2787.495 1661.225 2787.825 ;
        RECT 1666.415 2787.495 1666.745 2787.825 ;
        RECT 1672.855 2787.495 1673.185 2787.825 ;
        RECT 1678.375 2787.495 1678.705 2787.825 ;
        RECT 1683.895 2787.495 1684.225 2787.825 ;
        RECT 1695.855 2787.495 1696.185 2787.825 ;
        RECT 1702.295 2787.495 1702.625 2787.825 ;
        RECT 1708.735 2787.495 1709.065 2787.825 ;
        RECT 1713.335 2787.495 1713.665 2787.825 ;
        RECT 1719.775 2787.495 1720.105 2787.825 ;
        RECT 1730.815 2787.495 1731.145 2787.825 ;
        RECT 1737.255 2787.495 1737.585 2787.825 ;
        RECT 1743.695 2787.495 1744.025 2787.825 ;
        RECT 1748.295 2787.495 1748.625 2787.825 ;
        RECT 1754.735 2787.495 1755.065 2787.825 ;
        RECT 1760.255 2787.495 1760.585 2787.825 ;
        RECT 1772.215 2787.495 1772.545 2787.825 ;
        RECT 1777.735 2787.495 1778.065 2787.825 ;
        RECT 1783.255 2787.495 1783.585 2787.825 ;
        RECT 1789.695 2787.495 1790.025 2787.825 ;
        RECT 1795.215 2787.495 1795.545 2787.825 ;
        RECT 2231.295 2787.495 2231.625 2787.825 ;
        RECT 1691.310 2051.635 1691.610 2056.235 ;
        RECT 1691.930 2051.635 1692.230 2056.235 ;
        RECT 1697.150 2051.635 1697.450 2056.235 ;
        RECT 1697.770 2051.635 1698.070 2056.235 ;
        RECT 1702.990 2051.635 1703.290 2056.235 ;
        RECT 1703.610 2051.635 1703.910 2056.235 ;
        RECT 1708.830 2051.635 1709.130 2056.235 ;
        RECT 1709.450 2051.635 1709.750 2056.235 ;
        RECT 1714.670 2051.635 1714.970 2056.235 ;
        RECT 1715.290 2051.635 1715.590 2056.235 ;
        RECT 1720.510 2051.635 1720.810 2056.235 ;
        RECT 1721.130 2051.635 1721.430 2056.235 ;
        RECT 1726.350 2051.635 1726.650 2056.235 ;
        RECT 1726.970 2051.635 1727.270 2056.235 ;
        RECT 1732.190 2051.635 1732.490 2056.235 ;
        RECT 1732.810 2051.635 1733.110 2056.235 ;
        RECT 1738.030 2051.635 1738.330 2056.235 ;
        RECT 1738.650 2051.635 1738.950 2056.235 ;
        RECT 1743.870 2051.635 1744.170 2056.235 ;
        RECT 1744.490 2051.635 1744.790 2056.235 ;
        RECT 1749.710 2051.635 1750.010 2056.235 ;
        RECT 1750.330 2051.635 1750.630 2056.235 ;
        RECT 1755.550 2051.635 1755.850 2056.235 ;
        RECT 1756.170 2051.635 1756.470 2056.235 ;
        RECT 1761.390 2051.635 1761.690 2056.235 ;
        RECT 1762.010 2051.635 1762.310 2056.235 ;
        RECT 1767.230 2051.635 1767.530 2056.235 ;
        RECT 1767.850 2051.635 1768.150 2056.235 ;
        RECT 1773.070 2051.635 1773.370 2056.235 ;
        RECT 1773.690 2051.635 1773.990 2056.235 ;
        RECT 1778.910 2051.635 1779.210 2056.235 ;
        RECT 1779.530 2051.635 1779.830 2056.235 ;
        RECT 1784.750 2051.635 1785.050 2056.235 ;
        RECT 1785.370 2051.635 1785.670 2056.235 ;
        RECT 1790.590 2051.635 1790.890 2056.235 ;
        RECT 1791.210 2051.635 1791.510 2056.235 ;
        RECT 1796.430 2051.635 1796.730 2056.235 ;
        RECT 1797.050 2051.635 1797.350 2056.235 ;
        RECT 1802.270 2051.635 1802.570 2056.235 ;
        RECT 1802.890 2051.635 1803.190 2056.235 ;
        RECT 1808.110 2051.635 1808.410 2056.235 ;
        RECT 1808.730 2051.635 1809.030 2056.235 ;
        RECT 1813.950 2051.635 1814.250 2056.235 ;
        RECT 1814.570 2051.635 1814.870 2056.235 ;
        RECT 1819.790 2051.635 1820.090 2056.235 ;
        RECT 1820.410 2051.635 1820.710 2056.235 ;
        RECT 1825.630 2051.635 1825.930 2056.235 ;
        RECT 1826.250 2051.635 1826.550 2056.235 ;
        RECT 1831.470 2051.635 1831.770 2056.235 ;
        RECT 1832.090 2051.635 1832.390 2056.235 ;
        RECT 1837.310 2051.635 1837.610 2056.235 ;
        RECT 1837.930 2051.635 1838.230 2056.235 ;
        RECT 1843.150 2051.635 1843.450 2056.235 ;
        RECT 1843.770 2051.635 1844.070 2056.235 ;
        RECT 1848.990 2051.635 1849.290 2056.235 ;
        RECT 1849.610 2051.635 1849.910 2056.235 ;
        RECT 1854.830 2051.635 1855.130 2056.235 ;
        RECT 1855.450 2051.635 1855.750 2056.235 ;
        RECT 1860.670 2051.635 1860.970 2056.235 ;
        RECT 1861.290 2051.635 1861.590 2056.235 ;
        RECT 1866.510 2051.635 1866.810 2056.235 ;
        RECT 1867.130 2051.635 1867.430 2056.235 ;
        RECT 1872.350 2051.635 1872.650 2056.235 ;
        RECT 1872.970 2051.635 1873.270 2056.235 ;
        RECT 1878.810 2051.635 1879.110 2056.235 ;
        RECT 1884.650 2051.635 1884.950 2056.235 ;
        RECT 1890.490 2051.635 1890.790 2056.235 ;
        RECT 1896.330 2051.635 1896.630 2056.235 ;
        RECT 1902.170 2051.635 1902.470 2056.235 ;
        RECT 2294.025 2051.635 2294.325 2056.235 ;
        RECT 2300.265 2051.635 2300.565 2056.235 ;
        RECT 2306.505 2051.635 2306.805 2056.235 ;
        RECT 2312.745 2051.635 2313.045 2056.235 ;
        RECT 2318.985 2051.635 2319.285 2056.235 ;
        RECT 2325.225 2051.635 2325.525 2056.235 ;
        RECT 2331.465 2051.635 2331.765 2056.235 ;
        RECT 2337.705 2051.635 2338.005 2056.235 ;
        RECT 2343.945 2051.635 2344.245 2056.235 ;
        RECT 2350.185 2051.635 2350.485 2056.235 ;
        RECT 2356.425 2051.635 2356.725 2056.235 ;
        RECT 2362.665 2051.635 2362.965 2056.235 ;
        RECT 2368.905 2051.635 2369.205 2056.235 ;
        RECT 2375.145 2051.635 2375.445 2056.235 ;
        RECT 2381.385 2051.635 2381.685 2056.235 ;
        RECT 2387.625 2051.635 2387.925 2056.235 ;
        RECT 2393.865 2051.635 2394.165 2056.235 ;
        RECT 2400.105 2051.635 2400.405 2056.235 ;
        RECT 2406.345 2051.635 2406.645 2056.235 ;
        RECT 2412.585 2051.635 2412.885 2056.235 ;
        RECT 2418.825 2051.635 2419.125 2056.235 ;
        RECT 2425.065 2051.635 2425.365 2056.235 ;
        RECT 2431.305 2051.635 2431.605 2056.235 ;
        RECT 2437.545 2051.635 2437.845 2056.235 ;
        RECT 2443.785 2051.635 2444.085 2056.235 ;
        RECT 2450.025 2051.635 2450.325 2056.235 ;
        RECT 2456.265 2051.635 2456.565 2056.235 ;
        RECT 2462.505 2051.635 2462.805 2056.235 ;
        RECT 2468.745 2051.635 2469.045 2056.235 ;
        RECT 2474.985 2051.635 2475.285 2056.235 ;
        RECT 2481.225 2051.635 2481.525 2056.235 ;
        RECT 2487.465 2051.635 2487.765 2056.235 ;
        RECT 2542.890 2051.635 2543.190 2056.235 ;
        RECT 1417.095 1627.415 1417.425 1627.745 ;
      LAYER met4 ;
        RECT 1555.000 1605.000 1931.480 2051.235 ;
        RECT 2205.000 1605.000 2581.480 2051.235 ;
      LAYER met4 ;
        RECT 1593.290 1600.000 1593.590 1604.600 ;
        RECT 1648.715 1600.000 1649.015 1604.600 ;
        RECT 1654.955 1600.000 1655.255 1604.600 ;
        RECT 1661.195 1600.000 1661.495 1604.600 ;
        RECT 1667.435 1600.000 1667.735 1604.600 ;
        RECT 1673.675 1600.000 1673.975 1604.600 ;
        RECT 1679.915 1600.000 1680.215 1604.600 ;
        RECT 1686.155 1600.000 1686.455 1604.600 ;
        RECT 1692.395 1600.000 1692.695 1604.600 ;
        RECT 1698.635 1600.000 1698.935 1604.600 ;
        RECT 1704.875 1600.000 1705.175 1604.600 ;
        RECT 1711.115 1600.000 1711.415 1604.600 ;
        RECT 1717.355 1600.000 1717.655 1604.600 ;
        RECT 1723.595 1600.000 1723.895 1604.600 ;
        RECT 1729.835 1600.000 1730.135 1604.600 ;
        RECT 1736.075 1600.000 1736.375 1604.600 ;
        RECT 1742.315 1600.000 1742.615 1604.600 ;
        RECT 1748.555 1600.000 1748.855 1604.600 ;
        RECT 1754.795 1600.000 1755.095 1604.600 ;
        RECT 1761.035 1600.000 1761.335 1604.600 ;
        RECT 1767.275 1600.000 1767.575 1604.600 ;
        RECT 1773.515 1600.000 1773.815 1604.600 ;
        RECT 1779.755 1600.000 1780.055 1604.600 ;
        RECT 1785.995 1600.000 1786.295 1604.600 ;
        RECT 1792.235 1600.000 1792.535 1604.600 ;
        RECT 1798.475 1600.000 1798.775 1604.600 ;
        RECT 1804.715 1600.000 1805.015 1604.600 ;
        RECT 1810.955 1600.000 1811.255 1604.600 ;
        RECT 1817.195 1600.000 1817.495 1604.600 ;
        RECT 1823.435 1600.000 1823.735 1604.600 ;
        RECT 1829.675 1600.000 1829.975 1604.600 ;
        RECT 1835.915 1600.000 1836.215 1604.600 ;
        RECT 1842.155 1600.000 1842.455 1604.600 ;
        RECT 2234.010 1600.000 2234.310 1604.600 ;
        RECT 2239.850 1600.000 2240.150 1604.600 ;
        RECT 2245.690 1600.000 2245.990 1604.600 ;
        RECT 2251.530 1600.000 2251.830 1604.600 ;
        RECT 2257.370 1600.000 2257.670 1604.600 ;
        RECT 2263.210 1600.000 2263.510 1604.600 ;
        RECT 2263.830 1600.000 2264.130 1604.600 ;
        RECT 2269.050 1600.000 2269.350 1604.600 ;
        RECT 2269.670 1600.000 2269.970 1604.600 ;
        RECT 2274.890 1600.000 2275.190 1604.600 ;
        RECT 2275.510 1600.000 2275.810 1604.600 ;
        RECT 2280.730 1600.000 2281.030 1604.600 ;
        RECT 2281.350 1600.000 2281.650 1604.600 ;
        RECT 2286.570 1600.000 2286.870 1604.600 ;
        RECT 2287.190 1600.000 2287.490 1604.600 ;
        RECT 2292.410 1600.000 2292.710 1604.600 ;
        RECT 2293.030 1600.000 2293.330 1604.600 ;
        RECT 2298.250 1600.000 2298.550 1604.600 ;
        RECT 2298.870 1600.000 2299.170 1604.600 ;
        RECT 2304.090 1600.000 2304.390 1604.600 ;
        RECT 2304.710 1600.000 2305.010 1604.600 ;
        RECT 2309.930 1600.000 2310.230 1604.600 ;
        RECT 2310.550 1600.000 2310.850 1604.600 ;
        RECT 2315.770 1600.000 2316.070 1604.600 ;
        RECT 2316.390 1600.000 2316.690 1604.600 ;
        RECT 2321.610 1600.000 2321.910 1604.600 ;
        RECT 2322.230 1600.000 2322.530 1604.600 ;
        RECT 2327.450 1600.000 2327.750 1604.600 ;
        RECT 2328.070 1600.000 2328.370 1604.600 ;
        RECT 2333.290 1600.000 2333.590 1604.600 ;
        RECT 2333.910 1600.000 2334.210 1604.600 ;
        RECT 2339.130 1600.000 2339.430 1604.600 ;
        RECT 2339.750 1600.000 2340.050 1604.600 ;
        RECT 2344.970 1600.000 2345.270 1604.600 ;
        RECT 2345.590 1600.000 2345.890 1604.600 ;
        RECT 2350.810 1600.000 2351.110 1604.600 ;
        RECT 2351.430 1600.000 2351.730 1604.600 ;
        RECT 2356.650 1600.000 2356.950 1604.600 ;
        RECT 2357.270 1600.000 2357.570 1604.600 ;
        RECT 2362.490 1600.000 2362.790 1604.600 ;
        RECT 2363.110 1600.000 2363.410 1604.600 ;
        RECT 2368.330 1600.000 2368.630 1604.600 ;
        RECT 2368.950 1600.000 2369.250 1604.600 ;
        RECT 2374.170 1600.000 2374.470 1604.600 ;
        RECT 2374.790 1600.000 2375.090 1604.600 ;
        RECT 2380.010 1600.000 2380.310 1604.600 ;
        RECT 2380.630 1600.000 2380.930 1604.600 ;
        RECT 2385.850 1600.000 2386.150 1604.600 ;
        RECT 2386.470 1600.000 2386.770 1604.600 ;
        RECT 2391.690 1600.000 2391.990 1604.600 ;
        RECT 2392.310 1600.000 2392.610 1604.600 ;
        RECT 2397.530 1600.000 2397.830 1604.600 ;
        RECT 2398.150 1600.000 2398.450 1604.600 ;
        RECT 2403.370 1600.000 2403.670 1604.600 ;
        RECT 2403.990 1600.000 2404.290 1604.600 ;
        RECT 2409.210 1600.000 2409.510 1604.600 ;
        RECT 2409.830 1600.000 2410.130 1604.600 ;
        RECT 2415.050 1600.000 2415.350 1604.600 ;
        RECT 2415.670 1600.000 2415.970 1604.600 ;
        RECT 2420.890 1600.000 2421.190 1604.600 ;
        RECT 2421.510 1600.000 2421.810 1604.600 ;
        RECT 2426.730 1600.000 2427.030 1604.600 ;
        RECT 2427.350 1600.000 2427.650 1604.600 ;
        RECT 2432.570 1600.000 2432.870 1604.600 ;
        RECT 2433.190 1600.000 2433.490 1604.600 ;
        RECT 2438.410 1600.000 2438.710 1604.600 ;
        RECT 2439.030 1600.000 2439.330 1604.600 ;
        RECT 2444.250 1600.000 2444.550 1604.600 ;
        RECT 2444.870 1600.000 2445.170 1604.600 ;
        RECT 1588.020 1515.000 1591.020 1585.000 ;
        RECT 1624.020 1515.000 1627.020 1585.000 ;
        RECT 1642.020 1515.000 1645.020 1585.000 ;
        RECT 1660.020 1515.000 1663.020 1585.000 ;
        RECT 1678.020 1515.000 1681.020 1585.000 ;
        RECT 1768.020 1515.000 1771.020 1585.000 ;
        RECT 1804.020 1515.000 1807.020 1585.000 ;
        RECT 1822.020 1515.000 1825.020 1585.000 ;
        RECT 1840.020 1515.000 1843.020 1585.000 ;
        RECT 1858.020 1515.000 1861.020 1585.000 ;
        RECT 1948.020 1515.000 1951.020 1585.000 ;
        RECT 2182.020 1515.000 2185.020 1585.000 ;
        RECT 2200.020 1515.000 2203.020 1585.000 ;
        RECT 2218.020 1515.000 2221.020 1585.000 ;
        RECT 2308.020 1515.000 2311.020 1585.000 ;
        RECT 2344.020 1515.000 2347.020 1585.000 ;
        RECT 2362.020 1515.000 2365.020 1585.000 ;
        RECT 2380.020 1515.000 2383.020 1585.000 ;
        RECT 2398.020 1515.000 2401.020 1585.000 ;
        RECT 2488.020 1515.000 2491.020 1585.000 ;
        RECT 2524.020 1515.000 2527.020 1585.000 ;
        RECT 2542.020 1515.000 2545.020 1585.000 ;
        RECT 2560.020 1515.000 2563.020 1585.000 ;
        RECT 2578.020 1515.000 2581.020 1585.000 ;
      LAYER met4 ;
        RECT 1575.065 410.640 1647.370 1488.240 ;
        RECT 1649.770 410.640 2638.915 1488.240 ;
      LAYER met5 ;
        RECT 1351.140 2935.100 2588.300 2936.700 ;
        RECT 302.340 2894.300 2188.100 2895.900 ;
  END
END user_project_wrapper
END LIBRARY

