VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hs32_core1
  CLASS BLOCK ;
  FOREIGN hs32_core1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 1200.000 ;
  PIN cpu_addr_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 489.640 1100.000 490.240 ;
    END
  END cpu_addr_e[0]
  PIN cpu_addr_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 599.800 1100.000 600.400 ;
    END
  END cpu_addr_e[10]
  PIN cpu_addr_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 610.680 1100.000 611.280 ;
    END
  END cpu_addr_e[11]
  PIN cpu_addr_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 621.560 1100.000 622.160 ;
    END
  END cpu_addr_e[12]
  PIN cpu_addr_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 632.440 1100.000 633.040 ;
    END
  END cpu_addr_e[13]
  PIN cpu_addr_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 644.000 1100.000 644.600 ;
    END
  END cpu_addr_e[14]
  PIN cpu_addr_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 654.880 1100.000 655.480 ;
    END
  END cpu_addr_e[15]
  PIN cpu_addr_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 500.520 1100.000 501.120 ;
    END
  END cpu_addr_e[1]
  PIN cpu_addr_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 511.400 1100.000 512.000 ;
    END
  END cpu_addr_e[2]
  PIN cpu_addr_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 522.960 1100.000 523.560 ;
    END
  END cpu_addr_e[3]
  PIN cpu_addr_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 533.840 1100.000 534.440 ;
    END
  END cpu_addr_e[4]
  PIN cpu_addr_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 544.720 1100.000 545.320 ;
    END
  END cpu_addr_e[5]
  PIN cpu_addr_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 555.600 1100.000 556.200 ;
    END
  END cpu_addr_e[6]
  PIN cpu_addr_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 566.480 1100.000 567.080 ;
    END
  END cpu_addr_e[7]
  PIN cpu_addr_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 578.040 1100.000 578.640 ;
    END
  END cpu_addr_e[8]
  PIN cpu_addr_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 588.920 1100.000 589.520 ;
    END
  END cpu_addr_e[9]
  PIN cpu_addr_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.810 1196.000 337.090 1200.000 ;
    END
  END cpu_addr_n[0]
  PIN cpu_addr_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 440.770 1196.000 441.050 1200.000 ;
    END
  END cpu_addr_n[10]
  PIN cpu_addr_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.890 1196.000 451.170 1200.000 ;
    END
  END cpu_addr_n[11]
  PIN cpu_addr_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 461.470 1196.000 461.750 1200.000 ;
    END
  END cpu_addr_n[12]
  PIN cpu_addr_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.050 1196.000 472.330 1200.000 ;
    END
  END cpu_addr_n[13]
  PIN cpu_addr_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 482.170 1196.000 482.450 1200.000 ;
    END
  END cpu_addr_n[14]
  PIN cpu_addr_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.750 1196.000 493.030 1200.000 ;
    END
  END cpu_addr_n[15]
  PIN cpu_addr_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.390 1196.000 347.670 1200.000 ;
    END
  END cpu_addr_n[1]
  PIN cpu_addr_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.510 1196.000 357.790 1200.000 ;
    END
  END cpu_addr_n[2]
  PIN cpu_addr_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.090 1196.000 368.370 1200.000 ;
    END
  END cpu_addr_n[3]
  PIN cpu_addr_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.670 1196.000 378.950 1200.000 ;
    END
  END cpu_addr_n[4]
  PIN cpu_addr_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.790 1196.000 389.070 1200.000 ;
    END
  END cpu_addr_n[5]
  PIN cpu_addr_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 399.370 1196.000 399.650 1200.000 ;
    END
  END cpu_addr_n[6]
  PIN cpu_addr_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.490 1196.000 409.770 1200.000 ;
    END
  END cpu_addr_n[7]
  PIN cpu_addr_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.070 1196.000 420.350 1200.000 ;
    END
  END cpu_addr_n[8]
  PIN cpu_addr_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.190 1196.000 430.470 1200.000 ;
    END
  END cpu_addr_n[9]
  PIN cpu_dtr_e0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 27.240 1100.000 27.840 ;
    END
  END cpu_dtr_e0[0]
  PIN cpu_dtr_e0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 137.400 1100.000 138.000 ;
    END
  END cpu_dtr_e0[10]
  PIN cpu_dtr_e0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 148.280 1100.000 148.880 ;
    END
  END cpu_dtr_e0[11]
  PIN cpu_dtr_e0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 159.160 1100.000 159.760 ;
    END
  END cpu_dtr_e0[12]
  PIN cpu_dtr_e0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 170.040 1100.000 170.640 ;
    END
  END cpu_dtr_e0[13]
  PIN cpu_dtr_e0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 181.600 1100.000 182.200 ;
    END
  END cpu_dtr_e0[14]
  PIN cpu_dtr_e0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 192.480 1100.000 193.080 ;
    END
  END cpu_dtr_e0[15]
  PIN cpu_dtr_e0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 203.360 1100.000 203.960 ;
    END
  END cpu_dtr_e0[16]
  PIN cpu_dtr_e0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 214.240 1100.000 214.840 ;
    END
  END cpu_dtr_e0[17]
  PIN cpu_dtr_e0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 225.120 1100.000 225.720 ;
    END
  END cpu_dtr_e0[18]
  PIN cpu_dtr_e0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 236.680 1100.000 237.280 ;
    END
  END cpu_dtr_e0[19]
  PIN cpu_dtr_e0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 38.120 1100.000 38.720 ;
    END
  END cpu_dtr_e0[1]
  PIN cpu_dtr_e0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 247.560 1100.000 248.160 ;
    END
  END cpu_dtr_e0[20]
  PIN cpu_dtr_e0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 258.440 1100.000 259.040 ;
    END
  END cpu_dtr_e0[21]
  PIN cpu_dtr_e0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 269.320 1100.000 269.920 ;
    END
  END cpu_dtr_e0[22]
  PIN cpu_dtr_e0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 280.200 1100.000 280.800 ;
    END
  END cpu_dtr_e0[23]
  PIN cpu_dtr_e0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 291.760 1100.000 292.360 ;
    END
  END cpu_dtr_e0[24]
  PIN cpu_dtr_e0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 302.640 1100.000 303.240 ;
    END
  END cpu_dtr_e0[25]
  PIN cpu_dtr_e0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 313.520 1100.000 314.120 ;
    END
  END cpu_dtr_e0[26]
  PIN cpu_dtr_e0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 324.400 1100.000 325.000 ;
    END
  END cpu_dtr_e0[27]
  PIN cpu_dtr_e0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 335.280 1100.000 335.880 ;
    END
  END cpu_dtr_e0[28]
  PIN cpu_dtr_e0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 346.160 1100.000 346.760 ;
    END
  END cpu_dtr_e0[29]
  PIN cpu_dtr_e0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 49.000 1100.000 49.600 ;
    END
  END cpu_dtr_e0[2]
  PIN cpu_dtr_e0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 357.720 1100.000 358.320 ;
    END
  END cpu_dtr_e0[30]
  PIN cpu_dtr_e0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 368.600 1100.000 369.200 ;
    END
  END cpu_dtr_e0[31]
  PIN cpu_dtr_e0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 59.880 1100.000 60.480 ;
    END
  END cpu_dtr_e0[3]
  PIN cpu_dtr_e0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 71.440 1100.000 72.040 ;
    END
  END cpu_dtr_e0[4]
  PIN cpu_dtr_e0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 82.320 1100.000 82.920 ;
    END
  END cpu_dtr_e0[5]
  PIN cpu_dtr_e0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 93.200 1100.000 93.800 ;
    END
  END cpu_dtr_e0[6]
  PIN cpu_dtr_e0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 104.080 1100.000 104.680 ;
    END
  END cpu_dtr_e0[7]
  PIN cpu_dtr_e0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 114.960 1100.000 115.560 ;
    END
  END cpu_dtr_e0[8]
  PIN cpu_dtr_e0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 126.520 1100.000 127.120 ;
    END
  END cpu_dtr_e0[9]
  PIN cpu_dtr_e1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 841.880 1100.000 842.480 ;
    END
  END cpu_dtr_e1[0]
  PIN cpu_dtr_e1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 952.040 1100.000 952.640 ;
    END
  END cpu_dtr_e1[10]
  PIN cpu_dtr_e1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 962.920 1100.000 963.520 ;
    END
  END cpu_dtr_e1[11]
  PIN cpu_dtr_e1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 973.800 1100.000 974.400 ;
    END
  END cpu_dtr_e1[12]
  PIN cpu_dtr_e1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 985.360 1100.000 985.960 ;
    END
  END cpu_dtr_e1[13]
  PIN cpu_dtr_e1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 996.240 1100.000 996.840 ;
    END
  END cpu_dtr_e1[14]
  PIN cpu_dtr_e1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1007.120 1100.000 1007.720 ;
    END
  END cpu_dtr_e1[15]
  PIN cpu_dtr_e1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1018.000 1100.000 1018.600 ;
    END
  END cpu_dtr_e1[16]
  PIN cpu_dtr_e1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1028.880 1100.000 1029.480 ;
    END
  END cpu_dtr_e1[17]
  PIN cpu_dtr_e1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1040.440 1100.000 1041.040 ;
    END
  END cpu_dtr_e1[18]
  PIN cpu_dtr_e1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1051.320 1100.000 1051.920 ;
    END
  END cpu_dtr_e1[19]
  PIN cpu_dtr_e1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 852.760 1100.000 853.360 ;
    END
  END cpu_dtr_e1[1]
  PIN cpu_dtr_e1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1062.200 1100.000 1062.800 ;
    END
  END cpu_dtr_e1[20]
  PIN cpu_dtr_e1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1073.080 1100.000 1073.680 ;
    END
  END cpu_dtr_e1[21]
  PIN cpu_dtr_e1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1083.960 1100.000 1084.560 ;
    END
  END cpu_dtr_e1[22]
  PIN cpu_dtr_e1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1095.520 1100.000 1096.120 ;
    END
  END cpu_dtr_e1[23]
  PIN cpu_dtr_e1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1106.400 1100.000 1107.000 ;
    END
  END cpu_dtr_e1[24]
  PIN cpu_dtr_e1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1117.280 1100.000 1117.880 ;
    END
  END cpu_dtr_e1[25]
  PIN cpu_dtr_e1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1128.160 1100.000 1128.760 ;
    END
  END cpu_dtr_e1[26]
  PIN cpu_dtr_e1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1139.040 1100.000 1139.640 ;
    END
  END cpu_dtr_e1[27]
  PIN cpu_dtr_e1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1150.600 1100.000 1151.200 ;
    END
  END cpu_dtr_e1[28]
  PIN cpu_dtr_e1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1161.480 1100.000 1162.080 ;
    END
  END cpu_dtr_e1[29]
  PIN cpu_dtr_e1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 864.320 1100.000 864.920 ;
    END
  END cpu_dtr_e1[2]
  PIN cpu_dtr_e1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1172.360 1100.000 1172.960 ;
    END
  END cpu_dtr_e1[30]
  PIN cpu_dtr_e1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1183.240 1100.000 1183.840 ;
    END
  END cpu_dtr_e1[31]
  PIN cpu_dtr_e1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 875.200 1100.000 875.800 ;
    END
  END cpu_dtr_e1[3]
  PIN cpu_dtr_e1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 886.080 1100.000 886.680 ;
    END
  END cpu_dtr_e1[4]
  PIN cpu_dtr_e1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 896.960 1100.000 897.560 ;
    END
  END cpu_dtr_e1[5]
  PIN cpu_dtr_e1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 907.840 1100.000 908.440 ;
    END
  END cpu_dtr_e1[6]
  PIN cpu_dtr_e1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 918.720 1100.000 919.320 ;
    END
  END cpu_dtr_e1[7]
  PIN cpu_dtr_e1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 930.280 1100.000 930.880 ;
    END
  END cpu_dtr_e1[8]
  PIN cpu_dtr_e1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 941.160 1100.000 941.760 ;
    END
  END cpu_dtr_e1[9]
  PIN cpu_dtr_n0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 1196.000 5.430 1200.000 ;
    END
  END cpu_dtr_n0[0]
  PIN cpu_dtr_n0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.650 1196.000 108.930 1200.000 ;
    END
  END cpu_dtr_n0[10]
  PIN cpu_dtr_n0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.230 1196.000 119.510 1200.000 ;
    END
  END cpu_dtr_n0[11]
  PIN cpu_dtr_n0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.350 1196.000 129.630 1200.000 ;
    END
  END cpu_dtr_n0[12]
  PIN cpu_dtr_n0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.930 1196.000 140.210 1200.000 ;
    END
  END cpu_dtr_n0[13]
  PIN cpu_dtr_n0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.050 1196.000 150.330 1200.000 ;
    END
  END cpu_dtr_n0[14]
  PIN cpu_dtr_n0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.630 1196.000 160.910 1200.000 ;
    END
  END cpu_dtr_n0[15]
  PIN cpu_dtr_n0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.750 1196.000 171.030 1200.000 ;
    END
  END cpu_dtr_n0[16]
  PIN cpu_dtr_n0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.330 1196.000 181.610 1200.000 ;
    END
  END cpu_dtr_n0[17]
  PIN cpu_dtr_n0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.910 1196.000 192.190 1200.000 ;
    END
  END cpu_dtr_n0[18]
  PIN cpu_dtr_n0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.030 1196.000 202.310 1200.000 ;
    END
  END cpu_dtr_n0[19]
  PIN cpu_dtr_n0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 1196.000 15.550 1200.000 ;
    END
  END cpu_dtr_n0[1]
  PIN cpu_dtr_n0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 212.610 1196.000 212.890 1200.000 ;
    END
  END cpu_dtr_n0[20]
  PIN cpu_dtr_n0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.730 1196.000 223.010 1200.000 ;
    END
  END cpu_dtr_n0[21]
  PIN cpu_dtr_n0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.310 1196.000 233.590 1200.000 ;
    END
  END cpu_dtr_n0[22]
  PIN cpu_dtr_n0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 243.430 1196.000 243.710 1200.000 ;
    END
  END cpu_dtr_n0[23]
  PIN cpu_dtr_n0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.010 1196.000 254.290 1200.000 ;
    END
  END cpu_dtr_n0[24]
  PIN cpu_dtr_n0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.130 1196.000 264.410 1200.000 ;
    END
  END cpu_dtr_n0[25]
  PIN cpu_dtr_n0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.710 1196.000 274.990 1200.000 ;
    END
  END cpu_dtr_n0[26]
  PIN cpu_dtr_n0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 285.290 1196.000 285.570 1200.000 ;
    END
  END cpu_dtr_n0[27]
  PIN cpu_dtr_n0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 295.410 1196.000 295.690 1200.000 ;
    END
  END cpu_dtr_n0[28]
  PIN cpu_dtr_n0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.990 1196.000 306.270 1200.000 ;
    END
  END cpu_dtr_n0[29]
  PIN cpu_dtr_n0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 1196.000 26.130 1200.000 ;
    END
  END cpu_dtr_n0[2]
  PIN cpu_dtr_n0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.110 1196.000 316.390 1200.000 ;
    END
  END cpu_dtr_n0[30]
  PIN cpu_dtr_n0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.690 1196.000 326.970 1200.000 ;
    END
  END cpu_dtr_n0[31]
  PIN cpu_dtr_n0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 1196.000 36.250 1200.000 ;
    END
  END cpu_dtr_n0[3]
  PIN cpu_dtr_n0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 1196.000 46.830 1200.000 ;
    END
  END cpu_dtr_n0[4]
  PIN cpu_dtr_n0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 1196.000 56.950 1200.000 ;
    END
  END cpu_dtr_n0[5]
  PIN cpu_dtr_n0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.250 1196.000 67.530 1200.000 ;
    END
  END cpu_dtr_n0[6]
  PIN cpu_dtr_n0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 1196.000 77.650 1200.000 ;
    END
  END cpu_dtr_n0[7]
  PIN cpu_dtr_n0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.950 1196.000 88.230 1200.000 ;
    END
  END cpu_dtr_n0[8]
  PIN cpu_dtr_n0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.530 1196.000 98.810 1200.000 ;
    END
  END cpu_dtr_n0[9]
  PIN cpu_dtr_n1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 772.890 1196.000 773.170 1200.000 ;
    END
  END cpu_dtr_n1[0]
  PIN cpu_dtr_n1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.390 1196.000 876.670 1200.000 ;
    END
  END cpu_dtr_n1[10]
  PIN cpu_dtr_n1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.970 1196.000 887.250 1200.000 ;
    END
  END cpu_dtr_n1[11]
  PIN cpu_dtr_n1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 897.090 1196.000 897.370 1200.000 ;
    END
  END cpu_dtr_n1[12]
  PIN cpu_dtr_n1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.670 1196.000 907.950 1200.000 ;
    END
  END cpu_dtr_n1[13]
  PIN cpu_dtr_n1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 917.790 1196.000 918.070 1200.000 ;
    END
  END cpu_dtr_n1[14]
  PIN cpu_dtr_n1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 928.370 1196.000 928.650 1200.000 ;
    END
  END cpu_dtr_n1[15]
  PIN cpu_dtr_n1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.950 1196.000 939.230 1200.000 ;
    END
  END cpu_dtr_n1[16]
  PIN cpu_dtr_n1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.070 1196.000 949.350 1200.000 ;
    END
  END cpu_dtr_n1[17]
  PIN cpu_dtr_n1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 959.650 1196.000 959.930 1200.000 ;
    END
  END cpu_dtr_n1[18]
  PIN cpu_dtr_n1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.770 1196.000 970.050 1200.000 ;
    END
  END cpu_dtr_n1[19]
  PIN cpu_dtr_n1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.010 1196.000 783.290 1200.000 ;
    END
  END cpu_dtr_n1[1]
  PIN cpu_dtr_n1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 980.350 1196.000 980.630 1200.000 ;
    END
  END cpu_dtr_n1[20]
  PIN cpu_dtr_n1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 990.470 1196.000 990.750 1200.000 ;
    END
  END cpu_dtr_n1[21]
  PIN cpu_dtr_n1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.050 1196.000 1001.330 1200.000 ;
    END
  END cpu_dtr_n1[22]
  PIN cpu_dtr_n1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1011.170 1196.000 1011.450 1200.000 ;
    END
  END cpu_dtr_n1[23]
  PIN cpu_dtr_n1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1021.750 1196.000 1022.030 1200.000 ;
    END
  END cpu_dtr_n1[24]
  PIN cpu_dtr_n1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.330 1196.000 1032.610 1200.000 ;
    END
  END cpu_dtr_n1[25]
  PIN cpu_dtr_n1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1042.450 1196.000 1042.730 1200.000 ;
    END
  END cpu_dtr_n1[26]
  PIN cpu_dtr_n1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1053.030 1196.000 1053.310 1200.000 ;
    END
  END cpu_dtr_n1[27]
  PIN cpu_dtr_n1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.150 1196.000 1063.430 1200.000 ;
    END
  END cpu_dtr_n1[28]
  PIN cpu_dtr_n1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.730 1196.000 1074.010 1200.000 ;
    END
  END cpu_dtr_n1[29]
  PIN cpu_dtr_n1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.590 1196.000 793.870 1200.000 ;
    END
  END cpu_dtr_n1[2]
  PIN cpu_dtr_n1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.850 1196.000 1084.130 1200.000 ;
    END
  END cpu_dtr_n1[30]
  PIN cpu_dtr_n1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.430 1196.000 1094.710 1200.000 ;
    END
  END cpu_dtr_n1[31]
  PIN cpu_dtr_n1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.710 1196.000 803.990 1200.000 ;
    END
  END cpu_dtr_n1[3]
  PIN cpu_dtr_n1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 814.290 1196.000 814.570 1200.000 ;
    END
  END cpu_dtr_n1[4]
  PIN cpu_dtr_n1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.410 1196.000 824.690 1200.000 ;
    END
  END cpu_dtr_n1[5]
  PIN cpu_dtr_n1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.990 1196.000 835.270 1200.000 ;
    END
  END cpu_dtr_n1[6]
  PIN cpu_dtr_n1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 845.570 1196.000 845.850 1200.000 ;
    END
  END cpu_dtr_n1[7]
  PIN cpu_dtr_n1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.690 1196.000 855.970 1200.000 ;
    END
  END cpu_dtr_n1[8]
  PIN cpu_dtr_n1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.270 1196.000 866.550 1200.000 ;
    END
  END cpu_dtr_n1[9]
  PIN cpu_dtw_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 665.760 1100.000 666.360 ;
    END
  END cpu_dtw_e[0]
  PIN cpu_dtw_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 775.920 1100.000 776.520 ;
    END
  END cpu_dtw_e[10]
  PIN cpu_dtw_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 786.800 1100.000 787.400 ;
    END
  END cpu_dtw_e[11]
  PIN cpu_dtw_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 797.680 1100.000 798.280 ;
    END
  END cpu_dtw_e[12]
  PIN cpu_dtw_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 809.240 1100.000 809.840 ;
    END
  END cpu_dtw_e[13]
  PIN cpu_dtw_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 820.120 1100.000 820.720 ;
    END
  END cpu_dtw_e[14]
  PIN cpu_dtw_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 831.000 1100.000 831.600 ;
    END
  END cpu_dtw_e[15]
  PIN cpu_dtw_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 676.640 1100.000 677.240 ;
    END
  END cpu_dtw_e[1]
  PIN cpu_dtw_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 687.520 1100.000 688.120 ;
    END
  END cpu_dtw_e[2]
  PIN cpu_dtw_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 699.080 1100.000 699.680 ;
    END
  END cpu_dtw_e[3]
  PIN cpu_dtw_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 709.960 1100.000 710.560 ;
    END
  END cpu_dtw_e[4]
  PIN cpu_dtw_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 720.840 1100.000 721.440 ;
    END
  END cpu_dtw_e[5]
  PIN cpu_dtw_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 731.720 1100.000 732.320 ;
    END
  END cpu_dtw_e[6]
  PIN cpu_dtw_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 742.600 1100.000 743.200 ;
    END
  END cpu_dtw_e[7]
  PIN cpu_dtw_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 754.160 1100.000 754.760 ;
    END
  END cpu_dtw_e[8]
  PIN cpu_dtw_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 765.040 1100.000 765.640 ;
    END
  END cpu_dtw_e[9]
  PIN cpu_dtw_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 606.830 1196.000 607.110 1200.000 ;
    END
  END cpu_dtw_n[0]
  PIN cpu_dtw_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.330 1196.000 710.610 1200.000 ;
    END
  END cpu_dtw_n[10]
  PIN cpu_dtw_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 720.910 1196.000 721.190 1200.000 ;
    END
  END cpu_dtw_n[11]
  PIN cpu_dtw_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.030 1196.000 731.310 1200.000 ;
    END
  END cpu_dtw_n[12]
  PIN cpu_dtw_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 741.610 1196.000 741.890 1200.000 ;
    END
  END cpu_dtw_n[13]
  PIN cpu_dtw_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 752.190 1196.000 752.470 1200.000 ;
    END
  END cpu_dtw_n[14]
  PIN cpu_dtw_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 762.310 1196.000 762.590 1200.000 ;
    END
  END cpu_dtw_n[15]
  PIN cpu_dtw_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 616.950 1196.000 617.230 1200.000 ;
    END
  END cpu_dtw_n[1]
  PIN cpu_dtw_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.530 1196.000 627.810 1200.000 ;
    END
  END cpu_dtw_n[2]
  PIN cpu_dtw_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 637.650 1196.000 637.930 1200.000 ;
    END
  END cpu_dtw_n[3]
  PIN cpu_dtw_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 648.230 1196.000 648.510 1200.000 ;
    END
  END cpu_dtw_n[4]
  PIN cpu_dtw_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 658.810 1196.000 659.090 1200.000 ;
    END
  END cpu_dtw_n[5]
  PIN cpu_dtw_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 668.930 1196.000 669.210 1200.000 ;
    END
  END cpu_dtw_n[6]
  PIN cpu_dtw_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 679.510 1196.000 679.790 1200.000 ;
    END
  END cpu_dtw_n[7]
  PIN cpu_dtw_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.630 1196.000 689.910 1200.000 ;
    END
  END cpu_dtw_n[8]
  PIN cpu_dtw_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 700.210 1196.000 700.490 1200.000 ;
    END
  END cpu_dtw_n[9]
  PIN cpu_mask_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 379.480 1100.000 380.080 ;
    END
  END cpu_mask_e[0]
  PIN cpu_mask_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 390.360 1100.000 390.960 ;
    END
  END cpu_mask_e[1]
  PIN cpu_mask_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 401.240 1100.000 401.840 ;
    END
  END cpu_mask_e[2]
  PIN cpu_mask_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 412.800 1100.000 413.400 ;
    END
  END cpu_mask_e[3]
  PIN cpu_mask_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 423.680 1100.000 424.280 ;
    END
  END cpu_mask_e[4]
  PIN cpu_mask_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 434.560 1100.000 435.160 ;
    END
  END cpu_mask_e[5]
  PIN cpu_mask_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 445.440 1100.000 446.040 ;
    END
  END cpu_mask_e[6]
  PIN cpu_mask_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 456.320 1100.000 456.920 ;
    END
  END cpu_mask_e[7]
  PIN cpu_mask_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.870 1196.000 503.150 1200.000 ;
    END
  END cpu_mask_n[0]
  PIN cpu_mask_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 513.450 1196.000 513.730 1200.000 ;
    END
  END cpu_mask_n[1]
  PIN cpu_mask_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 523.570 1196.000 523.850 1200.000 ;
    END
  END cpu_mask_n[2]
  PIN cpu_mask_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.150 1196.000 534.430 1200.000 ;
    END
  END cpu_mask_n[3]
  PIN cpu_mask_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 544.270 1196.000 544.550 1200.000 ;
    END
  END cpu_mask_n[4]
  PIN cpu_mask_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 554.850 1196.000 555.130 1200.000 ;
    END
  END cpu_mask_n[5]
  PIN cpu_mask_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 565.430 1196.000 565.710 1200.000 ;
    END
  END cpu_mask_n[6]
  PIN cpu_mask_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 575.550 1196.000 575.830 1200.000 ;
    END
  END cpu_mask_n[7]
  PIN cpu_wen_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 467.880 1100.000 468.480 ;
    END
  END cpu_wen_e[0]
  PIN cpu_wen_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 478.760 1100.000 479.360 ;
    END
  END cpu_wen_e[1]
  PIN cpu_wen_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 586.130 1196.000 586.410 1200.000 ;
    END
  END cpu_wen_n[0]
  PIN cpu_wen_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 596.250 1196.000 596.530 1200.000 ;
    END
  END cpu_wen_n[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.800 4.000 447.400 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 762.320 4.000 762.920 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 4.000 794.880 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 857.520 4.000 858.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.800 4.000 889.400 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1015.280 4.000 1015.880 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1046.560 4.000 1047.160 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1078.520 4.000 1079.120 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.800 4.000 1110.400 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.760 4.000 1142.360 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 804.480 4.000 805.080 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 4.000 868.320 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.680 4.000 900.280 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.720 4.000 1089.320 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.680 4.000 1121.280 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.960 4.000 1152.560 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.920 4.000 1184.520 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 783.400 4.000 784.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.120 4.000 973.720 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1004.400 4.000 1005.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.880 4.000 1131.480 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.120 4.000 1194.720 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1065.450 0.000 1065.730 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1075.110 0.000 1075.390 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.430 0.000 1094.710 4.000 ;
    END
  END la_data_out[2]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 4.000 ;
    END
  END la_oen[1]
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 16.360 1100.000 16.960 ;
    END
  END one
  PIN ram_ce
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1194.120 1100.000 1194.720 ;
    END
  END ram_ce
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 802.790 0.000 803.070 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 861.210 0.000 861.490 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 919.170 0.000 919.450 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.610 0.000 948.890 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.590 0.000 977.870 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.030 0.000 1007.310 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.430 0.000 841.710 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 899.850 0.000 900.130 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.270 0.000 958.550 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 987.710 0.000 987.990 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 675.830 0.000 676.110 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 792.670 0.000 792.950 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.530 0.000 880.810 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 938.950 0.000 939.230 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.930 0.000 968.210 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.370 0.000 997.650 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1026.350 0.000 1026.630 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_we_i
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 5.480 1100.000 6.080 ;
    END
  END zero
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1188.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1094.340 1188.725 ;
      LAYER met1 ;
        RECT 5.130 4.460 1094.730 1189.280 ;
      LAYER met2 ;
        RECT 4.760 1195.720 4.870 1196.000 ;
        RECT 5.710 1195.720 14.990 1196.000 ;
        RECT 15.830 1195.720 25.570 1196.000 ;
        RECT 26.410 1195.720 35.690 1196.000 ;
        RECT 36.530 1195.720 46.270 1196.000 ;
        RECT 47.110 1195.720 56.390 1196.000 ;
        RECT 57.230 1195.720 66.970 1196.000 ;
        RECT 67.810 1195.720 77.090 1196.000 ;
        RECT 77.930 1195.720 87.670 1196.000 ;
        RECT 88.510 1195.720 98.250 1196.000 ;
        RECT 99.090 1195.720 108.370 1196.000 ;
        RECT 109.210 1195.720 118.950 1196.000 ;
        RECT 119.790 1195.720 129.070 1196.000 ;
        RECT 129.910 1195.720 139.650 1196.000 ;
        RECT 140.490 1195.720 149.770 1196.000 ;
        RECT 150.610 1195.720 160.350 1196.000 ;
        RECT 161.190 1195.720 170.470 1196.000 ;
        RECT 171.310 1195.720 181.050 1196.000 ;
        RECT 181.890 1195.720 191.630 1196.000 ;
        RECT 192.470 1195.720 201.750 1196.000 ;
        RECT 202.590 1195.720 212.330 1196.000 ;
        RECT 213.170 1195.720 222.450 1196.000 ;
        RECT 223.290 1195.720 233.030 1196.000 ;
        RECT 233.870 1195.720 243.150 1196.000 ;
        RECT 243.990 1195.720 253.730 1196.000 ;
        RECT 254.570 1195.720 263.850 1196.000 ;
        RECT 264.690 1195.720 274.430 1196.000 ;
        RECT 275.270 1195.720 285.010 1196.000 ;
        RECT 285.850 1195.720 295.130 1196.000 ;
        RECT 295.970 1195.720 305.710 1196.000 ;
        RECT 306.550 1195.720 315.830 1196.000 ;
        RECT 316.670 1195.720 326.410 1196.000 ;
        RECT 327.250 1195.720 336.530 1196.000 ;
        RECT 337.370 1195.720 347.110 1196.000 ;
        RECT 347.950 1195.720 357.230 1196.000 ;
        RECT 358.070 1195.720 367.810 1196.000 ;
        RECT 368.650 1195.720 378.390 1196.000 ;
        RECT 379.230 1195.720 388.510 1196.000 ;
        RECT 389.350 1195.720 399.090 1196.000 ;
        RECT 399.930 1195.720 409.210 1196.000 ;
        RECT 410.050 1195.720 419.790 1196.000 ;
        RECT 420.630 1195.720 429.910 1196.000 ;
        RECT 430.750 1195.720 440.490 1196.000 ;
        RECT 441.330 1195.720 450.610 1196.000 ;
        RECT 451.450 1195.720 461.190 1196.000 ;
        RECT 462.030 1195.720 471.770 1196.000 ;
        RECT 472.610 1195.720 481.890 1196.000 ;
        RECT 482.730 1195.720 492.470 1196.000 ;
        RECT 493.310 1195.720 502.590 1196.000 ;
        RECT 503.430 1195.720 513.170 1196.000 ;
        RECT 514.010 1195.720 523.290 1196.000 ;
        RECT 524.130 1195.720 533.870 1196.000 ;
        RECT 534.710 1195.720 543.990 1196.000 ;
        RECT 544.830 1195.720 554.570 1196.000 ;
        RECT 555.410 1195.720 565.150 1196.000 ;
        RECT 565.990 1195.720 575.270 1196.000 ;
        RECT 576.110 1195.720 585.850 1196.000 ;
        RECT 586.690 1195.720 595.970 1196.000 ;
        RECT 596.810 1195.720 606.550 1196.000 ;
        RECT 607.390 1195.720 616.670 1196.000 ;
        RECT 617.510 1195.720 627.250 1196.000 ;
        RECT 628.090 1195.720 637.370 1196.000 ;
        RECT 638.210 1195.720 647.950 1196.000 ;
        RECT 648.790 1195.720 658.530 1196.000 ;
        RECT 659.370 1195.720 668.650 1196.000 ;
        RECT 669.490 1195.720 679.230 1196.000 ;
        RECT 680.070 1195.720 689.350 1196.000 ;
        RECT 690.190 1195.720 699.930 1196.000 ;
        RECT 700.770 1195.720 710.050 1196.000 ;
        RECT 710.890 1195.720 720.630 1196.000 ;
        RECT 721.470 1195.720 730.750 1196.000 ;
        RECT 731.590 1195.720 741.330 1196.000 ;
        RECT 742.170 1195.720 751.910 1196.000 ;
        RECT 752.750 1195.720 762.030 1196.000 ;
        RECT 762.870 1195.720 772.610 1196.000 ;
        RECT 773.450 1195.720 782.730 1196.000 ;
        RECT 783.570 1195.720 793.310 1196.000 ;
        RECT 794.150 1195.720 803.430 1196.000 ;
        RECT 804.270 1195.720 814.010 1196.000 ;
        RECT 814.850 1195.720 824.130 1196.000 ;
        RECT 824.970 1195.720 834.710 1196.000 ;
        RECT 835.550 1195.720 845.290 1196.000 ;
        RECT 846.130 1195.720 855.410 1196.000 ;
        RECT 856.250 1195.720 865.990 1196.000 ;
        RECT 866.830 1195.720 876.110 1196.000 ;
        RECT 876.950 1195.720 886.690 1196.000 ;
        RECT 887.530 1195.720 896.810 1196.000 ;
        RECT 897.650 1195.720 907.390 1196.000 ;
        RECT 908.230 1195.720 917.510 1196.000 ;
        RECT 918.350 1195.720 928.090 1196.000 ;
        RECT 928.930 1195.720 938.670 1196.000 ;
        RECT 939.510 1195.720 948.790 1196.000 ;
        RECT 949.630 1195.720 959.370 1196.000 ;
        RECT 960.210 1195.720 969.490 1196.000 ;
        RECT 970.330 1195.720 980.070 1196.000 ;
        RECT 980.910 1195.720 990.190 1196.000 ;
        RECT 991.030 1195.720 1000.770 1196.000 ;
        RECT 1001.610 1195.720 1010.890 1196.000 ;
        RECT 1011.730 1195.720 1021.470 1196.000 ;
        RECT 1022.310 1195.720 1032.050 1196.000 ;
        RECT 1032.890 1195.720 1042.170 1196.000 ;
        RECT 1043.010 1195.720 1052.750 1196.000 ;
        RECT 1053.590 1195.720 1062.870 1196.000 ;
        RECT 1063.710 1195.720 1073.450 1196.000 ;
        RECT 1074.290 1195.720 1083.570 1196.000 ;
        RECT 1084.410 1195.720 1094.150 1196.000 ;
        RECT 1094.990 1195.720 1095.630 1196.000 ;
        RECT 4.760 4.280 1095.630 1195.720 ;
        RECT 5.250 4.000 14.070 4.280 ;
        RECT 14.910 4.000 23.730 4.280 ;
        RECT 24.570 4.000 33.390 4.280 ;
        RECT 34.230 4.000 43.050 4.280 ;
        RECT 43.890 4.000 52.710 4.280 ;
        RECT 53.550 4.000 62.370 4.280 ;
        RECT 63.210 4.000 72.490 4.280 ;
        RECT 73.330 4.000 82.150 4.280 ;
        RECT 82.990 4.000 91.810 4.280 ;
        RECT 92.650 4.000 101.470 4.280 ;
        RECT 102.310 4.000 111.130 4.280 ;
        RECT 111.970 4.000 120.790 4.280 ;
        RECT 121.630 4.000 130.910 4.280 ;
        RECT 131.750 4.000 140.570 4.280 ;
        RECT 141.410 4.000 150.230 4.280 ;
        RECT 151.070 4.000 159.890 4.280 ;
        RECT 160.730 4.000 169.550 4.280 ;
        RECT 170.390 4.000 179.210 4.280 ;
        RECT 180.050 4.000 189.330 4.280 ;
        RECT 190.170 4.000 198.990 4.280 ;
        RECT 199.830 4.000 208.650 4.280 ;
        RECT 209.490 4.000 218.310 4.280 ;
        RECT 219.150 4.000 227.970 4.280 ;
        RECT 228.810 4.000 237.630 4.280 ;
        RECT 238.470 4.000 247.290 4.280 ;
        RECT 248.130 4.000 257.410 4.280 ;
        RECT 258.250 4.000 267.070 4.280 ;
        RECT 267.910 4.000 276.730 4.280 ;
        RECT 277.570 4.000 286.390 4.280 ;
        RECT 287.230 4.000 296.050 4.280 ;
        RECT 296.890 4.000 305.710 4.280 ;
        RECT 306.550 4.000 315.830 4.280 ;
        RECT 316.670 4.000 325.490 4.280 ;
        RECT 326.330 4.000 335.150 4.280 ;
        RECT 335.990 4.000 344.810 4.280 ;
        RECT 345.650 4.000 354.470 4.280 ;
        RECT 355.310 4.000 364.130 4.280 ;
        RECT 364.970 4.000 374.250 4.280 ;
        RECT 375.090 4.000 383.910 4.280 ;
        RECT 384.750 4.000 393.570 4.280 ;
        RECT 394.410 4.000 403.230 4.280 ;
        RECT 404.070 4.000 412.890 4.280 ;
        RECT 413.730 4.000 422.550 4.280 ;
        RECT 423.390 4.000 432.670 4.280 ;
        RECT 433.510 4.000 442.330 4.280 ;
        RECT 443.170 4.000 451.990 4.280 ;
        RECT 452.830 4.000 461.650 4.280 ;
        RECT 462.490 4.000 471.310 4.280 ;
        RECT 472.150 4.000 480.970 4.280 ;
        RECT 481.810 4.000 490.630 4.280 ;
        RECT 491.470 4.000 500.750 4.280 ;
        RECT 501.590 4.000 510.410 4.280 ;
        RECT 511.250 4.000 520.070 4.280 ;
        RECT 520.910 4.000 529.730 4.280 ;
        RECT 530.570 4.000 539.390 4.280 ;
        RECT 540.230 4.000 549.050 4.280 ;
        RECT 549.890 4.000 559.170 4.280 ;
        RECT 560.010 4.000 568.830 4.280 ;
        RECT 569.670 4.000 578.490 4.280 ;
        RECT 579.330 4.000 588.150 4.280 ;
        RECT 588.990 4.000 597.810 4.280 ;
        RECT 598.650 4.000 607.470 4.280 ;
        RECT 608.310 4.000 617.590 4.280 ;
        RECT 618.430 4.000 627.250 4.280 ;
        RECT 628.090 4.000 636.910 4.280 ;
        RECT 637.750 4.000 646.570 4.280 ;
        RECT 647.410 4.000 656.230 4.280 ;
        RECT 657.070 4.000 665.890 4.280 ;
        RECT 666.730 4.000 675.550 4.280 ;
        RECT 676.390 4.000 685.670 4.280 ;
        RECT 686.510 4.000 695.330 4.280 ;
        RECT 696.170 4.000 704.990 4.280 ;
        RECT 705.830 4.000 714.650 4.280 ;
        RECT 715.490 4.000 724.310 4.280 ;
        RECT 725.150 4.000 733.970 4.280 ;
        RECT 734.810 4.000 744.090 4.280 ;
        RECT 744.930 4.000 753.750 4.280 ;
        RECT 754.590 4.000 763.410 4.280 ;
        RECT 764.250 4.000 773.070 4.280 ;
        RECT 773.910 4.000 782.730 4.280 ;
        RECT 783.570 4.000 792.390 4.280 ;
        RECT 793.230 4.000 802.510 4.280 ;
        RECT 803.350 4.000 812.170 4.280 ;
        RECT 813.010 4.000 821.830 4.280 ;
        RECT 822.670 4.000 831.490 4.280 ;
        RECT 832.330 4.000 841.150 4.280 ;
        RECT 841.990 4.000 850.810 4.280 ;
        RECT 851.650 4.000 860.930 4.280 ;
        RECT 861.770 4.000 870.590 4.280 ;
        RECT 871.430 4.000 880.250 4.280 ;
        RECT 881.090 4.000 889.910 4.280 ;
        RECT 890.750 4.000 899.570 4.280 ;
        RECT 900.410 4.000 909.230 4.280 ;
        RECT 910.070 4.000 918.890 4.280 ;
        RECT 919.730 4.000 929.010 4.280 ;
        RECT 929.850 4.000 938.670 4.280 ;
        RECT 939.510 4.000 948.330 4.280 ;
        RECT 949.170 4.000 957.990 4.280 ;
        RECT 958.830 4.000 967.650 4.280 ;
        RECT 968.490 4.000 977.310 4.280 ;
        RECT 978.150 4.000 987.430 4.280 ;
        RECT 988.270 4.000 997.090 4.280 ;
        RECT 997.930 4.000 1006.750 4.280 ;
        RECT 1007.590 4.000 1016.410 4.280 ;
        RECT 1017.250 4.000 1026.070 4.280 ;
        RECT 1026.910 4.000 1035.730 4.280 ;
        RECT 1036.570 4.000 1045.850 4.280 ;
        RECT 1046.690 4.000 1055.510 4.280 ;
        RECT 1056.350 4.000 1065.170 4.280 ;
        RECT 1066.010 4.000 1074.830 4.280 ;
        RECT 1075.670 4.000 1084.490 4.280 ;
        RECT 1085.330 4.000 1094.150 4.280 ;
        RECT 1094.990 4.000 1095.630 4.280 ;
      LAYER met3 ;
        RECT 4.400 1193.720 1095.600 1194.585 ;
        RECT 3.990 1184.920 1096.000 1193.720 ;
        RECT 4.400 1184.240 1096.000 1184.920 ;
        RECT 4.400 1183.520 1095.600 1184.240 ;
        RECT 3.990 1182.840 1095.600 1183.520 ;
        RECT 3.990 1174.040 1096.000 1182.840 ;
        RECT 4.400 1173.360 1096.000 1174.040 ;
        RECT 4.400 1172.640 1095.600 1173.360 ;
        RECT 3.990 1171.960 1095.600 1172.640 ;
        RECT 3.990 1163.840 1096.000 1171.960 ;
        RECT 4.400 1162.480 1096.000 1163.840 ;
        RECT 4.400 1162.440 1095.600 1162.480 ;
        RECT 3.990 1161.080 1095.600 1162.440 ;
        RECT 3.990 1152.960 1096.000 1161.080 ;
        RECT 4.400 1151.600 1096.000 1152.960 ;
        RECT 4.400 1151.560 1095.600 1151.600 ;
        RECT 3.990 1150.200 1095.600 1151.560 ;
        RECT 3.990 1142.760 1096.000 1150.200 ;
        RECT 4.400 1141.360 1096.000 1142.760 ;
        RECT 3.990 1140.040 1096.000 1141.360 ;
        RECT 3.990 1138.640 1095.600 1140.040 ;
        RECT 3.990 1131.880 1096.000 1138.640 ;
        RECT 4.400 1130.480 1096.000 1131.880 ;
        RECT 3.990 1129.160 1096.000 1130.480 ;
        RECT 3.990 1127.760 1095.600 1129.160 ;
        RECT 3.990 1121.680 1096.000 1127.760 ;
        RECT 4.400 1120.280 1096.000 1121.680 ;
        RECT 3.990 1118.280 1096.000 1120.280 ;
        RECT 3.990 1116.880 1095.600 1118.280 ;
        RECT 3.990 1110.800 1096.000 1116.880 ;
        RECT 4.400 1109.400 1096.000 1110.800 ;
        RECT 3.990 1107.400 1096.000 1109.400 ;
        RECT 3.990 1106.000 1095.600 1107.400 ;
        RECT 3.990 1100.600 1096.000 1106.000 ;
        RECT 4.400 1099.200 1096.000 1100.600 ;
        RECT 3.990 1096.520 1096.000 1099.200 ;
        RECT 3.990 1095.120 1095.600 1096.520 ;
        RECT 3.990 1089.720 1096.000 1095.120 ;
        RECT 4.400 1088.320 1096.000 1089.720 ;
        RECT 3.990 1084.960 1096.000 1088.320 ;
        RECT 3.990 1083.560 1095.600 1084.960 ;
        RECT 3.990 1079.520 1096.000 1083.560 ;
        RECT 4.400 1078.120 1096.000 1079.520 ;
        RECT 3.990 1074.080 1096.000 1078.120 ;
        RECT 3.990 1072.680 1095.600 1074.080 ;
        RECT 3.990 1068.640 1096.000 1072.680 ;
        RECT 4.400 1067.240 1096.000 1068.640 ;
        RECT 3.990 1063.200 1096.000 1067.240 ;
        RECT 3.990 1061.800 1095.600 1063.200 ;
        RECT 3.990 1058.440 1096.000 1061.800 ;
        RECT 4.400 1057.040 1096.000 1058.440 ;
        RECT 3.990 1052.320 1096.000 1057.040 ;
        RECT 3.990 1050.920 1095.600 1052.320 ;
        RECT 3.990 1047.560 1096.000 1050.920 ;
        RECT 4.400 1046.160 1096.000 1047.560 ;
        RECT 3.990 1041.440 1096.000 1046.160 ;
        RECT 3.990 1040.040 1095.600 1041.440 ;
        RECT 3.990 1037.360 1096.000 1040.040 ;
        RECT 4.400 1035.960 1096.000 1037.360 ;
        RECT 3.990 1029.880 1096.000 1035.960 ;
        RECT 3.990 1028.480 1095.600 1029.880 ;
        RECT 3.990 1026.480 1096.000 1028.480 ;
        RECT 4.400 1025.080 1096.000 1026.480 ;
        RECT 3.990 1019.000 1096.000 1025.080 ;
        RECT 3.990 1017.600 1095.600 1019.000 ;
        RECT 3.990 1016.280 1096.000 1017.600 ;
        RECT 4.400 1014.880 1096.000 1016.280 ;
        RECT 3.990 1008.120 1096.000 1014.880 ;
        RECT 3.990 1006.720 1095.600 1008.120 ;
        RECT 3.990 1005.400 1096.000 1006.720 ;
        RECT 4.400 1004.000 1096.000 1005.400 ;
        RECT 3.990 997.240 1096.000 1004.000 ;
        RECT 3.990 995.840 1095.600 997.240 ;
        RECT 3.990 995.200 1096.000 995.840 ;
        RECT 4.400 993.800 1096.000 995.200 ;
        RECT 3.990 986.360 1096.000 993.800 ;
        RECT 3.990 984.960 1095.600 986.360 ;
        RECT 3.990 984.320 1096.000 984.960 ;
        RECT 4.400 982.920 1096.000 984.320 ;
        RECT 3.990 974.800 1096.000 982.920 ;
        RECT 3.990 974.120 1095.600 974.800 ;
        RECT 4.400 973.400 1095.600 974.120 ;
        RECT 4.400 972.720 1096.000 973.400 ;
        RECT 3.990 963.920 1096.000 972.720 ;
        RECT 3.990 963.240 1095.600 963.920 ;
        RECT 4.400 962.520 1095.600 963.240 ;
        RECT 4.400 961.840 1096.000 962.520 ;
        RECT 3.990 953.040 1096.000 961.840 ;
        RECT 4.400 951.640 1095.600 953.040 ;
        RECT 3.990 942.160 1096.000 951.640 ;
        RECT 4.400 940.760 1095.600 942.160 ;
        RECT 3.990 931.960 1096.000 940.760 ;
        RECT 4.400 931.280 1096.000 931.960 ;
        RECT 4.400 930.560 1095.600 931.280 ;
        RECT 3.990 929.880 1095.600 930.560 ;
        RECT 3.990 921.080 1096.000 929.880 ;
        RECT 4.400 919.720 1096.000 921.080 ;
        RECT 4.400 919.680 1095.600 919.720 ;
        RECT 3.990 918.320 1095.600 919.680 ;
        RECT 3.990 910.880 1096.000 918.320 ;
        RECT 4.400 909.480 1096.000 910.880 ;
        RECT 3.990 908.840 1096.000 909.480 ;
        RECT 3.990 907.440 1095.600 908.840 ;
        RECT 3.990 900.680 1096.000 907.440 ;
        RECT 4.400 899.280 1096.000 900.680 ;
        RECT 3.990 897.960 1096.000 899.280 ;
        RECT 3.990 896.560 1095.600 897.960 ;
        RECT 3.990 889.800 1096.000 896.560 ;
        RECT 4.400 888.400 1096.000 889.800 ;
        RECT 3.990 887.080 1096.000 888.400 ;
        RECT 3.990 885.680 1095.600 887.080 ;
        RECT 3.990 879.600 1096.000 885.680 ;
        RECT 4.400 878.200 1096.000 879.600 ;
        RECT 3.990 876.200 1096.000 878.200 ;
        RECT 3.990 874.800 1095.600 876.200 ;
        RECT 3.990 868.720 1096.000 874.800 ;
        RECT 4.400 867.320 1096.000 868.720 ;
        RECT 3.990 865.320 1096.000 867.320 ;
        RECT 3.990 863.920 1095.600 865.320 ;
        RECT 3.990 858.520 1096.000 863.920 ;
        RECT 4.400 857.120 1096.000 858.520 ;
        RECT 3.990 853.760 1096.000 857.120 ;
        RECT 3.990 852.360 1095.600 853.760 ;
        RECT 3.990 847.640 1096.000 852.360 ;
        RECT 4.400 846.240 1096.000 847.640 ;
        RECT 3.990 842.880 1096.000 846.240 ;
        RECT 3.990 841.480 1095.600 842.880 ;
        RECT 3.990 837.440 1096.000 841.480 ;
        RECT 4.400 836.040 1096.000 837.440 ;
        RECT 3.990 832.000 1096.000 836.040 ;
        RECT 3.990 830.600 1095.600 832.000 ;
        RECT 3.990 826.560 1096.000 830.600 ;
        RECT 4.400 825.160 1096.000 826.560 ;
        RECT 3.990 821.120 1096.000 825.160 ;
        RECT 3.990 819.720 1095.600 821.120 ;
        RECT 3.990 816.360 1096.000 819.720 ;
        RECT 4.400 814.960 1096.000 816.360 ;
        RECT 3.990 810.240 1096.000 814.960 ;
        RECT 3.990 808.840 1095.600 810.240 ;
        RECT 3.990 805.480 1096.000 808.840 ;
        RECT 4.400 804.080 1096.000 805.480 ;
        RECT 3.990 798.680 1096.000 804.080 ;
        RECT 3.990 797.280 1095.600 798.680 ;
        RECT 3.990 795.280 1096.000 797.280 ;
        RECT 4.400 793.880 1096.000 795.280 ;
        RECT 3.990 787.800 1096.000 793.880 ;
        RECT 3.990 786.400 1095.600 787.800 ;
        RECT 3.990 784.400 1096.000 786.400 ;
        RECT 4.400 783.000 1096.000 784.400 ;
        RECT 3.990 776.920 1096.000 783.000 ;
        RECT 3.990 775.520 1095.600 776.920 ;
        RECT 3.990 774.200 1096.000 775.520 ;
        RECT 4.400 772.800 1096.000 774.200 ;
        RECT 3.990 766.040 1096.000 772.800 ;
        RECT 3.990 764.640 1095.600 766.040 ;
        RECT 3.990 763.320 1096.000 764.640 ;
        RECT 4.400 761.920 1096.000 763.320 ;
        RECT 3.990 755.160 1096.000 761.920 ;
        RECT 3.990 753.760 1095.600 755.160 ;
        RECT 3.990 753.120 1096.000 753.760 ;
        RECT 4.400 751.720 1096.000 753.120 ;
        RECT 3.990 743.600 1096.000 751.720 ;
        RECT 3.990 742.240 1095.600 743.600 ;
        RECT 4.400 742.200 1095.600 742.240 ;
        RECT 4.400 740.840 1096.000 742.200 ;
        RECT 3.990 732.720 1096.000 740.840 ;
        RECT 3.990 732.040 1095.600 732.720 ;
        RECT 4.400 731.320 1095.600 732.040 ;
        RECT 4.400 730.640 1096.000 731.320 ;
        RECT 3.990 721.840 1096.000 730.640 ;
        RECT 3.990 721.160 1095.600 721.840 ;
        RECT 4.400 720.440 1095.600 721.160 ;
        RECT 4.400 719.760 1096.000 720.440 ;
        RECT 3.990 710.960 1096.000 719.760 ;
        RECT 4.400 709.560 1095.600 710.960 ;
        RECT 3.990 700.080 1096.000 709.560 ;
        RECT 4.400 698.680 1095.600 700.080 ;
        RECT 3.990 689.880 1096.000 698.680 ;
        RECT 4.400 688.520 1096.000 689.880 ;
        RECT 4.400 688.480 1095.600 688.520 ;
        RECT 3.990 687.120 1095.600 688.480 ;
        RECT 3.990 679.000 1096.000 687.120 ;
        RECT 4.400 677.640 1096.000 679.000 ;
        RECT 4.400 677.600 1095.600 677.640 ;
        RECT 3.990 676.240 1095.600 677.600 ;
        RECT 3.990 668.800 1096.000 676.240 ;
        RECT 4.400 667.400 1096.000 668.800 ;
        RECT 3.990 666.760 1096.000 667.400 ;
        RECT 3.990 665.360 1095.600 666.760 ;
        RECT 3.990 657.920 1096.000 665.360 ;
        RECT 4.400 656.520 1096.000 657.920 ;
        RECT 3.990 655.880 1096.000 656.520 ;
        RECT 3.990 654.480 1095.600 655.880 ;
        RECT 3.990 647.720 1096.000 654.480 ;
        RECT 4.400 646.320 1096.000 647.720 ;
        RECT 3.990 645.000 1096.000 646.320 ;
        RECT 3.990 643.600 1095.600 645.000 ;
        RECT 3.990 636.840 1096.000 643.600 ;
        RECT 4.400 635.440 1096.000 636.840 ;
        RECT 3.990 633.440 1096.000 635.440 ;
        RECT 3.990 632.040 1095.600 633.440 ;
        RECT 3.990 626.640 1096.000 632.040 ;
        RECT 4.400 625.240 1096.000 626.640 ;
        RECT 3.990 622.560 1096.000 625.240 ;
        RECT 3.990 621.160 1095.600 622.560 ;
        RECT 3.990 615.760 1096.000 621.160 ;
        RECT 4.400 614.360 1096.000 615.760 ;
        RECT 3.990 611.680 1096.000 614.360 ;
        RECT 3.990 610.280 1095.600 611.680 ;
        RECT 3.990 605.560 1096.000 610.280 ;
        RECT 4.400 604.160 1096.000 605.560 ;
        RECT 3.990 600.800 1096.000 604.160 ;
        RECT 3.990 599.400 1095.600 600.800 ;
        RECT 3.990 595.360 1096.000 599.400 ;
        RECT 4.400 593.960 1096.000 595.360 ;
        RECT 3.990 589.920 1096.000 593.960 ;
        RECT 3.990 588.520 1095.600 589.920 ;
        RECT 3.990 584.480 1096.000 588.520 ;
        RECT 4.400 583.080 1096.000 584.480 ;
        RECT 3.990 579.040 1096.000 583.080 ;
        RECT 3.990 577.640 1095.600 579.040 ;
        RECT 3.990 574.280 1096.000 577.640 ;
        RECT 4.400 572.880 1096.000 574.280 ;
        RECT 3.990 567.480 1096.000 572.880 ;
        RECT 3.990 566.080 1095.600 567.480 ;
        RECT 3.990 563.400 1096.000 566.080 ;
        RECT 4.400 562.000 1096.000 563.400 ;
        RECT 3.990 556.600 1096.000 562.000 ;
        RECT 3.990 555.200 1095.600 556.600 ;
        RECT 3.990 553.200 1096.000 555.200 ;
        RECT 4.400 551.800 1096.000 553.200 ;
        RECT 3.990 545.720 1096.000 551.800 ;
        RECT 3.990 544.320 1095.600 545.720 ;
        RECT 3.990 542.320 1096.000 544.320 ;
        RECT 4.400 540.920 1096.000 542.320 ;
        RECT 3.990 534.840 1096.000 540.920 ;
        RECT 3.990 533.440 1095.600 534.840 ;
        RECT 3.990 532.120 1096.000 533.440 ;
        RECT 4.400 530.720 1096.000 532.120 ;
        RECT 3.990 523.960 1096.000 530.720 ;
        RECT 3.990 522.560 1095.600 523.960 ;
        RECT 3.990 521.240 1096.000 522.560 ;
        RECT 4.400 519.840 1096.000 521.240 ;
        RECT 3.990 512.400 1096.000 519.840 ;
        RECT 3.990 511.040 1095.600 512.400 ;
        RECT 4.400 511.000 1095.600 511.040 ;
        RECT 4.400 509.640 1096.000 511.000 ;
        RECT 3.990 501.520 1096.000 509.640 ;
        RECT 3.990 500.160 1095.600 501.520 ;
        RECT 4.400 500.120 1095.600 500.160 ;
        RECT 4.400 498.760 1096.000 500.120 ;
        RECT 3.990 490.640 1096.000 498.760 ;
        RECT 3.990 489.960 1095.600 490.640 ;
        RECT 4.400 489.240 1095.600 489.960 ;
        RECT 4.400 488.560 1096.000 489.240 ;
        RECT 3.990 479.760 1096.000 488.560 ;
        RECT 3.990 479.080 1095.600 479.760 ;
        RECT 4.400 478.360 1095.600 479.080 ;
        RECT 4.400 477.680 1096.000 478.360 ;
        RECT 3.990 468.880 1096.000 477.680 ;
        RECT 4.400 467.480 1095.600 468.880 ;
        RECT 3.990 458.000 1096.000 467.480 ;
        RECT 4.400 457.320 1096.000 458.000 ;
        RECT 4.400 456.600 1095.600 457.320 ;
        RECT 3.990 455.920 1095.600 456.600 ;
        RECT 3.990 447.800 1096.000 455.920 ;
        RECT 4.400 446.440 1096.000 447.800 ;
        RECT 4.400 446.400 1095.600 446.440 ;
        RECT 3.990 445.040 1095.600 446.400 ;
        RECT 3.990 436.920 1096.000 445.040 ;
        RECT 4.400 435.560 1096.000 436.920 ;
        RECT 4.400 435.520 1095.600 435.560 ;
        RECT 3.990 434.160 1095.600 435.520 ;
        RECT 3.990 426.720 1096.000 434.160 ;
        RECT 4.400 425.320 1096.000 426.720 ;
        RECT 3.990 424.680 1096.000 425.320 ;
        RECT 3.990 423.280 1095.600 424.680 ;
        RECT 3.990 415.840 1096.000 423.280 ;
        RECT 4.400 414.440 1096.000 415.840 ;
        RECT 3.990 413.800 1096.000 414.440 ;
        RECT 3.990 412.400 1095.600 413.800 ;
        RECT 3.990 405.640 1096.000 412.400 ;
        RECT 4.400 404.240 1096.000 405.640 ;
        RECT 3.990 402.240 1096.000 404.240 ;
        RECT 3.990 400.840 1095.600 402.240 ;
        RECT 3.990 394.760 1096.000 400.840 ;
        RECT 4.400 393.360 1096.000 394.760 ;
        RECT 3.990 391.360 1096.000 393.360 ;
        RECT 3.990 389.960 1095.600 391.360 ;
        RECT 3.990 384.560 1096.000 389.960 ;
        RECT 4.400 383.160 1096.000 384.560 ;
        RECT 3.990 380.480 1096.000 383.160 ;
        RECT 3.990 379.080 1095.600 380.480 ;
        RECT 3.990 373.680 1096.000 379.080 ;
        RECT 4.400 372.280 1096.000 373.680 ;
        RECT 3.990 369.600 1096.000 372.280 ;
        RECT 3.990 368.200 1095.600 369.600 ;
        RECT 3.990 363.480 1096.000 368.200 ;
        RECT 4.400 362.080 1096.000 363.480 ;
        RECT 3.990 358.720 1096.000 362.080 ;
        RECT 3.990 357.320 1095.600 358.720 ;
        RECT 3.990 352.600 1096.000 357.320 ;
        RECT 4.400 351.200 1096.000 352.600 ;
        RECT 3.990 347.160 1096.000 351.200 ;
        RECT 3.990 345.760 1095.600 347.160 ;
        RECT 3.990 342.400 1096.000 345.760 ;
        RECT 4.400 341.000 1096.000 342.400 ;
        RECT 3.990 336.280 1096.000 341.000 ;
        RECT 3.990 334.880 1095.600 336.280 ;
        RECT 3.990 331.520 1096.000 334.880 ;
        RECT 4.400 330.120 1096.000 331.520 ;
        RECT 3.990 325.400 1096.000 330.120 ;
        RECT 3.990 324.000 1095.600 325.400 ;
        RECT 3.990 321.320 1096.000 324.000 ;
        RECT 4.400 319.920 1096.000 321.320 ;
        RECT 3.990 314.520 1096.000 319.920 ;
        RECT 3.990 313.120 1095.600 314.520 ;
        RECT 3.990 310.440 1096.000 313.120 ;
        RECT 4.400 309.040 1096.000 310.440 ;
        RECT 3.990 303.640 1096.000 309.040 ;
        RECT 3.990 302.240 1095.600 303.640 ;
        RECT 3.990 300.240 1096.000 302.240 ;
        RECT 4.400 298.840 1096.000 300.240 ;
        RECT 3.990 292.760 1096.000 298.840 ;
        RECT 3.990 291.360 1095.600 292.760 ;
        RECT 3.990 290.040 1096.000 291.360 ;
        RECT 4.400 288.640 1096.000 290.040 ;
        RECT 3.990 281.200 1096.000 288.640 ;
        RECT 3.990 279.800 1095.600 281.200 ;
        RECT 3.990 279.160 1096.000 279.800 ;
        RECT 4.400 277.760 1096.000 279.160 ;
        RECT 3.990 270.320 1096.000 277.760 ;
        RECT 3.990 268.960 1095.600 270.320 ;
        RECT 4.400 268.920 1095.600 268.960 ;
        RECT 4.400 267.560 1096.000 268.920 ;
        RECT 3.990 259.440 1096.000 267.560 ;
        RECT 3.990 258.080 1095.600 259.440 ;
        RECT 4.400 258.040 1095.600 258.080 ;
        RECT 4.400 256.680 1096.000 258.040 ;
        RECT 3.990 248.560 1096.000 256.680 ;
        RECT 3.990 247.880 1095.600 248.560 ;
        RECT 4.400 247.160 1095.600 247.880 ;
        RECT 4.400 246.480 1096.000 247.160 ;
        RECT 3.990 237.680 1096.000 246.480 ;
        RECT 3.990 237.000 1095.600 237.680 ;
        RECT 4.400 236.280 1095.600 237.000 ;
        RECT 4.400 235.600 1096.000 236.280 ;
        RECT 3.990 226.800 1096.000 235.600 ;
        RECT 4.400 226.120 1096.000 226.800 ;
        RECT 4.400 225.400 1095.600 226.120 ;
        RECT 3.990 224.720 1095.600 225.400 ;
        RECT 3.990 215.920 1096.000 224.720 ;
        RECT 4.400 215.240 1096.000 215.920 ;
        RECT 4.400 214.520 1095.600 215.240 ;
        RECT 3.990 213.840 1095.600 214.520 ;
        RECT 3.990 205.720 1096.000 213.840 ;
        RECT 4.400 204.360 1096.000 205.720 ;
        RECT 4.400 204.320 1095.600 204.360 ;
        RECT 3.990 202.960 1095.600 204.320 ;
        RECT 3.990 194.840 1096.000 202.960 ;
        RECT 4.400 193.480 1096.000 194.840 ;
        RECT 4.400 193.440 1095.600 193.480 ;
        RECT 3.990 192.080 1095.600 193.440 ;
        RECT 3.990 184.640 1096.000 192.080 ;
        RECT 4.400 183.240 1096.000 184.640 ;
        RECT 3.990 182.600 1096.000 183.240 ;
        RECT 3.990 181.200 1095.600 182.600 ;
        RECT 3.990 173.760 1096.000 181.200 ;
        RECT 4.400 172.360 1096.000 173.760 ;
        RECT 3.990 171.040 1096.000 172.360 ;
        RECT 3.990 169.640 1095.600 171.040 ;
        RECT 3.990 163.560 1096.000 169.640 ;
        RECT 4.400 162.160 1096.000 163.560 ;
        RECT 3.990 160.160 1096.000 162.160 ;
        RECT 3.990 158.760 1095.600 160.160 ;
        RECT 3.990 152.680 1096.000 158.760 ;
        RECT 4.400 151.280 1096.000 152.680 ;
        RECT 3.990 149.280 1096.000 151.280 ;
        RECT 3.990 147.880 1095.600 149.280 ;
        RECT 3.990 142.480 1096.000 147.880 ;
        RECT 4.400 141.080 1096.000 142.480 ;
        RECT 3.990 138.400 1096.000 141.080 ;
        RECT 3.990 137.000 1095.600 138.400 ;
        RECT 3.990 131.600 1096.000 137.000 ;
        RECT 4.400 130.200 1096.000 131.600 ;
        RECT 3.990 127.520 1096.000 130.200 ;
        RECT 3.990 126.120 1095.600 127.520 ;
        RECT 3.990 121.400 1096.000 126.120 ;
        RECT 4.400 120.000 1096.000 121.400 ;
        RECT 3.990 115.960 1096.000 120.000 ;
        RECT 3.990 114.560 1095.600 115.960 ;
        RECT 3.990 110.520 1096.000 114.560 ;
        RECT 4.400 109.120 1096.000 110.520 ;
        RECT 3.990 105.080 1096.000 109.120 ;
        RECT 3.990 103.680 1095.600 105.080 ;
        RECT 3.990 100.320 1096.000 103.680 ;
        RECT 4.400 98.920 1096.000 100.320 ;
        RECT 3.990 94.200 1096.000 98.920 ;
        RECT 3.990 92.800 1095.600 94.200 ;
        RECT 3.990 89.440 1096.000 92.800 ;
        RECT 4.400 88.040 1096.000 89.440 ;
        RECT 3.990 83.320 1096.000 88.040 ;
        RECT 3.990 81.920 1095.600 83.320 ;
        RECT 3.990 79.240 1096.000 81.920 ;
        RECT 4.400 77.840 1096.000 79.240 ;
        RECT 3.990 72.440 1096.000 77.840 ;
        RECT 3.990 71.040 1095.600 72.440 ;
        RECT 3.990 68.360 1096.000 71.040 ;
        RECT 4.400 66.960 1096.000 68.360 ;
        RECT 3.990 60.880 1096.000 66.960 ;
        RECT 3.990 59.480 1095.600 60.880 ;
        RECT 3.990 58.160 1096.000 59.480 ;
        RECT 4.400 56.760 1096.000 58.160 ;
        RECT 3.990 50.000 1096.000 56.760 ;
        RECT 3.990 48.600 1095.600 50.000 ;
        RECT 3.990 47.280 1096.000 48.600 ;
        RECT 4.400 45.880 1096.000 47.280 ;
        RECT 3.990 39.120 1096.000 45.880 ;
        RECT 3.990 37.720 1095.600 39.120 ;
        RECT 3.990 37.080 1096.000 37.720 ;
        RECT 4.400 35.680 1096.000 37.080 ;
        RECT 3.990 28.240 1096.000 35.680 ;
        RECT 3.990 26.840 1095.600 28.240 ;
        RECT 3.990 26.200 1096.000 26.840 ;
        RECT 4.400 24.800 1096.000 26.200 ;
        RECT 3.990 17.360 1096.000 24.800 ;
        RECT 3.990 16.000 1095.600 17.360 ;
        RECT 4.400 15.960 1095.600 16.000 ;
        RECT 4.400 14.600 1096.000 15.960 ;
        RECT 3.990 6.480 1096.000 14.600 ;
        RECT 3.990 5.800 1095.600 6.480 ;
        RECT 4.400 5.080 1095.600 5.800 ;
        RECT 4.400 4.400 1096.000 5.080 ;
        RECT 3.990 4.255 1096.000 4.400 ;
      LAYER met4 ;
        RECT 14.095 10.640 20.640 1188.880 ;
        RECT 23.040 10.640 97.440 1188.880 ;
        RECT 99.840 10.640 1088.065 1188.880 ;
  END
END hs32_core1
END LIBRARY

