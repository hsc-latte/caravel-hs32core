magic
tech sky130A
magscale 1 2
timestamp 1608929960
<< metal1 >>
rect 170306 700884 170312 700936
rect 170364 700924 170370 700936
rect 171042 700924 171048 700936
rect 170364 700896 171048 700924
rect 170364 700884 170370 700896
rect 171042 700884 171048 700896
rect 171100 700884 171106 700936
rect 478506 700816 478512 700868
rect 478564 700856 478570 700868
rect 519078 700856 519084 700868
rect 478564 700828 519084 700856
rect 478564 700816 478570 700828
rect 519078 700816 519084 700828
rect 519136 700816 519142 700868
rect 413646 700748 413652 700800
rect 413704 700788 413710 700800
rect 519170 700788 519176 700800
rect 413704 700760 519176 700788
rect 413704 700748 413710 700760
rect 519170 700748 519176 700760
rect 519228 700748 519234 700800
rect 348786 700680 348792 700732
rect 348844 700720 348850 700732
rect 520274 700720 520280 700732
rect 348844 700692 520280 700720
rect 348844 700680 348850 700692
rect 520274 700680 520280 700692
rect 520332 700680 520338 700732
rect 283834 700612 283840 700664
rect 283892 700652 283898 700664
rect 520366 700652 520372 700664
rect 283892 700624 520372 700652
rect 283892 700612 283898 700624
rect 520366 700612 520372 700624
rect 520424 700612 520430 700664
rect 267642 700544 267648 700596
rect 267700 700584 267706 700596
rect 519262 700584 519268 700596
rect 267700 700556 519268 700584
rect 267700 700544 267706 700556
rect 519262 700544 519268 700556
rect 519320 700544 519326 700596
rect 218974 700476 218980 700528
rect 219032 700516 219038 700528
rect 519446 700516 519452 700528
rect 219032 700488 519452 700516
rect 219032 700476 219038 700488
rect 519446 700476 519452 700488
rect 519504 700476 519510 700528
rect 202782 700408 202788 700460
rect 202840 700448 202846 700460
rect 519354 700448 519360 700460
rect 202840 700420 519360 700448
rect 202840 700408 202846 700420
rect 519354 700408 519360 700420
rect 519412 700408 519418 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 154114 700340 154120 700392
rect 154172 700380 154178 700392
rect 520458 700380 520464 700392
rect 154172 700352 520464 700380
rect 154172 700340 154178 700352
rect 520458 700340 520464 700352
rect 520516 700340 520522 700392
rect 137830 700272 137836 700324
rect 137888 700312 137894 700324
rect 519538 700312 519544 700324
rect 137888 700284 519544 700312
rect 137888 700272 137894 700284
rect 519538 700272 519544 700284
rect 519596 700272 519602 700324
rect 531958 700272 531964 700324
rect 532016 700312 532022 700324
rect 559650 700312 559656 700324
rect 532016 700284 559656 700312
rect 532016 700272 532022 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 462314 700068 462320 700120
rect 462372 700108 462378 700120
rect 463602 700108 463608 700120
rect 462372 700080 463608 700108
rect 462372 700068 462378 700080
rect 463602 700068 463608 700080
rect 463660 700068 463666 700120
rect 397454 699932 397460 699984
rect 397512 699972 397518 699984
rect 398742 699972 398748 699984
rect 397512 699944 398748 699972
rect 397512 699932 397518 699944
rect 398742 699932 398748 699944
rect 398800 699932 398806 699984
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300578 699700 300584 699712
rect 300176 699672 300584 699700
rect 300176 699660 300182 699672
rect 300578 699660 300584 699672
rect 300636 699660 300642 699712
rect 364978 699660 364984 699712
rect 365036 699700 365042 699712
rect 365622 699700 365628 699712
rect 365036 699672 365628 699700
rect 365036 699660 365042 699672
rect 365622 699660 365628 699672
rect 365680 699660 365686 699712
rect 429838 699660 429844 699712
rect 429896 699700 429902 699712
rect 430482 699700 430488 699712
rect 429896 699672 430488 699700
rect 429896 699660 429902 699672
rect 430482 699660 430488 699672
rect 430540 699660 430546 699712
rect 494790 699660 494796 699712
rect 494848 699700 494854 699712
rect 495342 699700 495348 699712
rect 494848 699672 495348 699700
rect 494848 699660 494854 699672
rect 495342 699660 495348 699672
rect 495400 699660 495406 699712
rect 542722 698232 542728 698284
rect 542780 698272 542786 698284
rect 543550 698272 543556 698284
rect 542780 698244 543556 698272
rect 542780 698232 542786 698244
rect 543550 698232 543556 698244
rect 543608 698232 543614 698284
rect 545758 696940 545764 696992
rect 545816 696980 545822 696992
rect 580166 696980 580172 696992
rect 545816 696952 580172 696980
rect 545816 696940 545822 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 542538 694084 542544 694136
rect 542596 694124 542602 694136
rect 542722 694124 542728 694136
rect 542596 694096 542728 694124
rect 542596 694084 542602 694096
rect 542722 694084 542728 694096
rect 542780 694084 542786 694136
rect 560938 685856 560944 685908
rect 560996 685896 561002 685908
rect 580166 685896 580172 685908
rect 560996 685868 580172 685896
rect 560996 685856 561002 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 542446 684496 542452 684548
rect 542504 684536 542510 684548
rect 542538 684536 542544 684548
rect 542504 684508 542544 684536
rect 542504 684496 542510 684508
rect 542538 684496 542544 684508
rect 542596 684496 542602 684548
rect 529198 673480 529204 673532
rect 529256 673520 529262 673532
rect 580166 673520 580172 673532
rect 529256 673492 580172 673520
rect 529256 673480 529262 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 542538 666544 542544 666596
rect 542596 666584 542602 666596
rect 542814 666584 542820 666596
rect 542596 666556 542820 666584
rect 542596 666544 542602 666556
rect 542814 666544 542820 666556
rect 542872 666544 542878 666596
rect 542538 661716 542544 661768
rect 542596 661756 542602 661768
rect 542814 661756 542820 661768
rect 542596 661728 542820 661756
rect 542596 661716 542602 661728
rect 542814 661716 542820 661728
rect 542872 661716 542878 661768
rect 542538 656888 542544 656940
rect 542596 656928 542602 656940
rect 542630 656928 542636 656940
rect 542596 656900 542636 656928
rect 542596 656888 542602 656900
rect 542630 656888 542636 656900
rect 542688 656888 542694 656940
rect 540238 650020 540244 650072
rect 540296 650060 540302 650072
rect 580166 650060 580172 650072
rect 540296 650032 580172 650060
rect 540296 650020 540302 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 542538 647232 542544 647284
rect 542596 647272 542602 647284
rect 542630 647272 542636 647284
rect 542596 647244 542636 647272
rect 542596 647232 542602 647244
rect 542630 647232 542636 647244
rect 542688 647232 542694 647284
rect 542538 640364 542544 640416
rect 542596 640404 542602 640416
rect 542630 640404 542636 640416
rect 542596 640376 542636 640404
rect 542596 640364 542602 640376
rect 542630 640364 542636 640376
rect 542688 640364 542694 640416
rect 558178 638936 558184 638988
rect 558236 638976 558242 638988
rect 580166 638976 580172 638988
rect 558236 638948 580172 638976
rect 558236 638936 558242 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 542446 630640 542452 630692
rect 542504 630680 542510 630692
rect 542630 630680 542636 630692
rect 542504 630652 542636 630680
rect 542504 630640 542510 630652
rect 542630 630640 542636 630652
rect 542688 630640 542694 630692
rect 525058 626560 525064 626612
rect 525116 626600 525122 626612
rect 580166 626600 580172 626612
rect 525116 626572 580172 626600
rect 525116 626560 525122 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 488534 613368 488540 613420
rect 488592 613408 488598 613420
rect 493962 613408 493968 613420
rect 488592 613380 493968 613408
rect 488592 613368 488598 613380
rect 493962 613368 493968 613380
rect 494020 613368 494026 613420
rect 373626 612756 373632 612808
rect 373684 612796 373690 612808
rect 379606 612796 379612 612808
rect 373684 612768 379612 612796
rect 373684 612756 373690 612768
rect 379606 612756 379612 612768
rect 379664 612796 379670 612808
rect 488534 612796 488540 612808
rect 379664 612768 488540 612796
rect 379664 612756 379670 612768
rect 488534 612756 488540 612768
rect 488592 612756 488598 612808
rect 493962 612756 493968 612808
rect 494020 612796 494026 612808
rect 499574 612796 499580 612808
rect 494020 612768 499580 612796
rect 494020 612756 494026 612768
rect 499574 612756 499580 612768
rect 499632 612756 499638 612808
rect 542446 611328 542452 611380
rect 542504 611368 542510 611380
rect 542630 611368 542636 611380
rect 542504 611340 542636 611368
rect 542504 611328 542510 611340
rect 542630 611328 542636 611340
rect 542688 611328 542694 611380
rect 495342 610852 495348 610904
rect 495400 610892 495406 610904
rect 520550 610892 520556 610904
rect 495400 610864 520556 610892
rect 495400 610852 495406 610864
rect 520550 610852 520556 610864
rect 520608 610852 520614 610904
rect 463602 610784 463608 610836
rect 463660 610824 463666 610836
rect 519630 610824 519636 610836
rect 463660 610796 519636 610824
rect 463660 610784 463666 610796
rect 519630 610784 519636 610796
rect 519688 610784 519694 610836
rect 430482 610716 430488 610768
rect 430540 610756 430546 610768
rect 520642 610756 520648 610768
rect 430540 610728 520648 610756
rect 430540 610716 430546 610728
rect 520642 610716 520648 610728
rect 520700 610716 520706 610768
rect 365622 610648 365628 610700
rect 365680 610688 365686 610700
rect 520734 610688 520740 610700
rect 365680 610660 520740 610688
rect 365680 610648 365686 610660
rect 520734 610648 520740 610660
rect 520792 610648 520798 610700
rect 332502 610580 332508 610632
rect 332560 610620 332566 610632
rect 519722 610620 519728 610632
rect 332560 610592 519728 610620
rect 332560 610580 332566 610592
rect 519722 610580 519728 610592
rect 519780 610580 519786 610632
rect 379974 610376 379980 610428
rect 380032 610416 380038 610428
rect 496446 610416 496452 610428
rect 380032 610388 496452 610416
rect 380032 610376 380038 610388
rect 496446 610376 496452 610388
rect 496504 610376 496510 610428
rect 3418 610308 3424 610360
rect 3476 610348 3482 610360
rect 520826 610348 520832 610360
rect 3476 610320 520832 610348
rect 3476 610308 3482 610320
rect 520826 610308 520832 610320
rect 520884 610308 520890 610360
rect 542446 608540 542452 608592
rect 542504 608580 542510 608592
rect 542538 608580 542544 608592
rect 542504 608552 542544 608580
rect 542504 608540 542510 608552
rect 542538 608540 542544 608552
rect 542596 608540 542602 608592
rect 389082 605820 389088 605872
rect 389140 605860 389146 605872
rect 416774 605860 416780 605872
rect 389140 605832 416780 605860
rect 389140 605820 389146 605832
rect 416774 605820 416780 605832
rect 416832 605820 416838 605872
rect 387702 604460 387708 604512
rect 387760 604500 387766 604512
rect 416774 604500 416780 604512
rect 387760 604472 416780 604500
rect 387760 604460 387766 604472
rect 416774 604460 416780 604472
rect 416832 604460 416838 604512
rect 384942 603100 384948 603152
rect 385000 603140 385006 603152
rect 416774 603140 416780 603152
rect 385000 603112 416780 603140
rect 385000 603100 385006 603112
rect 416774 603100 416780 603112
rect 416832 603100 416838 603152
rect 538858 603100 538864 603152
rect 538916 603140 538922 603152
rect 580166 603140 580172 603152
rect 538916 603112 580172 603140
rect 538916 603100 538922 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 383562 601672 383568 601724
rect 383620 601712 383626 601724
rect 416774 601712 416780 601724
rect 383620 601684 416780 601712
rect 383620 601672 383626 601684
rect 416774 601672 416780 601684
rect 416832 601672 416838 601724
rect 542446 601672 542452 601724
rect 542504 601712 542510 601724
rect 542722 601712 542728 601724
rect 542504 601684 542728 601712
rect 542504 601672 542510 601684
rect 542722 601672 542728 601684
rect 542780 601672 542786 601724
rect 380802 600312 380808 600364
rect 380860 600352 380866 600364
rect 416774 600352 416780 600364
rect 380860 600324 416780 600352
rect 380860 600312 380866 600324
rect 416774 600312 416780 600324
rect 416832 600312 416838 600364
rect 378042 598952 378048 599004
rect 378100 598992 378106 599004
rect 416774 598992 416780 599004
rect 378100 598964 416780 598992
rect 378100 598952 378106 598964
rect 416774 598952 416780 598964
rect 416832 598952 416838 599004
rect 542538 598884 542544 598936
rect 542596 598924 542602 598936
rect 542722 598924 542728 598936
rect 542596 598896 542728 598924
rect 542596 598884 542602 598896
rect 542722 598884 542728 598896
rect 542780 598884 542786 598936
rect 410518 597524 410524 597576
rect 410576 597564 410582 597576
rect 416774 597564 416780 597576
rect 410576 597536 416780 597564
rect 410576 597524 410582 597536
rect 416774 597524 416780 597536
rect 416832 597524 416838 597576
rect 556798 592016 556804 592068
rect 556856 592056 556862 592068
rect 580166 592056 580172 592068
rect 556856 592028 580172 592056
rect 556856 592016 556862 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 542538 589296 542544 589348
rect 542596 589336 542602 589348
rect 542814 589336 542820 589348
rect 542596 589308 542820 589336
rect 542596 589296 542602 589308
rect 542814 589296 542820 589308
rect 542872 589296 542878 589348
rect 542814 582468 542820 582480
rect 542740 582440 542820 582468
rect 542740 582344 542768 582440
rect 542814 582428 542820 582440
rect 542872 582428 542878 582480
rect 542722 582292 542728 582344
rect 542780 582292 542786 582344
rect 523678 579640 523684 579692
rect 523736 579680 523742 579692
rect 580166 579680 580172 579692
rect 523736 579652 580172 579680
rect 523736 579640 523742 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 542446 563116 542452 563168
rect 542504 563116 542510 563168
rect 542464 563032 542492 563116
rect 542446 562980 542452 563032
rect 542504 562980 542510 563032
rect 537478 556180 537484 556232
rect 537536 556220 537542 556232
rect 580166 556220 580172 556232
rect 537536 556192 580172 556220
rect 537536 556180 537542 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 542354 553392 542360 553444
rect 542412 553432 542418 553444
rect 542412 553404 542492 553432
rect 542412 553392 542418 553404
rect 542464 553376 542492 553404
rect 542446 553324 542452 553376
rect 542504 553324 542510 553376
rect 542354 550604 542360 550656
rect 542412 550644 542418 550656
rect 542446 550644 542452 550656
rect 542412 550616 542452 550644
rect 542412 550604 542418 550616
rect 542446 550604 542452 550616
rect 542504 550604 542510 550656
rect 555418 545096 555424 545148
rect 555476 545136 555482 545148
rect 580166 545136 580172 545148
rect 555476 545108 580172 545136
rect 555476 545096 555482 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 542354 543736 542360 543788
rect 542412 543736 542418 543788
rect 542372 543640 542400 543736
rect 542446 543640 542452 543652
rect 542372 543612 542452 543640
rect 542446 543600 542452 543612
rect 542504 543600 542510 543652
rect 411162 539588 411168 539640
rect 411220 539628 411226 539640
rect 416774 539628 416780 539640
rect 411220 539600 416780 539628
rect 411220 539588 411226 539600
rect 416774 539588 416780 539600
rect 416832 539588 416838 539640
rect 379514 538228 379520 538280
rect 379572 538268 379578 538280
rect 379790 538268 379796 538280
rect 379572 538240 379796 538268
rect 379572 538228 379578 538240
rect 379790 538228 379796 538240
rect 379848 538228 379854 538280
rect 409138 538228 409144 538280
rect 409196 538268 409202 538280
rect 416774 538268 416780 538280
rect 409196 538240 416780 538268
rect 409196 538228 409202 538240
rect 416774 538228 416780 538240
rect 416832 538228 416838 538280
rect 379514 536052 379520 536104
rect 379572 536092 379578 536104
rect 379790 536092 379796 536104
rect 379572 536064 379796 536092
rect 379572 536052 379578 536064
rect 379790 536052 379796 536064
rect 379848 536052 379854 536104
rect 542446 534012 542452 534064
rect 542504 534052 542510 534064
rect 542630 534052 542636 534064
rect 542504 534024 542636 534052
rect 542504 534012 542510 534024
rect 542630 534012 542636 534024
rect 542688 534012 542694 534064
rect 523770 532720 523776 532772
rect 523828 532760 523834 532772
rect 580166 532760 580172 532772
rect 523828 532732 580172 532760
rect 523828 532720 523834 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 542630 524424 542636 524476
rect 542688 524424 542694 524476
rect 542648 524396 542676 524424
rect 542722 524396 542728 524408
rect 542648 524368 542728 524396
rect 542722 524356 542728 524368
rect 542780 524356 542786 524408
rect 408494 521568 408500 521620
rect 408552 521608 408558 521620
rect 409138 521608 409144 521620
rect 408552 521580 409144 521608
rect 408552 521568 408558 521580
rect 409138 521568 409144 521580
rect 409196 521568 409202 521620
rect 297266 520888 297272 520940
rect 297324 520928 297330 520940
rect 408494 520928 408500 520940
rect 297324 520900 408500 520928
rect 297324 520888 297330 520900
rect 408494 520888 408500 520900
rect 408552 520888 408558 520940
rect 379606 519528 379612 519580
rect 379664 519568 379670 519580
rect 379790 519568 379796 519580
rect 379664 519540 379796 519568
rect 379664 519528 379670 519540
rect 379790 519528 379796 519540
rect 379848 519528 379854 519580
rect 318702 518848 318708 518900
rect 318760 518888 318766 518900
rect 327166 518888 327172 518900
rect 318760 518860 327172 518888
rect 318760 518848 318766 518860
rect 327166 518848 327172 518860
rect 327224 518848 327230 518900
rect 317322 518780 317328 518832
rect 317380 518820 317386 518832
rect 325418 518820 325424 518832
rect 317380 518792 325424 518820
rect 317380 518780 317386 518792
rect 325418 518780 325424 518792
rect 325476 518780 325482 518832
rect 331214 518780 331220 518832
rect 331272 518820 331278 518832
rect 340506 518820 340512 518832
rect 331272 518792 340512 518820
rect 331272 518780 331278 518792
rect 340506 518780 340512 518792
rect 340564 518780 340570 518832
rect 369854 518780 369860 518832
rect 369912 518820 369918 518832
rect 379422 518820 379428 518832
rect 369912 518792 379428 518820
rect 369912 518780 369918 518792
rect 379422 518780 379428 518792
rect 379480 518780 379486 518832
rect 379514 518780 379520 518832
rect 379572 518820 379578 518832
rect 388990 518820 388996 518832
rect 379572 518792 388996 518820
rect 379572 518780 379578 518792
rect 388990 518780 388996 518792
rect 389048 518780 389054 518832
rect 393314 518780 393320 518832
rect 393372 518820 393378 518832
rect 402882 518820 402888 518832
rect 393372 518792 402888 518820
rect 393372 518780 393378 518792
rect 402882 518780 402888 518792
rect 402940 518780 402946 518832
rect 451274 518780 451280 518832
rect 451332 518820 451338 518832
rect 459554 518820 459560 518832
rect 451332 518792 459560 518820
rect 451332 518780 451338 518792
rect 459554 518780 459560 518792
rect 459612 518780 459618 518832
rect 307570 518712 307576 518764
rect 307628 518752 307634 518764
rect 324314 518752 324320 518764
rect 307628 518724 324320 518752
rect 307628 518712 307634 518724
rect 324314 518712 324320 518724
rect 324372 518712 324378 518764
rect 326430 518712 326436 518764
rect 326488 518752 326494 518764
rect 335538 518752 335544 518764
rect 326488 518724 335544 518752
rect 326488 518712 326494 518724
rect 335538 518712 335544 518724
rect 335596 518752 335602 518764
rect 345474 518752 345480 518764
rect 335596 518724 345480 518752
rect 335596 518712 335602 518724
rect 345474 518712 345480 518724
rect 345532 518752 345538 518764
rect 441614 518752 441620 518764
rect 345532 518724 441620 518752
rect 345532 518712 345538 518724
rect 441614 518712 441620 518724
rect 441672 518712 441678 518764
rect 443178 518712 443184 518764
rect 443236 518752 443242 518764
rect 452562 518752 452568 518764
rect 443236 518724 452568 518752
rect 443236 518712 443242 518724
rect 452562 518712 452568 518724
rect 452620 518752 452626 518764
rect 460934 518752 460940 518764
rect 452620 518724 460940 518752
rect 452620 518712 452626 518724
rect 460934 518712 460940 518724
rect 460992 518712 460998 518764
rect 314562 518644 314568 518696
rect 314620 518684 314626 518696
rect 323118 518684 323124 518696
rect 314620 518656 323124 518684
rect 314620 518644 314626 518656
rect 323118 518644 323124 518656
rect 323176 518684 323182 518696
rect 332318 518684 332324 518696
rect 323176 518656 332324 518684
rect 323176 518644 323182 518656
rect 332318 518644 332324 518656
rect 332376 518684 332382 518696
rect 332376 518656 337148 518684
rect 332376 518644 332382 518656
rect 320082 518576 320088 518628
rect 320140 518616 320146 518628
rect 328914 518616 328920 518628
rect 320140 518588 328920 518616
rect 320140 518576 320146 518588
rect 328914 518576 328920 518588
rect 328972 518616 328978 518628
rect 337120 518616 337148 518656
rect 337194 518644 337200 518696
rect 337252 518684 337258 518696
rect 346486 518684 346492 518696
rect 337252 518656 346492 518684
rect 337252 518644 337258 518656
rect 346486 518644 346492 518656
rect 346544 518684 346550 518696
rect 442994 518684 443000 518696
rect 346544 518656 443000 518684
rect 346544 518644 346550 518656
rect 442994 518644 443000 518656
rect 443052 518644 443058 518696
rect 453666 518644 453672 518696
rect 453724 518684 453730 518696
rect 462314 518684 462320 518696
rect 453724 518656 462320 518684
rect 453724 518644 453730 518656
rect 462314 518644 462320 518656
rect 462372 518644 462378 518696
rect 341610 518616 341616 518628
rect 328972 518588 337056 518616
rect 337120 518588 341616 518616
rect 328972 518576 328978 518588
rect 317322 518508 317328 518560
rect 317380 518548 317386 518560
rect 326430 518548 326436 518560
rect 317380 518520 326436 518548
rect 317380 518508 317386 518520
rect 326430 518508 326436 518520
rect 326488 518508 326494 518560
rect 327166 518508 327172 518560
rect 327224 518548 327230 518560
rect 336642 518548 336648 518560
rect 327224 518520 336648 518548
rect 327224 518508 327230 518520
rect 336642 518508 336648 518520
rect 336700 518508 336706 518560
rect 337028 518548 337056 518588
rect 341610 518576 341616 518588
rect 341668 518616 341674 518628
rect 342162 518616 342168 518628
rect 341668 518588 342168 518616
rect 341668 518576 341674 518588
rect 342162 518576 342168 518588
rect 342220 518576 342226 518628
rect 347774 518576 347780 518628
rect 347832 518616 347838 518628
rect 348602 518616 348608 518628
rect 347832 518588 348608 518616
rect 347832 518576 347838 518588
rect 348602 518576 348608 518588
rect 348660 518616 348666 518628
rect 350534 518616 350540 518628
rect 348660 518588 350540 518616
rect 348660 518576 348666 518588
rect 350534 518576 350540 518588
rect 350592 518576 350598 518628
rect 357434 518576 357440 518628
rect 357492 518616 357498 518628
rect 362218 518616 362224 518628
rect 357492 518588 362224 518616
rect 357492 518576 357498 518588
rect 362218 518576 362224 518588
rect 362276 518576 362282 518628
rect 379422 518576 379428 518628
rect 379480 518616 379486 518628
rect 379514 518616 379520 518628
rect 379480 518588 379520 518616
rect 379480 518576 379486 518588
rect 379514 518576 379520 518588
rect 379572 518576 379578 518628
rect 402882 518576 402888 518628
rect 402940 518616 402946 518628
rect 432506 518616 432512 518628
rect 402940 518588 432512 518616
rect 402940 518576 402946 518588
rect 432506 518576 432512 518588
rect 432564 518576 432570 518628
rect 446582 518576 446588 518628
rect 446640 518616 446646 518628
rect 456058 518616 456064 518628
rect 446640 518588 456064 518616
rect 446640 518576 446646 518588
rect 456058 518576 456064 518588
rect 456116 518616 456122 518628
rect 465074 518616 465080 518628
rect 456116 518588 465080 518616
rect 456116 518576 456122 518588
rect 465074 518576 465080 518588
rect 465132 518576 465138 518628
rect 338114 518548 338120 518560
rect 337028 518520 338120 518548
rect 338114 518508 338120 518520
rect 338172 518548 338178 518560
rect 347682 518548 347688 518560
rect 338172 518520 347688 518548
rect 338172 518508 338178 518520
rect 347682 518508 347688 518520
rect 347740 518548 347746 518560
rect 445754 518548 445760 518560
rect 347740 518520 445760 518548
rect 347740 518508 347746 518520
rect 445754 518508 445760 518520
rect 445812 518508 445818 518560
rect 447410 518508 447416 518560
rect 447468 518548 447474 518560
rect 456886 518548 456892 518560
rect 447468 518520 456892 518548
rect 447468 518508 447474 518520
rect 456886 518508 456892 518520
rect 456944 518508 456950 518560
rect 315942 518440 315948 518492
rect 316000 518480 316006 518492
rect 324406 518480 324412 518492
rect 316000 518452 324412 518480
rect 316000 518440 316006 518452
rect 324406 518440 324412 518452
rect 324464 518480 324470 518492
rect 324464 518452 325372 518480
rect 324464 518440 324470 518452
rect 292482 518372 292488 518424
rect 292540 518412 292546 518424
rect 316034 518412 316040 518424
rect 292540 518384 316040 518412
rect 292540 518372 292546 518384
rect 316034 518372 316040 518384
rect 316092 518372 316098 518424
rect 325344 518412 325372 518452
rect 325418 518440 325424 518492
rect 325476 518480 325482 518492
rect 334158 518480 334164 518492
rect 325476 518452 334164 518480
rect 325476 518440 325482 518452
rect 334158 518440 334164 518452
rect 334216 518480 334222 518492
rect 335170 518480 335176 518492
rect 334216 518452 335176 518480
rect 334216 518440 334222 518452
rect 335170 518440 335176 518452
rect 335228 518440 335234 518492
rect 362218 518440 362224 518492
rect 362276 518480 362282 518492
rect 369854 518480 369860 518492
rect 362276 518452 369860 518480
rect 362276 518440 362282 518452
rect 369854 518440 369860 518452
rect 369912 518440 369918 518492
rect 388990 518440 388996 518492
rect 389048 518480 389054 518492
rect 393314 518480 393320 518492
rect 389048 518452 393320 518480
rect 389048 518440 389054 518452
rect 393314 518440 393320 518452
rect 393372 518440 393378 518492
rect 448790 518440 448796 518492
rect 448848 518480 448854 518492
rect 458266 518480 458272 518492
rect 448848 518452 458272 518480
rect 448848 518440 448854 518452
rect 458266 518440 458272 518452
rect 458324 518480 458330 518492
rect 466546 518480 466552 518492
rect 458324 518452 466552 518480
rect 458324 518440 458330 518452
rect 466546 518440 466552 518452
rect 466604 518440 466610 518492
rect 333422 518412 333428 518424
rect 325344 518384 333428 518412
rect 333422 518372 333428 518384
rect 333480 518412 333486 518424
rect 342990 518412 342996 518424
rect 333480 518384 342996 518412
rect 333480 518372 333486 518384
rect 342990 518372 342996 518384
rect 343048 518412 343054 518424
rect 343542 518412 343548 518424
rect 343048 518384 343548 518412
rect 343048 518372 343054 518384
rect 343542 518372 343548 518384
rect 343600 518372 343606 518424
rect 350534 518372 350540 518424
rect 350592 518412 350598 518424
rect 357434 518412 357440 518424
rect 350592 518384 357440 518412
rect 350592 518372 350598 518384
rect 357434 518372 357440 518384
rect 357492 518372 357498 518424
rect 373902 518372 373908 518424
rect 373960 518412 373966 518424
rect 426434 518412 426440 518424
rect 373960 518384 426440 518412
rect 373960 518372 373966 518384
rect 426434 518372 426440 518384
rect 426492 518372 426498 518424
rect 445386 518372 445392 518424
rect 445444 518412 445450 518424
rect 455322 518412 455328 518424
rect 445444 518384 455328 518412
rect 445444 518372 445450 518384
rect 455322 518372 455328 518384
rect 455380 518372 455386 518424
rect 456886 518372 456892 518424
rect 456944 518412 456950 518424
rect 466454 518412 466460 518424
rect 456944 518384 466460 518412
rect 456944 518372 456950 518384
rect 466454 518372 466460 518384
rect 466512 518372 466518 518424
rect 295242 518304 295248 518356
rect 295300 518344 295306 518356
rect 317414 518344 317420 518356
rect 295300 518316 317420 518344
rect 295300 518304 295306 518316
rect 317414 518304 317420 518316
rect 317472 518304 317478 518356
rect 321094 518304 321100 518356
rect 321152 518344 321158 518356
rect 330110 518344 330116 518356
rect 321152 518316 330116 518344
rect 321152 518304 321158 518316
rect 330110 518304 330116 518316
rect 330168 518344 330174 518356
rect 339954 518344 339960 518356
rect 330168 518316 339960 518344
rect 330168 518304 330174 518316
rect 339954 518304 339960 518316
rect 340012 518344 340018 518356
rect 347774 518344 347780 518356
rect 340012 518316 347780 518344
rect 340012 518304 340018 518316
rect 347774 518304 347780 518316
rect 347832 518304 347838 518356
rect 362862 518304 362868 518356
rect 362920 518344 362926 518356
rect 430574 518344 430580 518356
rect 362920 518316 430580 518344
rect 362920 518304 362926 518316
rect 430574 518304 430580 518316
rect 430632 518304 430638 518356
rect 432506 518304 432512 518356
rect 432564 518344 432570 518356
rect 447134 518344 447140 518356
rect 432564 518316 447140 518344
rect 432564 518304 432570 518316
rect 447134 518304 447140 518316
rect 447192 518304 447198 518356
rect 449894 518304 449900 518356
rect 449952 518344 449958 518356
rect 459554 518344 459560 518356
rect 449952 518316 459560 518344
rect 449952 518304 449958 518316
rect 459554 518304 459560 518316
rect 459612 518344 459618 518356
rect 467834 518344 467840 518356
rect 459612 518316 467840 518344
rect 459612 518304 459618 518316
rect 467834 518304 467840 518316
rect 467892 518304 467898 518356
rect 313182 518236 313188 518288
rect 313240 518276 313246 518288
rect 321738 518276 321744 518288
rect 313240 518248 321744 518276
rect 313240 518236 313246 518248
rect 321738 518236 321744 518248
rect 321796 518276 321802 518288
rect 331214 518276 331220 518288
rect 321796 518248 331220 518276
rect 321796 518236 321802 518248
rect 331214 518236 331220 518248
rect 331272 518236 331278 518288
rect 335170 518236 335176 518288
rect 335228 518276 335234 518288
rect 344186 518276 344192 518288
rect 335228 518248 344192 518276
rect 335228 518236 335234 518248
rect 344186 518236 344192 518248
rect 344244 518276 344250 518288
rect 344922 518276 344928 518288
rect 344244 518248 344928 518276
rect 344244 518236 344250 518248
rect 344922 518236 344928 518248
rect 344980 518236 344986 518288
rect 361482 518236 361488 518288
rect 361540 518276 361546 518288
rect 429286 518276 429292 518288
rect 361540 518248 429292 518276
rect 361540 518236 361546 518248
rect 429286 518236 429292 518248
rect 429344 518236 429350 518288
rect 432598 518236 432604 518288
rect 432656 518276 432662 518288
rect 442074 518276 442080 518288
rect 432656 518248 442080 518276
rect 432656 518236 432662 518248
rect 442074 518236 442080 518248
rect 442132 518276 442138 518288
rect 442132 518248 442212 518276
rect 442132 518236 442138 518248
rect 303614 518168 303620 518220
rect 303672 518208 303678 518220
rect 423674 518208 423680 518220
rect 303672 518180 423680 518208
rect 303672 518168 303678 518180
rect 423674 518168 423680 518180
rect 423732 518168 423738 518220
rect 442184 518208 442212 518248
rect 444282 518236 444288 518288
rect 444340 518276 444346 518288
rect 453666 518276 453672 518288
rect 444340 518248 453672 518276
rect 444340 518236 444346 518248
rect 453666 518236 453672 518248
rect 453724 518236 453730 518288
rect 455322 518236 455328 518288
rect 455380 518276 455386 518288
rect 463694 518276 463700 518288
rect 455380 518248 463700 518276
rect 455380 518236 455386 518248
rect 463694 518236 463700 518248
rect 463752 518236 463758 518288
rect 451274 518208 451280 518220
rect 442184 518180 451280 518208
rect 451274 518168 451280 518180
rect 451332 518168 451338 518220
rect 306282 518100 306288 518152
rect 306340 518140 306346 518152
rect 322934 518140 322940 518152
rect 306340 518112 322940 518140
rect 306340 518100 306346 518112
rect 322934 518100 322940 518112
rect 322992 518100 322998 518152
rect 358722 518100 358728 518152
rect 358780 518140 358786 518152
rect 429194 518140 429200 518152
rect 358780 518112 429200 518140
rect 358780 518100 358786 518112
rect 429194 518100 429200 518112
rect 429252 518100 429258 518152
rect 303522 518032 303528 518084
rect 303580 518072 303586 518084
rect 321830 518072 321836 518084
rect 303580 518044 321836 518072
rect 303580 518032 303586 518044
rect 321830 518032 321836 518044
rect 321888 518032 321894 518084
rect 355962 518032 355968 518084
rect 356020 518072 356026 518084
rect 425606 518072 425612 518084
rect 356020 518044 425612 518072
rect 356020 518032 356026 518044
rect 425606 518032 425612 518044
rect 425664 518032 425670 518084
rect 435910 518032 435916 518084
rect 435968 518072 435974 518084
rect 444282 518072 444288 518084
rect 435968 518044 444288 518072
rect 435968 518032 435974 518044
rect 444282 518032 444288 518044
rect 444340 518032 444346 518084
rect 299382 517964 299388 518016
rect 299440 518004 299446 518016
rect 318794 518004 318800 518016
rect 299440 517976 318800 518004
rect 299440 517964 299446 517976
rect 318794 517964 318800 517976
rect 318852 517964 318858 518016
rect 327074 518004 327080 518016
rect 323412 517976 327080 518004
rect 296622 517896 296628 517948
rect 296680 517936 296686 517948
rect 317506 517936 317512 517948
rect 296680 517908 317512 517936
rect 296680 517896 296686 517908
rect 317506 517896 317512 517908
rect 317564 517896 317570 517948
rect 285582 517828 285588 517880
rect 285640 517868 285646 517880
rect 312078 517868 312084 517880
rect 285640 517840 312084 517868
rect 285640 517828 285646 517840
rect 312078 517828 312084 517840
rect 312136 517828 312142 517880
rect 314562 517828 314568 517880
rect 314620 517868 314626 517880
rect 323412 517868 323440 517976
rect 327074 517964 327080 517976
rect 327132 517964 327138 518016
rect 340506 517964 340512 518016
rect 340564 518004 340570 518016
rect 431954 518004 431960 518016
rect 340564 517976 431960 518004
rect 340564 517964 340570 517976
rect 431954 517964 431960 517976
rect 432012 517964 432018 518016
rect 331214 517936 331220 517948
rect 314620 517840 323440 517868
rect 326356 517908 331220 517936
rect 314620 517828 314626 517840
rect 300670 517760 300676 517812
rect 300728 517800 300734 517812
rect 320174 517800 320180 517812
rect 300728 517772 320180 517800
rect 300728 517760 300734 517772
rect 320174 517760 320180 517772
rect 320232 517760 320238 517812
rect 321462 517760 321468 517812
rect 321520 517800 321526 517812
rect 326356 517800 326384 517908
rect 331214 517896 331220 517908
rect 331272 517896 331278 517948
rect 343542 517896 343548 517948
rect 343600 517936 343606 517948
rect 436094 517936 436100 517948
rect 343600 517908 436100 517936
rect 343600 517896 343606 517908
rect 436094 517896 436100 517908
rect 436152 517896 436158 517948
rect 436738 517896 436744 517948
rect 436796 517936 436802 517948
rect 437290 517936 437296 517948
rect 436796 517908 437296 517936
rect 436796 517896 436802 517908
rect 437290 517896 437296 517908
rect 437348 517936 437354 517948
rect 446582 517936 446588 517948
rect 437348 517908 446588 517936
rect 437348 517896 437354 517908
rect 446582 517896 446588 517908
rect 446640 517896 446646 517948
rect 332594 517868 332600 517880
rect 321520 517772 326384 517800
rect 326448 517840 332600 517868
rect 321520 517760 321526 517772
rect 280890 517692 280896 517744
rect 280948 517732 280954 517744
rect 303614 517732 303620 517744
rect 280948 517704 303620 517732
rect 280948 517692 280954 517704
rect 303614 517692 303620 517704
rect 303672 517692 303678 517744
rect 310422 517692 310428 517744
rect 310480 517732 310486 517744
rect 310480 517704 322796 517732
rect 310480 517692 310486 517704
rect 288342 517624 288348 517676
rect 288400 517664 288406 517676
rect 313274 517664 313280 517676
rect 288400 517636 313280 517664
rect 288400 517624 288406 517636
rect 313274 517624 313280 517636
rect 313332 517624 313338 517676
rect 322768 517664 322796 517704
rect 322842 517692 322848 517744
rect 322900 517732 322906 517744
rect 326448 517732 326476 517840
rect 332594 517828 332600 517840
rect 332652 517828 332658 517880
rect 433886 517828 433892 517880
rect 433944 517868 433950 517880
rect 443178 517868 443184 517880
rect 433944 517840 443184 517868
rect 433944 517828 433950 517840
rect 443178 517828 443184 517840
rect 443236 517828 443242 517880
rect 438118 517760 438124 517812
rect 438176 517800 438182 517812
rect 447410 517800 447416 517812
rect 438176 517772 447416 517800
rect 438176 517760 438182 517772
rect 447410 517760 447416 517772
rect 447468 517760 447474 517812
rect 322900 517704 326476 517732
rect 322900 517692 322906 517704
rect 328362 517692 328368 517744
rect 328420 517732 328426 517744
rect 333974 517732 333980 517744
rect 328420 517704 333980 517732
rect 328420 517692 328426 517704
rect 333974 517692 333980 517704
rect 334032 517692 334038 517744
rect 440878 517692 440884 517744
rect 440936 517732 440942 517744
rect 449894 517732 449900 517744
rect 440936 517704 449900 517732
rect 440936 517692 440942 517704
rect 449894 517692 449900 517704
rect 449952 517692 449958 517744
rect 324314 517664 324320 517676
rect 322768 517636 324320 517664
rect 324314 517624 324320 517636
rect 324372 517624 324378 517676
rect 326338 517624 326344 517676
rect 326396 517664 326402 517676
rect 329834 517664 329840 517676
rect 326396 517636 329840 517664
rect 326396 517624 326402 517636
rect 329834 517624 329840 517636
rect 329892 517624 329898 517676
rect 330478 517624 330484 517676
rect 330536 517664 330542 517676
rect 335722 517664 335728 517676
rect 330536 517636 335728 517664
rect 330536 517624 330542 517636
rect 335722 517624 335728 517636
rect 335780 517624 335786 517676
rect 344922 517624 344928 517676
rect 344980 517664 344986 517676
rect 438854 517664 438860 517676
rect 344980 517636 438860 517664
rect 344980 517624 344986 517636
rect 438854 517624 438860 517636
rect 438912 517624 438918 517676
rect 439498 517624 439504 517676
rect 439556 517664 439562 517676
rect 448790 517664 448796 517676
rect 439556 517636 448796 517664
rect 439556 517624 439562 517636
rect 448790 517624 448796 517636
rect 448848 517624 448854 517676
rect 289722 517556 289728 517608
rect 289780 517596 289786 517608
rect 314654 517596 314660 517608
rect 289780 517568 314660 517596
rect 289780 517556 289786 517568
rect 314654 517556 314660 517568
rect 314712 517556 314718 517608
rect 317322 517556 317328 517608
rect 317380 517596 317386 517608
rect 317380 517568 325832 517596
rect 317380 517556 317386 517568
rect 311802 517488 311808 517540
rect 311860 517528 311866 517540
rect 325694 517528 325700 517540
rect 311860 517500 325700 517528
rect 311860 517488 311866 517500
rect 325694 517488 325700 517500
rect 325752 517488 325758 517540
rect 325804 517528 325832 517568
rect 327718 517556 327724 517608
rect 327776 517596 327782 517608
rect 332594 517596 332600 517608
rect 327776 517568 332600 517596
rect 327776 517556 327782 517568
rect 332594 517556 332600 517568
rect 332652 517556 332658 517608
rect 333882 517556 333888 517608
rect 333940 517596 333946 517608
rect 338114 517596 338120 517608
rect 333940 517568 338120 517596
rect 333940 517556 333946 517568
rect 338114 517556 338120 517568
rect 338172 517556 338178 517608
rect 342162 517556 342168 517608
rect 342220 517596 342226 517608
rect 434714 517596 434720 517608
rect 342220 517568 434720 517596
rect 342220 517556 342226 517568
rect 434714 517556 434720 517568
rect 434772 517556 434778 517608
rect 436646 517556 436652 517608
rect 436704 517596 436710 517608
rect 436922 517596 436928 517608
rect 436704 517568 436928 517596
rect 436704 517556 436710 517568
rect 436922 517556 436928 517568
rect 436980 517596 436986 517608
rect 445386 517596 445392 517608
rect 436980 517568 445392 517596
rect 436980 517556 436986 517568
rect 445386 517556 445392 517568
rect 445444 517556 445450 517608
rect 328454 517528 328460 517540
rect 325804 517500 328460 517528
rect 328454 517488 328460 517500
rect 328512 517488 328518 517540
rect 333238 517488 333244 517540
rect 333296 517528 333302 517540
rect 336734 517528 336740 517540
rect 333296 517500 336740 517528
rect 333296 517488 333302 517500
rect 336734 517488 336740 517500
rect 336792 517488 336798 517540
rect 337378 517488 337384 517540
rect 337436 517528 337442 517540
rect 339494 517528 339500 517540
rect 337436 517500 339500 517528
rect 337436 517488 337442 517500
rect 339494 517488 339500 517500
rect 339552 517488 339558 517540
rect 379606 514020 379612 514072
rect 379664 514060 379670 514072
rect 379790 514060 379796 514072
rect 379664 514032 379796 514060
rect 379664 514020 379670 514032
rect 379790 514020 379796 514032
rect 379848 514020 379854 514072
rect 542538 511980 542544 512032
rect 542596 512020 542602 512032
rect 542814 512020 542820 512032
rect 542596 511992 542820 512020
rect 542596 511980 542602 511992
rect 542814 511980 542820 511992
rect 542872 511980 542878 512032
rect 433794 511912 433800 511964
rect 433852 511952 433858 511964
rect 433886 511952 433892 511964
rect 433852 511924 433892 511952
rect 433852 511912 433858 511924
rect 433886 511912 433892 511924
rect 433944 511912 433950 511964
rect 3326 509260 3332 509312
rect 3384 509300 3390 509312
rect 519998 509300 520004 509312
rect 3384 509272 520004 509300
rect 3384 509260 3390 509272
rect 519998 509260 520004 509272
rect 520056 509260 520062 509312
rect 536098 509260 536104 509312
rect 536156 509300 536162 509312
rect 580166 509300 580172 509312
rect 536156 509272 580172 509300
rect 536156 509260 536162 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 433794 502324 433800 502376
rect 433852 502364 433858 502376
rect 434070 502364 434076 502376
rect 433852 502336 434076 502364
rect 433852 502324 433858 502336
rect 434070 502324 434076 502336
rect 434128 502324 434134 502376
rect 542630 502324 542636 502376
rect 542688 502364 542694 502376
rect 542814 502364 542820 502376
rect 542688 502336 542820 502364
rect 542688 502324 542694 502336
rect 542814 502324 542820 502336
rect 542872 502324 542878 502376
rect 379606 499536 379612 499588
rect 379664 499576 379670 499588
rect 379790 499576 379796 499588
rect 379664 499548 379796 499576
rect 379664 499536 379670 499548
rect 379790 499536 379796 499548
rect 379848 499536 379854 499588
rect 554038 498176 554044 498228
rect 554096 498216 554102 498228
rect 580166 498216 580172 498228
rect 554096 498188 580172 498216
rect 554096 498176 554102 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 3418 495456 3424 495508
rect 3476 495496 3482 495508
rect 521286 495496 521292 495508
rect 3476 495468 521292 495496
rect 3476 495456 3482 495468
rect 521286 495456 521292 495468
rect 521344 495456 521350 495508
rect 379606 494708 379612 494760
rect 379664 494748 379670 494760
rect 379790 494748 379796 494760
rect 379664 494720 379796 494748
rect 379664 494708 379670 494720
rect 379790 494708 379796 494720
rect 379848 494708 379854 494760
rect 433610 492600 433616 492652
rect 433668 492640 433674 492652
rect 433886 492640 433892 492652
rect 433668 492612 433892 492640
rect 433668 492600 433674 492612
rect 433886 492600 433892 492612
rect 433944 492600 433950 492652
rect 542538 492600 542544 492652
rect 542596 492640 542602 492652
rect 542630 492640 542636 492652
rect 542596 492612 542636 492640
rect 542596 492600 542602 492612
rect 542630 492600 542636 492612
rect 542688 492600 542694 492652
rect 523862 485800 523868 485852
rect 523920 485840 523926 485852
rect 580166 485840 580172 485852
rect 523920 485812 580172 485840
rect 523920 485800 523926 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 542538 485732 542544 485784
rect 542596 485772 542602 485784
rect 542630 485772 542636 485784
rect 542596 485744 542636 485772
rect 542596 485732 542602 485744
rect 542630 485732 542636 485744
rect 542688 485732 542694 485784
rect 297818 482944 297824 482996
rect 297876 482984 297882 482996
rect 299566 482984 299572 482996
rect 297876 482956 299572 482984
rect 297876 482944 297882 482956
rect 299566 482944 299572 482956
rect 299624 482944 299630 482996
rect 307662 482944 307668 482996
rect 307720 482984 307726 482996
rect 307720 482956 383240 482984
rect 307720 482944 307726 482956
rect 297450 482876 297456 482928
rect 297508 482916 297514 482928
rect 383212 482916 383240 482956
rect 428826 482944 428832 482996
rect 428884 482984 428890 482996
rect 439498 482984 439504 482996
rect 428884 482956 439504 482984
rect 428884 482944 428890 482956
rect 439498 482944 439504 482956
rect 439556 482944 439562 482996
rect 455322 482944 455328 482996
rect 455380 482984 455386 482996
rect 492030 482984 492036 482996
rect 455380 482956 492036 482984
rect 455380 482944 455386 482956
rect 492030 482944 492036 482956
rect 492088 482944 492094 482996
rect 390738 482916 390744 482928
rect 297508 482888 383056 482916
rect 383212 482888 390744 482916
rect 297508 482876 297514 482888
rect 283466 482808 283472 482860
rect 283524 482848 283530 482860
rect 379698 482848 379704 482860
rect 283524 482820 379704 482848
rect 283524 482808 283530 482820
rect 379698 482808 379704 482820
rect 379756 482808 379762 482860
rect 383028 482848 383056 482888
rect 390738 482876 390744 482888
rect 390796 482876 390802 482928
rect 426158 482876 426164 482928
rect 426216 482916 426222 482928
rect 438118 482916 438124 482928
rect 426216 482888 438124 482916
rect 426216 482876 426222 482888
rect 438118 482876 438124 482888
rect 438176 482876 438182 482928
rect 453850 482876 453856 482928
rect 453908 482916 453914 482928
rect 489914 482916 489920 482928
rect 453908 482888 489920 482916
rect 453908 482876 453914 482888
rect 489914 482876 489920 482888
rect 489972 482876 489978 482928
rect 387610 482848 387616 482860
rect 383028 482820 387616 482848
rect 387610 482808 387616 482820
rect 387668 482808 387674 482860
rect 433242 482808 433248 482860
rect 433300 482848 433306 482860
rect 450262 482848 450268 482860
rect 433300 482820 450268 482848
rect 433300 482808 433306 482820
rect 450262 482808 450268 482820
rect 450320 482808 450326 482860
rect 458082 482808 458088 482860
rect 458140 482848 458146 482860
rect 496446 482848 496452 482860
rect 458140 482820 496452 482848
rect 458140 482808 458146 482820
rect 496446 482808 496452 482820
rect 496504 482808 496510 482860
rect 297542 482740 297548 482792
rect 297600 482780 297606 482792
rect 387334 482780 387340 482792
rect 297600 482752 387340 482780
rect 297600 482740 297606 482752
rect 387334 482740 387340 482752
rect 387392 482740 387398 482792
rect 434622 482740 434628 482792
rect 434680 482780 434686 482792
rect 452654 482780 452660 482792
rect 434680 482752 452660 482780
rect 434680 482740 434686 482752
rect 452654 482740 452660 482752
rect 452712 482740 452718 482792
rect 456702 482740 456708 482792
rect 456760 482780 456766 482792
rect 494238 482780 494244 482792
rect 456760 482752 494244 482780
rect 456760 482740 456766 482752
rect 494238 482740 494244 482752
rect 494296 482740 494302 482792
rect 281350 482672 281356 482724
rect 281408 482712 281414 482724
rect 379790 482712 379796 482724
rect 281408 482684 379796 482712
rect 281408 482672 281414 482684
rect 379790 482672 379796 482684
rect 379848 482672 379854 482724
rect 382642 482672 382648 482724
rect 382700 482712 382706 482724
rect 383562 482712 383568 482724
rect 382700 482684 383568 482712
rect 382700 482672 382706 482684
rect 383562 482672 383568 482684
rect 383620 482672 383626 482724
rect 386966 482672 386972 482724
rect 387024 482712 387030 482724
rect 387702 482712 387708 482724
rect 387024 482684 387708 482712
rect 387024 482672 387030 482684
rect 387702 482672 387708 482684
rect 387760 482672 387766 482724
rect 436002 482672 436008 482724
rect 436060 482712 436066 482724
rect 454586 482712 454592 482724
rect 436060 482684 454592 482712
rect 436060 482672 436066 482684
rect 454586 482672 454592 482684
rect 454644 482672 454650 482724
rect 459462 482672 459468 482724
rect 459520 482712 459526 482724
rect 498654 482712 498660 482724
rect 459520 482684 498660 482712
rect 459520 482672 459526 482684
rect 498654 482672 498660 482684
rect 498712 482672 498718 482724
rect 297634 482604 297640 482656
rect 297692 482644 297698 482656
rect 397454 482644 397460 482656
rect 297692 482616 397460 482644
rect 297692 482604 297698 482616
rect 397454 482604 397460 482616
rect 397512 482604 397518 482656
rect 437382 482604 437388 482656
rect 437440 482644 437446 482656
rect 456886 482644 456892 482656
rect 437440 482616 456892 482644
rect 437440 482604 437446 482616
rect 456886 482604 456892 482616
rect 456944 482604 456950 482656
rect 460842 482604 460848 482656
rect 460900 482644 460906 482656
rect 500954 482644 500960 482656
rect 460900 482616 500960 482644
rect 460900 482604 460906 482616
rect 500954 482604 500960 482616
rect 501012 482604 501018 482656
rect 287882 482536 287888 482588
rect 287940 482576 287946 482588
rect 288342 482576 288348 482588
rect 287940 482548 288348 482576
rect 287940 482536 287946 482548
rect 288342 482536 288348 482548
rect 288400 482536 288406 482588
rect 294506 482536 294512 482588
rect 294564 482576 294570 482588
rect 295242 482576 295248 482588
rect 294564 482548 295248 482576
rect 294564 482536 294570 482548
rect 295242 482536 295248 482548
rect 295300 482536 295306 482588
rect 298922 482536 298928 482588
rect 298980 482576 298986 482588
rect 299382 482576 299388 482588
rect 298980 482548 299388 482576
rect 298980 482536 298986 482548
rect 299382 482536 299388 482548
rect 299440 482536 299446 482588
rect 399570 482576 399576 482588
rect 299492 482548 399576 482576
rect 297726 482468 297732 482520
rect 297784 482508 297790 482520
rect 299492 482508 299520 482548
rect 399570 482536 399576 482548
rect 399628 482536 399634 482588
rect 424410 482536 424416 482588
rect 424468 482576 424474 482588
rect 436738 482576 436744 482588
rect 424468 482548 436744 482576
rect 424468 482536 424474 482548
rect 436738 482536 436744 482548
rect 436796 482536 436802 482588
rect 438670 482536 438676 482588
rect 438728 482576 438734 482588
rect 459002 482576 459008 482588
rect 438728 482548 459008 482576
rect 438728 482536 438734 482548
rect 459002 482536 459008 482548
rect 459060 482536 459066 482588
rect 460750 482536 460756 482588
rect 460808 482576 460814 482588
rect 503070 482576 503076 482588
rect 460808 482548 503076 482576
rect 460808 482536 460814 482548
rect 503070 482536 503076 482548
rect 503128 482536 503134 482588
rect 297784 482480 299520 482508
rect 297784 482468 297790 482480
rect 299566 482468 299572 482520
rect 299624 482508 299630 482520
rect 401778 482508 401784 482520
rect 299624 482480 401784 482508
rect 299624 482468 299630 482480
rect 401778 482468 401784 482480
rect 401836 482468 401842 482520
rect 419994 482468 420000 482520
rect 420052 482508 420058 482520
rect 435358 482508 435364 482520
rect 420052 482480 435364 482508
rect 420052 482468 420058 482480
rect 435358 482468 435364 482480
rect 435416 482468 435422 482520
rect 438762 482468 438768 482520
rect 438820 482508 438826 482520
rect 461210 482508 461216 482520
rect 438820 482480 461216 482508
rect 438820 482468 438826 482480
rect 461210 482468 461216 482480
rect 461268 482468 461274 482520
rect 462222 482468 462228 482520
rect 462280 482508 462286 482520
rect 505278 482508 505284 482520
rect 462280 482480 505284 482508
rect 462280 482468 462286 482480
rect 505278 482468 505284 482480
rect 505336 482468 505342 482520
rect 297910 482400 297916 482452
rect 297968 482440 297974 482452
rect 403986 482440 403992 482452
rect 297968 482412 403992 482440
rect 297968 482400 297974 482412
rect 403986 482400 403992 482412
rect 404044 482400 404050 482452
rect 422202 482400 422208 482452
rect 422260 482440 422266 482452
rect 436922 482440 436928 482452
rect 422260 482412 436928 482440
rect 422260 482400 422266 482412
rect 436922 482400 436928 482412
rect 436980 482400 436986 482452
rect 440142 482400 440148 482452
rect 440200 482440 440206 482452
rect 463694 482440 463700 482452
rect 440200 482412 463700 482440
rect 440200 482400 440206 482412
rect 463694 482400 463700 482412
rect 463752 482400 463758 482452
rect 464982 482400 464988 482452
rect 465040 482440 465046 482452
rect 509694 482440 509700 482452
rect 465040 482412 509700 482440
rect 465040 482400 465046 482412
rect 509694 482400 509700 482412
rect 509752 482400 509758 482452
rect 298002 482332 298008 482384
rect 298060 482372 298066 482384
rect 406194 482372 406200 482384
rect 298060 482344 406200 482372
rect 298060 482332 298066 482344
rect 406194 482332 406200 482344
rect 406252 482332 406258 482384
rect 417786 482332 417792 482384
rect 417844 482372 417850 482384
rect 433794 482372 433800 482384
rect 417844 482344 433800 482372
rect 417844 482332 417850 482344
rect 433794 482332 433800 482344
rect 433852 482332 433858 482384
rect 441522 482332 441528 482384
rect 441580 482372 441586 482384
rect 465626 482372 465632 482384
rect 441580 482344 465632 482372
rect 441580 482332 441586 482344
rect 465626 482332 465632 482344
rect 465684 482332 465690 482384
rect 466362 482332 466368 482384
rect 466420 482372 466426 482384
rect 511994 482372 512000 482384
rect 466420 482344 512000 482372
rect 466420 482332 466426 482344
rect 511994 482332 512000 482344
rect 512052 482332 512058 482384
rect 297358 482264 297364 482316
rect 297416 482304 297422 482316
rect 412818 482304 412824 482316
rect 297416 482276 412824 482304
rect 297416 482264 297422 482276
rect 412818 482264 412824 482276
rect 412876 482264 412882 482316
rect 415210 482264 415216 482316
rect 415268 482304 415274 482316
rect 432598 482304 432604 482316
rect 415268 482276 432604 482304
rect 415268 482264 415274 482276
rect 432598 482264 432604 482276
rect 432656 482264 432662 482316
rect 442902 482264 442908 482316
rect 442960 482304 442966 482316
rect 467834 482304 467840 482316
rect 442960 482276 467840 482304
rect 442960 482264 442966 482276
rect 467834 482264 467840 482276
rect 467892 482264 467898 482316
rect 469122 482264 469128 482316
rect 469180 482304 469186 482316
rect 516318 482304 516324 482316
rect 469180 482276 516324 482304
rect 469180 482264 469186 482276
rect 516318 482264 516324 482276
rect 516376 482264 516382 482316
rect 305546 482196 305552 482248
rect 305604 482236 305610 482248
rect 306282 482236 306288 482248
rect 305604 482208 306288 482236
rect 305604 482196 305610 482208
rect 306282 482196 306288 482208
rect 306340 482196 306346 482248
rect 309962 482196 309968 482248
rect 310020 482236 310026 482248
rect 310422 482236 310428 482248
rect 310020 482208 310428 482236
rect 310020 482196 310026 482208
rect 310422 482196 310428 482208
rect 310480 482196 310486 482248
rect 311710 482196 311716 482248
rect 311768 482236 311774 482248
rect 371234 482236 371240 482248
rect 311768 482208 371240 482236
rect 311768 482196 311774 482208
rect 371234 482196 371240 482208
rect 371292 482196 371298 482248
rect 376018 482196 376024 482248
rect 376076 482236 376082 482248
rect 410518 482236 410524 482248
rect 376076 482208 410524 482236
rect 376076 482196 376082 482208
rect 410518 482196 410524 482208
rect 410576 482196 410582 482248
rect 431034 482196 431040 482248
rect 431092 482236 431098 482248
rect 440878 482236 440884 482248
rect 431092 482208 440884 482236
rect 431092 482196 431098 482208
rect 440878 482196 440884 482208
rect 440936 482196 440942 482248
rect 453942 482196 453948 482248
rect 454000 482236 454006 482248
rect 487614 482236 487620 482248
rect 454000 482208 487620 482236
rect 454000 482196 454006 482208
rect 487614 482196 487620 482208
rect 487672 482196 487678 482248
rect 310238 482128 310244 482180
rect 310296 482168 310302 482180
rect 368750 482168 368756 482180
rect 310296 482140 368756 482168
rect 310296 482128 310302 482140
rect 368750 482128 368756 482140
rect 368808 482128 368814 482180
rect 387610 482128 387616 482180
rect 387668 482168 387674 482180
rect 392946 482168 392952 482180
rect 387668 482140 392952 482168
rect 387668 482128 387674 482140
rect 392946 482128 392952 482140
rect 393004 482128 393010 482180
rect 452562 482128 452568 482180
rect 452620 482168 452626 482180
rect 485774 482168 485780 482180
rect 452620 482140 485780 482168
rect 452620 482128 452626 482140
rect 485774 482128 485780 482140
rect 485832 482128 485838 482180
rect 310330 482060 310336 482112
rect 310388 482100 310394 482112
rect 366542 482100 366548 482112
rect 310388 482072 366548 482100
rect 310388 482060 310394 482072
rect 366542 482060 366548 482072
rect 366600 482060 366606 482112
rect 451182 482060 451188 482112
rect 451240 482100 451246 482112
rect 483290 482100 483296 482112
rect 451240 482072 483296 482100
rect 451240 482060 451246 482072
rect 483290 482060 483296 482072
rect 483348 482060 483354 482112
rect 309042 481992 309048 482044
rect 309100 482032 309106 482044
rect 364334 482032 364340 482044
rect 309100 482004 364340 482032
rect 309100 481992 309106 482004
rect 364334 481992 364340 482004
rect 364392 481992 364398 482044
rect 448422 481992 448428 482044
rect 448480 482032 448486 482044
rect 478874 482032 478880 482044
rect 448480 482004 478880 482032
rect 448480 481992 448486 482004
rect 478874 481992 478880 482004
rect 478932 481992 478938 482044
rect 316494 481924 316500 481976
rect 316552 481964 316558 481976
rect 317322 481964 317328 481976
rect 316552 481936 317328 481964
rect 316552 481924 316558 481936
rect 317322 481924 317328 481936
rect 317380 481924 317386 481976
rect 320910 481924 320916 481976
rect 320968 481964 320974 481976
rect 321462 481964 321468 481976
rect 320968 481936 321468 481964
rect 320968 481924 320974 481936
rect 321462 481924 321468 481936
rect 321520 481924 321526 481976
rect 327534 481924 327540 481976
rect 327592 481964 327598 481976
rect 328362 481964 328368 481976
rect 327592 481936 328368 481964
rect 327592 481924 327598 481936
rect 328362 481924 328368 481936
rect 328420 481924 328426 481976
rect 329742 481924 329748 481976
rect 329800 481964 329806 481976
rect 330478 481964 330484 481976
rect 329800 481936 330484 481964
rect 329800 481924 329806 481936
rect 330478 481924 330484 481936
rect 330536 481924 330542 481976
rect 331950 481924 331956 481976
rect 332008 481964 332014 481976
rect 333238 481964 333244 481976
rect 332008 481936 333244 481964
rect 332008 481924 332014 481936
rect 333238 481924 333244 481936
rect 333296 481924 333302 481976
rect 336366 481924 336372 481976
rect 336424 481964 336430 481976
rect 337378 481964 337384 481976
rect 336424 481936 337384 481964
rect 336424 481924 336430 481936
rect 337378 481924 337384 481936
rect 337436 481924 337442 481976
rect 338574 481924 338580 481976
rect 338632 481964 338638 481976
rect 339402 481964 339408 481976
rect 338632 481936 339408 481964
rect 338632 481924 338638 481936
rect 339402 481924 339408 481936
rect 339460 481924 339466 481976
rect 346302 481924 346308 481976
rect 346360 481964 346366 481976
rect 346762 481964 346768 481976
rect 346360 481936 346768 481964
rect 346360 481924 346366 481936
rect 346762 481924 346768 481936
rect 346820 481924 346826 481976
rect 348418 481924 348424 481976
rect 348476 481964 348482 481976
rect 349154 481964 349160 481976
rect 348476 481936 349160 481964
rect 348476 481924 348482 481936
rect 349154 481924 349160 481936
rect 349212 481924 349218 481976
rect 349246 481924 349252 481976
rect 349304 481964 349310 481976
rect 351086 481964 351092 481976
rect 349304 481936 351092 481964
rect 349304 481924 349310 481936
rect 351086 481924 351092 481936
rect 351144 481924 351150 481976
rect 358262 481924 358268 481976
rect 358320 481964 358326 481976
rect 358722 481964 358728 481976
rect 358320 481936 358728 481964
rect 358320 481924 358326 481936
rect 358722 481924 358728 481936
rect 358780 481924 358786 481976
rect 449802 481924 449808 481976
rect 449860 481964 449866 481976
rect 481082 481964 481088 481976
rect 449860 481936 481088 481964
rect 449860 481924 449866 481936
rect 481082 481924 481088 481936
rect 481140 481924 481146 481976
rect 325326 481856 325332 481908
rect 325384 481896 325390 481908
rect 327718 481896 327724 481908
rect 325384 481868 327724 481896
rect 325384 481856 325390 481868
rect 327718 481856 327724 481868
rect 327776 481856 327782 481908
rect 360562 481856 360568 481908
rect 360620 481896 360626 481908
rect 361482 481896 361488 481908
rect 360620 481868 361488 481896
rect 360620 481856 360626 481868
rect 361482 481856 361488 481868
rect 361540 481856 361546 481908
rect 445570 481856 445576 481908
rect 445628 481896 445634 481908
rect 474734 481896 474740 481908
rect 445628 481868 474740 481896
rect 445628 481856 445634 481868
rect 474734 481856 474740 481868
rect 474792 481856 474798 481908
rect 318702 481788 318708 481840
rect 318760 481828 318766 481840
rect 326338 481828 326344 481840
rect 318760 481800 326344 481828
rect 318760 481788 318766 481800
rect 326338 481788 326344 481800
rect 326396 481788 326402 481840
rect 348970 481788 348976 481840
rect 349028 481828 349034 481840
rect 353294 481828 353300 481840
rect 349028 481800 353300 481828
rect 349028 481788 349034 481800
rect 353294 481788 353300 481800
rect 353352 481788 353358 481840
rect 447042 481788 447048 481840
rect 447100 481828 447106 481840
rect 476666 481828 476672 481840
rect 447100 481800 476672 481828
rect 447100 481788 447106 481800
rect 476666 481788 476672 481800
rect 476724 481788 476730 481840
rect 445662 481720 445668 481772
rect 445720 481760 445726 481772
rect 472250 481760 472256 481772
rect 445720 481732 472256 481760
rect 445720 481720 445726 481732
rect 472250 481720 472256 481732
rect 472308 481720 472314 481772
rect 444282 481652 444288 481704
rect 444340 481692 444346 481704
rect 470042 481692 470048 481704
rect 444340 481664 470048 481692
rect 444340 481652 444346 481664
rect 470042 481652 470048 481664
rect 470100 481652 470106 481704
rect 2958 480224 2964 480276
rect 3016 480264 3022 480276
rect 520182 480264 520188 480276
rect 3016 480236 520188 480264
rect 3016 480224 3022 480236
rect 520182 480224 520188 480236
rect 520240 480224 520246 480276
rect 387334 480088 387340 480140
rect 387392 480128 387398 480140
rect 395476 480128 395482 480140
rect 387392 480100 395482 480128
rect 387392 480088 387398 480100
rect 395476 480088 395482 480100
rect 395534 480088 395540 480140
rect 367186 479816 367192 479868
rect 367244 479856 367250 479868
rect 369946 479856 369952 479868
rect 367244 479828 369952 479856
rect 367244 479816 367250 479828
rect 369946 479816 369952 479828
rect 370004 479816 370010 479868
rect 398742 479816 398748 479868
rect 398800 479856 398806 479868
rect 520090 479856 520096 479868
rect 398800 479828 520096 479856
rect 398800 479816 398806 479828
rect 520090 479816 520096 479828
rect 520148 479816 520154 479868
rect 300578 479748 300584 479800
rect 300636 479788 300642 479800
rect 520918 479788 520924 479800
rect 300636 479760 520924 479788
rect 300636 479748 300642 479760
rect 520918 479748 520924 479760
rect 520976 479748 520982 479800
rect 235902 479680 235908 479732
rect 235960 479720 235966 479732
rect 521010 479720 521016 479732
rect 235960 479692 521016 479720
rect 235960 479680 235966 479692
rect 521010 479680 521016 479692
rect 521068 479680 521074 479732
rect 171042 479612 171048 479664
rect 171100 479652 171106 479664
rect 521102 479652 521108 479664
rect 171100 479624 521108 479652
rect 171100 479612 171106 479624
rect 521102 479612 521108 479624
rect 521160 479612 521166 479664
rect 106182 479544 106188 479596
rect 106240 479584 106246 479596
rect 521194 479584 521200 479596
rect 106240 479556 521200 479584
rect 106240 479544 106246 479556
rect 521194 479544 521200 479556
rect 521252 479544 521258 479596
rect 3602 479476 3608 479528
rect 3660 479516 3666 479528
rect 521378 479516 521384 479528
rect 3660 479488 521384 479516
rect 3660 479476 3666 479488
rect 521378 479476 521384 479488
rect 521436 479476 521442 479528
rect 50982 479408 50988 479460
rect 51040 479448 51046 479460
rect 57790 479448 57796 479460
rect 51040 479420 57796 479448
rect 51040 479408 51046 479420
rect 57790 479408 57796 479420
rect 57848 479408 57854 479460
rect 128262 479408 128268 479460
rect 128320 479448 128326 479460
rect 135162 479448 135168 479460
rect 128320 479420 135168 479448
rect 128320 479408 128326 479420
rect 135162 479408 135168 479420
rect 135220 479408 135226 479460
rect 278866 479408 278872 479460
rect 278924 479448 278930 479460
rect 283558 479448 283564 479460
rect 278924 479420 283564 479448
rect 278924 479408 278930 479420
rect 283558 479408 283564 479420
rect 283616 479408 283622 479460
rect 466362 479408 466368 479460
rect 466420 479448 466426 479460
rect 473262 479448 473268 479460
rect 466420 479420 473268 479448
rect 466420 479408 466426 479420
rect 473262 479408 473268 479420
rect 473320 479408 473326 479460
rect 147582 479340 147588 479392
rect 147640 479380 147646 479392
rect 154482 479380 154488 479392
rect 147640 479352 154488 479380
rect 147640 479340 147646 479352
rect 154482 479340 154488 479352
rect 154540 479340 154546 479392
rect 166902 479340 166908 479392
rect 166960 479380 166966 479392
rect 173802 479380 173808 479392
rect 166960 479352 173808 479380
rect 166960 479340 166966 479352
rect 173802 479340 173808 479352
rect 173860 479340 173866 479392
rect 186222 479340 186228 479392
rect 186280 479380 186286 479392
rect 193122 479380 193128 479392
rect 186280 479352 193128 479380
rect 186280 479340 186286 479352
rect 193122 479340 193128 479352
rect 193180 479340 193186 479392
rect 205542 479340 205548 479392
rect 205600 479380 205606 479392
rect 212442 479380 212448 479392
rect 205600 479352 212448 479380
rect 205600 479340 205606 479352
rect 212442 479340 212448 479352
rect 212500 479340 212506 479392
rect 224862 479340 224868 479392
rect 224920 479380 224926 479392
rect 231762 479380 231768 479392
rect 224920 479352 231768 479380
rect 224920 479340 224926 479352
rect 231762 479340 231768 479352
rect 231820 479340 231826 479392
rect 244182 479340 244188 479392
rect 244240 479380 244246 479392
rect 251082 479380 251088 479392
rect 244240 479352 251088 479380
rect 244240 479340 244246 479352
rect 251082 479340 251088 479352
rect 251140 479340 251146 479392
rect 485682 479340 485688 479392
rect 485740 479380 485746 479392
rect 492582 479380 492588 479392
rect 485740 479352 492588 479380
rect 485740 479340 485746 479352
rect 492582 479340 492588 479352
rect 492640 479340 492646 479392
rect 57974 479272 57980 479324
rect 58032 479312 58038 479324
rect 61838 479312 61844 479324
rect 58032 479284 61844 479312
rect 58032 479272 58038 479284
rect 61838 479272 61844 479284
rect 61896 479272 61902 479324
rect 309134 479272 309140 479324
rect 309192 479312 309198 479324
rect 316770 479312 316776 479324
rect 309192 479284 316776 479312
rect 309192 479272 309198 479284
rect 316770 479272 316776 479284
rect 316828 479272 316834 479324
rect 279694 479136 279700 479188
rect 279752 479176 279758 479188
rect 519906 479176 519912 479188
rect 279752 479148 519912 479176
rect 279752 479136 279758 479148
rect 519906 479136 519912 479148
rect 519964 479136 519970 479188
rect 279602 479068 279608 479120
rect 279660 479108 279666 479120
rect 521562 479108 521568 479120
rect 279660 479080 521568 479108
rect 279660 479068 279666 479080
rect 521562 479068 521568 479080
rect 521620 479068 521626 479120
rect 279970 479000 279976 479052
rect 280028 479040 280034 479052
rect 523126 479040 523132 479052
rect 280028 479012 523132 479040
rect 280028 479000 280034 479012
rect 523126 479000 523132 479012
rect 523184 479000 523190 479052
rect 135162 478932 135168 478984
rect 135220 478972 135226 478984
rect 277394 478972 277400 478984
rect 135220 478944 277400 478972
rect 135220 478932 135226 478944
rect 277394 478932 277400 478944
rect 277452 478932 277458 478984
rect 279878 478932 279884 478984
rect 279936 478972 279942 478984
rect 523034 478972 523040 478984
rect 279936 478944 523040 478972
rect 279936 478932 279942 478944
rect 523034 478932 523040 478944
rect 523092 478932 523098 478984
rect 3418 478864 3424 478916
rect 3476 478904 3482 478916
rect 519814 478904 519820 478916
rect 3476 478876 519820 478904
rect 3476 478864 3482 478876
rect 519814 478864 519820 478876
rect 519872 478864 519878 478916
rect 520090 478728 520096 478780
rect 520148 478728 520154 478780
rect 519906 478660 519912 478712
rect 519964 478700 519970 478712
rect 520108 478700 520136 478728
rect 519964 478672 520136 478700
rect 519964 478660 519970 478672
rect 279142 478524 279148 478576
rect 279200 478564 279206 478576
rect 520182 478564 520188 478576
rect 279200 478536 520188 478564
rect 279200 478524 279206 478536
rect 520182 478524 520188 478536
rect 520240 478524 520246 478576
rect 280062 478456 280068 478508
rect 280120 478496 280126 478508
rect 521470 478496 521476 478508
rect 280120 478468 521476 478496
rect 280120 478456 280126 478468
rect 521470 478456 521476 478468
rect 521528 478456 521534 478508
rect 279786 478388 279792 478440
rect 279844 478428 279850 478440
rect 522666 478428 522672 478440
rect 279844 478400 522672 478428
rect 279844 478388 279850 478400
rect 522666 478388 522672 478400
rect 522724 478388 522730 478440
rect 279510 478320 279516 478372
rect 279568 478360 279574 478372
rect 522850 478360 522856 478372
rect 279568 478332 522856 478360
rect 279568 478320 279574 478332
rect 522850 478320 522856 478332
rect 522908 478320 522914 478372
rect 3786 478252 3792 478304
rect 3844 478292 3850 478304
rect 522482 478292 522488 478304
rect 3844 478264 522488 478292
rect 3844 478252 3850 478264
rect 522482 478252 522488 478264
rect 522540 478252 522546 478304
rect 3510 478184 3516 478236
rect 3568 478224 3574 478236
rect 522298 478224 522304 478236
rect 3568 478196 522304 478224
rect 3568 478184 3574 478196
rect 522298 478184 522304 478196
rect 522356 478184 522362 478236
rect 3694 478116 3700 478168
rect 3752 478156 3758 478168
rect 522574 478156 522580 478168
rect 3752 478128 522580 478156
rect 3752 478116 3758 478128
rect 522574 478116 522580 478128
rect 522632 478116 522638 478168
rect 279234 478048 279240 478100
rect 279292 478088 279298 478100
rect 522758 478088 522764 478100
rect 279292 478060 522764 478088
rect 279292 478048 279298 478060
rect 522758 478048 522764 478060
rect 522816 478048 522822 478100
rect 279418 477980 279424 478032
rect 279476 478020 279482 478032
rect 522390 478020 522396 478032
rect 279476 477992 522396 478020
rect 279476 477980 279482 477992
rect 522390 477980 522396 477992
rect 522448 477980 522454 478032
rect 279326 477912 279332 477964
rect 279384 477952 279390 477964
rect 524414 477952 524420 477964
rect 279384 477924 524420 477952
rect 279384 477912 279390 477924
rect 524414 477912 524420 477924
rect 524472 477912 524478 477964
rect 133782 476076 133788 476128
rect 133840 476116 133846 476128
rect 277394 476116 277400 476128
rect 133840 476088 277400 476116
rect 133840 476076 133846 476088
rect 277394 476076 277400 476088
rect 277452 476076 277458 476128
rect 542446 476076 542452 476128
rect 542504 476116 542510 476128
rect 542630 476116 542636 476128
rect 542504 476088 542636 476116
rect 542504 476076 542510 476088
rect 542630 476076 542636 476088
rect 542688 476076 542694 476128
rect 132402 473356 132408 473408
rect 132460 473396 132466 473408
rect 278682 473396 278688 473408
rect 132460 473368 278688 473396
rect 132460 473356 132466 473368
rect 278682 473356 278688 473368
rect 278740 473356 278746 473408
rect 542538 473288 542544 473340
rect 542596 473328 542602 473340
rect 542630 473328 542636 473340
rect 542596 473300 542636 473328
rect 542596 473288 542602 473300
rect 542630 473288 542636 473300
rect 542688 473288 542694 473340
rect 131022 471996 131028 472048
rect 131080 472036 131086 472048
rect 278682 472036 278688 472048
rect 131080 472008 278688 472036
rect 131080 471996 131086 472008
rect 278682 471996 278688 472008
rect 278740 471996 278746 472048
rect 129642 469208 129648 469260
rect 129700 469248 129706 469260
rect 277854 469248 277860 469260
rect 129700 469220 277860 469248
rect 129700 469208 129706 469220
rect 277854 469208 277860 469220
rect 277912 469208 277918 469260
rect 128262 467848 128268 467900
rect 128320 467888 128326 467900
rect 278682 467888 278688 467900
rect 128320 467860 278688 467888
rect 128320 467848 128326 467860
rect 278682 467848 278688 467860
rect 278740 467848 278746 467900
rect 542630 466460 542636 466472
rect 542556 466432 542636 466460
rect 542556 466404 542584 466432
rect 542630 466420 542636 466432
rect 542688 466420 542694 466472
rect 542538 466352 542544 466404
rect 542596 466352 542602 466404
rect 126882 465060 126888 465112
rect 126940 465100 126946 465112
rect 278682 465100 278688 465112
rect 126940 465072 278688 465100
rect 126940 465060 126946 465072
rect 278682 465060 278688 465072
rect 278740 465060 278746 465112
rect 125502 463700 125508 463752
rect 125560 463740 125566 463752
rect 278682 463740 278688 463752
rect 125560 463712 278688 463740
rect 125560 463700 125566 463712
rect 278682 463700 278688 463712
rect 278740 463700 278746 463752
rect 549898 462340 549904 462392
rect 549956 462380 549962 462392
rect 580166 462380 580172 462392
rect 549956 462352 580172 462380
rect 549956 462340 549962 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 125410 460912 125416 460964
rect 125468 460952 125474 460964
rect 278682 460952 278688 460964
rect 125468 460924 278688 460952
rect 125468 460912 125474 460924
rect 278682 460912 278688 460924
rect 278740 460912 278746 460964
rect 124122 459552 124128 459604
rect 124180 459592 124186 459604
rect 278682 459592 278688 459604
rect 124180 459564 278688 459592
rect 124180 459552 124186 459564
rect 278682 459552 278688 459564
rect 278740 459552 278746 459604
rect 122742 456764 122748 456816
rect 122800 456804 122806 456816
rect 278682 456804 278688 456816
rect 122800 456776 278688 456804
rect 122800 456764 122806 456776
rect 278682 456764 278688 456776
rect 278740 456764 278746 456816
rect 121362 455404 121368 455456
rect 121420 455444 121426 455456
rect 278682 455444 278688 455456
rect 121420 455416 278688 455444
rect 121420 455404 121426 455416
rect 278682 455404 278688 455416
rect 278740 455404 278746 455456
rect 119982 452616 119988 452668
rect 120040 452656 120046 452668
rect 278682 452656 278688 452668
rect 120040 452628 278688 452656
rect 120040 452616 120046 452628
rect 278682 452616 278688 452628
rect 278740 452616 278746 452668
rect 3510 452548 3516 452600
rect 3568 452588 3574 452600
rect 279142 452588 279148 452600
rect 3568 452560 279148 452588
rect 3568 452548 3574 452560
rect 279142 452548 279148 452560
rect 279200 452548 279206 452600
rect 118602 451256 118608 451308
rect 118660 451296 118666 451308
rect 278682 451296 278688 451308
rect 118660 451268 278688 451296
rect 118660 451256 118666 451268
rect 278682 451256 278688 451268
rect 278740 451256 278746 451308
rect 563698 451256 563704 451308
rect 563756 451296 563762 451308
rect 580166 451296 580172 451308
rect 563756 451268 580172 451296
rect 563756 451256 563762 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 117222 448536 117228 448588
rect 117280 448576 117286 448588
rect 278682 448576 278688 448588
rect 117280 448548 278688 448576
rect 117280 448536 117286 448548
rect 278682 448536 278688 448548
rect 278740 448536 278746 448588
rect 542354 447108 542360 447160
rect 542412 447108 542418 447160
rect 542372 447080 542400 447108
rect 542446 447080 542452 447092
rect 542372 447052 542452 447080
rect 542446 447040 542452 447052
rect 542504 447040 542510 447092
rect 117130 445748 117136 445800
rect 117188 445788 117194 445800
rect 278682 445788 278688 445800
rect 117188 445760 278688 445788
rect 117188 445748 117194 445760
rect 278682 445748 278688 445760
rect 278740 445748 278746 445800
rect 115842 444388 115848 444440
rect 115900 444428 115906 444440
rect 278682 444428 278688 444440
rect 115900 444400 278688 444428
rect 115900 444388 115906 444400
rect 278682 444388 278688 444400
rect 278740 444388 278746 444440
rect 542170 444320 542176 444372
rect 542228 444360 542234 444372
rect 542446 444360 542452 444372
rect 542228 444332 542452 444360
rect 542228 444320 542234 444332
rect 542446 444320 542452 444332
rect 542504 444320 542510 444372
rect 114462 441600 114468 441652
rect 114520 441640 114526 441652
rect 277854 441640 277860 441652
rect 114520 441612 277860 441640
rect 114520 441600 114526 441612
rect 277854 441600 277860 441612
rect 277912 441600 277918 441652
rect 113082 440240 113088 440292
rect 113140 440280 113146 440292
rect 278682 440280 278688 440292
rect 113140 440252 278688 440280
rect 113140 440240 113146 440252
rect 278682 440240 278688 440252
rect 278740 440240 278746 440292
rect 534718 438880 534724 438932
rect 534776 438920 534782 438932
rect 580166 438920 580172 438932
rect 534776 438892 580172 438920
rect 534776 438880 534782 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3510 438812 3516 438864
rect 3568 438852 3574 438864
rect 279234 438852 279240 438864
rect 3568 438824 279240 438852
rect 3568 438812 3574 438824
rect 279234 438812 279240 438824
rect 279292 438812 279298 438864
rect 522206 437628 522212 437640
rect 519832 437600 522212 437628
rect 519832 437504 519860 437600
rect 522206 437588 522212 437600
rect 522264 437588 522270 437640
rect 111702 437452 111708 437504
rect 111760 437492 111766 437504
rect 278682 437492 278688 437504
rect 111760 437464 278688 437492
rect 111760 437452 111766 437464
rect 278682 437452 278688 437464
rect 278740 437452 278746 437504
rect 519814 437452 519820 437504
rect 519872 437452 519878 437504
rect 522206 437452 522212 437504
rect 522264 437492 522270 437504
rect 522942 437492 522948 437504
rect 522264 437464 522948 437492
rect 522264 437452 522270 437464
rect 522942 437452 522948 437464
rect 523000 437452 523006 437504
rect 110322 436092 110328 436144
rect 110380 436132 110386 436144
rect 278038 436132 278044 436144
rect 110380 436104 278044 436132
rect 110380 436092 110386 436104
rect 278038 436092 278044 436104
rect 278096 436092 278102 436144
rect 108942 433304 108948 433356
rect 109000 433344 109006 433356
rect 278682 433344 278688 433356
rect 109000 433316 278688 433344
rect 109000 433304 109006 433316
rect 278682 433304 278688 433316
rect 278740 433304 278746 433356
rect 107562 431944 107568 431996
rect 107620 431984 107626 431996
rect 278682 431984 278688 431996
rect 107620 431956 278688 431984
rect 107620 431944 107626 431956
rect 278682 431944 278688 431956
rect 278740 431944 278746 431996
rect 107470 429156 107476 429208
rect 107528 429196 107534 429208
rect 277670 429196 277676 429208
rect 107528 429168 277676 429196
rect 107528 429156 107534 429168
rect 277670 429156 277676 429168
rect 277728 429156 277734 429208
rect 106182 427796 106188 427848
rect 106240 427836 106246 427848
rect 278682 427836 278688 427848
rect 106240 427808 278688 427836
rect 106240 427796 106246 427808
rect 278682 427796 278688 427808
rect 278740 427796 278746 427848
rect 542354 427796 542360 427848
rect 542412 427796 542418 427848
rect 542372 427768 542400 427796
rect 542446 427768 542452 427780
rect 542372 427740 542452 427768
rect 542446 427728 542452 427740
rect 542504 427728 542510 427780
rect 104802 425076 104808 425128
rect 104860 425116 104866 425128
rect 278682 425116 278688 425128
rect 104860 425088 278688 425116
rect 104860 425076 104866 425088
rect 278682 425076 278688 425088
rect 278740 425076 278746 425128
rect 3234 425008 3240 425060
rect 3292 425048 3298 425060
rect 279326 425048 279332 425060
rect 3292 425020 279332 425048
rect 3292 425008 3298 425020
rect 279326 425008 279332 425020
rect 279384 425008 279390 425060
rect 542170 425008 542176 425060
rect 542228 425048 542234 425060
rect 542446 425048 542452 425060
rect 542228 425020 542452 425048
rect 542228 425008 542234 425020
rect 542446 425008 542452 425020
rect 542504 425008 542510 425060
rect 103422 423648 103428 423700
rect 103480 423688 103486 423700
rect 278682 423688 278688 423700
rect 103480 423660 278688 423688
rect 103480 423648 103486 423660
rect 278682 423648 278688 423660
rect 278740 423648 278746 423700
rect 102042 420928 102048 420980
rect 102100 420968 102106 420980
rect 278682 420968 278688 420980
rect 102100 420940 278688 420968
rect 102100 420928 102106 420940
rect 278682 420928 278688 420940
rect 278740 420928 278746 420980
rect 522666 420044 522672 420096
rect 522724 420084 522730 420096
rect 524414 420084 524420 420096
rect 522724 420056 524420 420084
rect 522724 420044 522730 420056
rect 524414 420044 524420 420056
rect 524472 420044 524478 420096
rect 100662 418140 100668 418192
rect 100720 418180 100726 418192
rect 278682 418180 278688 418192
rect 100720 418152 278688 418180
rect 100720 418140 100726 418152
rect 278682 418140 278688 418152
rect 278740 418140 278746 418192
rect 99282 416780 99288 416832
rect 99340 416820 99346 416832
rect 278682 416820 278688 416832
rect 99340 416792 278688 416820
rect 99340 416780 99346 416792
rect 278682 416780 278688 416792
rect 278740 416780 278746 416832
rect 547138 415420 547144 415472
rect 547196 415460 547202 415472
rect 580166 415460 580172 415472
rect 547196 415432 580172 415460
rect 547196 415420 547202 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 99190 413992 99196 414044
rect 99248 414032 99254 414044
rect 277854 414032 277860 414044
rect 99248 414004 277860 414032
rect 99248 413992 99254 414004
rect 277854 413992 277860 414004
rect 277912 413992 277918 414044
rect 97902 412632 97908 412684
rect 97960 412672 97966 412684
rect 278682 412672 278688 412684
rect 97960 412644 278688 412672
rect 97960 412632 97966 412644
rect 278682 412632 278688 412644
rect 278740 412632 278746 412684
rect 96522 409844 96528 409896
rect 96580 409884 96586 409896
rect 278682 409884 278688 409896
rect 96580 409856 278688 409884
rect 96580 409844 96586 409856
rect 278682 409844 278688 409856
rect 278740 409844 278746 409896
rect 95142 408484 95148 408536
rect 95200 408524 95206 408536
rect 278682 408524 278688 408536
rect 95200 408496 278688 408524
rect 95200 408484 95206 408496
rect 278682 408484 278688 408496
rect 278740 408484 278746 408536
rect 542354 408484 542360 408536
rect 542412 408484 542418 408536
rect 542372 408388 542400 408484
rect 542446 408388 542452 408400
rect 542372 408360 542452 408388
rect 542446 408348 542452 408360
rect 542504 408348 542510 408400
rect 93762 405696 93768 405748
rect 93820 405736 93826 405748
rect 278682 405736 278688 405748
rect 93820 405708 278688 405736
rect 93820 405696 93826 405708
rect 278682 405696 278688 405708
rect 278740 405696 278746 405748
rect 92382 404336 92388 404388
rect 92440 404376 92446 404388
rect 278682 404376 278688 404388
rect 92440 404348 278688 404376
rect 92440 404336 92446 404348
rect 278682 404336 278688 404348
rect 278740 404336 278746 404388
rect 542078 404268 542084 404320
rect 542136 404308 542142 404320
rect 542446 404308 542452 404320
rect 542136 404280 542452 404308
rect 542136 404268 542142 404280
rect 542446 404268 542452 404280
rect 542504 404268 542510 404320
rect 91002 401616 91008 401668
rect 91060 401656 91066 401668
rect 278406 401656 278412 401668
rect 91060 401628 278412 401656
rect 91060 401616 91066 401628
rect 278406 401616 278412 401628
rect 278464 401616 278470 401668
rect 90910 400188 90916 400240
rect 90968 400228 90974 400240
rect 278682 400228 278688 400240
rect 90968 400200 278688 400228
rect 90968 400188 90974 400200
rect 278682 400188 278688 400200
rect 278740 400188 278746 400240
rect 89622 397468 89628 397520
rect 89680 397508 89686 397520
rect 278682 397508 278688 397520
rect 89680 397480 278688 397508
rect 89680 397468 89686 397480
rect 278682 397468 278688 397480
rect 278740 397468 278746 397520
rect 88242 396040 88248 396092
rect 88300 396080 88306 396092
rect 278682 396080 278688 396092
rect 88300 396052 278688 396080
rect 88300 396040 88306 396052
rect 278682 396040 278688 396052
rect 278740 396040 278746 396092
rect 3142 395972 3148 396024
rect 3200 396012 3206 396024
rect 280062 396012 280068 396024
rect 3200 395984 280068 396012
rect 3200 395972 3206 395984
rect 280062 395972 280068 395984
rect 280120 395972 280126 396024
rect 86862 393320 86868 393372
rect 86920 393360 86926 393372
rect 278682 393360 278688 393372
rect 86920 393332 278688 393360
rect 86920 393320 86926 393332
rect 278682 393320 278688 393332
rect 278740 393320 278746 393372
rect 542170 393252 542176 393304
rect 542228 393292 542234 393304
rect 542354 393292 542360 393304
rect 542228 393264 542360 393292
rect 542228 393252 542234 393264
rect 542354 393252 542360 393264
rect 542412 393252 542418 393304
rect 523954 391960 523960 392012
rect 524012 392000 524018 392012
rect 579890 392000 579896 392012
rect 524012 391972 579896 392000
rect 524012 391960 524018 391972
rect 579890 391960 579896 391972
rect 579948 391960 579954 392012
rect 85482 390532 85488 390584
rect 85540 390572 85546 390584
rect 278314 390572 278320 390584
rect 85540 390544 278320 390572
rect 85540 390532 85546 390544
rect 278314 390532 278320 390544
rect 278372 390532 278378 390584
rect 84102 389172 84108 389224
rect 84160 389212 84166 389224
rect 278682 389212 278688 389224
rect 84160 389184 278688 389212
rect 84160 389172 84166 389184
rect 278682 389172 278688 389184
rect 278740 389172 278746 389224
rect 82722 386384 82728 386436
rect 82780 386424 82786 386436
rect 277854 386424 277860 386436
rect 82780 386396 277860 386424
rect 82780 386384 82786 386396
rect 277854 386384 277860 386396
rect 277912 386384 277918 386436
rect 82630 385024 82636 385076
rect 82688 385064 82694 385076
rect 277670 385064 277676 385076
rect 82688 385036 277676 385064
rect 82688 385024 82694 385036
rect 277670 385024 277676 385036
rect 277728 385024 277734 385076
rect 542170 383664 542176 383716
rect 542228 383704 542234 383716
rect 542446 383704 542452 383716
rect 542228 383676 542452 383704
rect 542228 383664 542234 383676
rect 542446 383664 542452 383676
rect 542504 383664 542510 383716
rect 81342 382236 81348 382288
rect 81400 382276 81406 382288
rect 278682 382276 278688 382288
rect 81400 382248 278688 382276
rect 81400 382236 81406 382248
rect 278682 382236 278688 382248
rect 278740 382236 278746 382288
rect 79962 380876 79968 380928
rect 80020 380916 80026 380928
rect 278038 380916 278044 380928
rect 80020 380888 278044 380916
rect 80020 380876 80026 380888
rect 278038 380876 278044 380888
rect 278096 380876 278102 380928
rect 3510 380808 3516 380860
rect 3568 380848 3574 380860
rect 279970 380848 279976 380860
rect 3568 380820 279976 380848
rect 3568 380808 3574 380820
rect 279970 380808 279976 380820
rect 280028 380808 280034 380860
rect 542446 379448 542452 379500
rect 542504 379488 542510 379500
rect 542630 379488 542636 379500
rect 542504 379460 542636 379488
rect 542504 379448 542510 379460
rect 542630 379448 542636 379460
rect 542688 379448 542694 379500
rect 78582 378156 78588 378208
rect 78640 378196 78646 378208
rect 278682 378196 278688 378208
rect 78640 378168 278688 378196
rect 78640 378156 78646 378168
rect 278682 378156 278688 378168
rect 278740 378156 278746 378208
rect 77202 376728 77208 376780
rect 77260 376768 77266 376780
rect 278682 376768 278688 376780
rect 77260 376740 278688 376768
rect 77260 376728 77266 376740
rect 278682 376728 278688 376740
rect 278740 376728 278746 376780
rect 75822 374008 75828 374060
rect 75880 374048 75886 374060
rect 278406 374048 278412 374060
rect 75880 374020 278412 374048
rect 75880 374008 75886 374020
rect 278406 374008 278412 374020
rect 278464 374008 278470 374060
rect 74442 372580 74448 372632
rect 74500 372620 74506 372632
rect 278038 372620 278044 372632
rect 74500 372592 278044 372620
rect 74500 372580 74506 372592
rect 278038 372580 278044 372592
rect 278096 372580 278102 372632
rect 73062 369860 73068 369912
rect 73120 369900 73126 369912
rect 278314 369900 278320 369912
rect 73120 369872 278320 369900
rect 73120 369860 73126 369872
rect 278314 369860 278320 369872
rect 278372 369860 278378 369912
rect 72970 368500 72976 368552
rect 73028 368540 73034 368552
rect 278682 368540 278688 368552
rect 73028 368512 278688 368540
rect 73028 368500 73034 368512
rect 278682 368500 278688 368512
rect 278740 368500 278746 368552
rect 3510 367004 3516 367056
rect 3568 367044 3574 367056
rect 279878 367044 279884 367056
rect 3568 367016 279884 367044
rect 3568 367004 3574 367016
rect 279878 367004 279884 367016
rect 279936 367004 279942 367056
rect 542446 367004 542452 367056
rect 542504 367044 542510 367056
rect 542722 367044 542728 367056
rect 542504 367016 542728 367044
rect 542504 367004 542510 367016
rect 542722 367004 542728 367016
rect 542780 367004 542786 367056
rect 71682 365712 71688 365764
rect 71740 365752 71746 365764
rect 278682 365752 278688 365764
rect 71740 365724 278688 365752
rect 71740 365712 71746 365724
rect 278682 365712 278688 365724
rect 278740 365712 278746 365764
rect 70302 362924 70308 362976
rect 70360 362964 70366 362976
rect 277854 362964 277860 362976
rect 70360 362936 277860 362964
rect 70360 362924 70366 362936
rect 277854 362924 277860 362936
rect 277912 362924 277918 362976
rect 68922 361564 68928 361616
rect 68980 361604 68986 361616
rect 278682 361604 278688 361616
rect 68980 361576 278688 361604
rect 68980 361564 68986 361576
rect 278682 361564 278688 361576
rect 278740 361564 278746 361616
rect 67542 358776 67548 358828
rect 67600 358816 67606 358828
rect 277854 358816 277860 358828
rect 67600 358788 277860 358816
rect 67600 358776 67606 358788
rect 277854 358776 277860 358788
rect 277912 358776 277918 358828
rect 66162 357416 66168 357468
rect 66220 357456 66226 357468
rect 278682 357456 278688 357468
rect 66220 357428 278688 357456
rect 66220 357416 66226 357428
rect 278682 357416 278688 357428
rect 278740 357416 278746 357468
rect 542446 357416 542452 357468
rect 542504 357456 542510 357468
rect 542538 357456 542544 357468
rect 542504 357428 542544 357456
rect 542504 357416 542510 357428
rect 542538 357416 542544 357428
rect 542596 357416 542602 357468
rect 64782 354696 64788 354748
rect 64840 354736 64846 354748
rect 278682 354736 278688 354748
rect 64840 354708 278688 354736
rect 64840 354696 64846 354708
rect 278682 354696 278688 354708
rect 278740 354696 278746 354748
rect 64690 353268 64696 353320
rect 64748 353308 64754 353320
rect 278038 353308 278044 353320
rect 64748 353280 278044 353308
rect 64748 353268 64754 353280
rect 278038 353268 278044 353280
rect 278096 353268 278102 353320
rect 63402 350548 63408 350600
rect 63460 350588 63466 350600
rect 278682 350588 278688 350600
rect 63460 350560 278688 350588
rect 63460 350548 63466 350560
rect 278682 350548 278688 350560
rect 278740 350548 278746 350600
rect 542538 350548 542544 350600
rect 542596 350548 542602 350600
rect 542556 350520 542584 350548
rect 542722 350520 542728 350532
rect 542556 350492 542728 350520
rect 542722 350480 542728 350492
rect 542780 350480 542786 350532
rect 62022 349120 62028 349172
rect 62080 349160 62086 349172
rect 278682 349160 278688 349172
rect 62080 349132 278688 349160
rect 62080 349120 62086 349132
rect 278682 349120 278688 349132
rect 278740 349120 278746 349172
rect 60642 346400 60648 346452
rect 60700 346440 60706 346452
rect 278682 346440 278688 346452
rect 60700 346412 278688 346440
rect 60700 346400 60706 346412
rect 278682 346400 278688 346412
rect 278740 346400 278746 346452
rect 59262 345040 59268 345092
rect 59320 345080 59326 345092
rect 278682 345080 278688 345092
rect 59320 345052 278688 345080
rect 59320 345040 59326 345052
rect 278682 345040 278688 345052
rect 278740 345040 278746 345092
rect 57882 342252 57888 342304
rect 57940 342292 57946 342304
rect 278314 342292 278320 342304
rect 57940 342264 278320 342292
rect 57940 342252 57946 342264
rect 278314 342252 278320 342264
rect 278372 342252 278378 342304
rect 56502 340892 56508 340944
rect 56560 340932 56566 340944
rect 278682 340932 278688 340944
rect 56560 340904 278688 340932
rect 56560 340892 56566 340904
rect 278682 340892 278688 340904
rect 278740 340892 278746 340944
rect 522942 340824 522948 340876
rect 523000 340864 523006 340876
rect 542722 340864 542728 340876
rect 523000 340836 542728 340864
rect 523000 340824 523006 340836
rect 542722 340824 542728 340836
rect 542780 340824 542786 340876
rect 56410 338104 56416 338156
rect 56468 338144 56474 338156
rect 278682 338144 278688 338156
rect 56468 338116 278688 338144
rect 56468 338104 56474 338116
rect 278682 338104 278688 338116
rect 278740 338104 278746 338156
rect 3510 338036 3516 338088
rect 3568 338076 3574 338088
rect 279786 338076 279792 338088
rect 3568 338048 279792 338076
rect 3568 338036 3574 338048
rect 279786 338036 279792 338048
rect 279844 338036 279850 338088
rect 522942 337900 522948 337952
rect 523000 337940 523006 337952
rect 527174 337940 527180 337952
rect 523000 337912 527180 337940
rect 523000 337900 523006 337912
rect 527174 337900 527180 337912
rect 527232 337900 527238 337952
rect 522574 336676 522580 336728
rect 522632 336716 522638 336728
rect 531958 336716 531964 336728
rect 522632 336688 531964 336716
rect 522632 336676 522638 336688
rect 531958 336676 531964 336688
rect 532016 336676 532022 336728
rect 55122 335316 55128 335368
rect 55180 335356 55186 335368
rect 277854 335356 277860 335368
rect 55180 335328 277860 335356
rect 55180 335316 55186 335328
rect 277854 335316 277860 335328
rect 277912 335316 277918 335368
rect 53742 333956 53748 334008
rect 53800 333996 53806 334008
rect 278682 333996 278688 334008
rect 53800 333968 278688 333996
rect 53800 333956 53806 333968
rect 278682 333956 278688 333968
rect 278740 333956 278746 334008
rect 522942 333888 522948 333940
rect 523000 333928 523006 333940
rect 560938 333928 560944 333940
rect 523000 333900 560944 333928
rect 523000 333888 523006 333900
rect 560938 333888 560944 333900
rect 560996 333888 561002 333940
rect 522574 332528 522580 332580
rect 522632 332568 522638 332580
rect 545758 332568 545764 332580
rect 522632 332540 545764 332568
rect 522632 332528 522638 332540
rect 545758 332528 545764 332540
rect 545816 332528 545822 332580
rect 52362 331236 52368 331288
rect 52420 331276 52426 331288
rect 278682 331276 278688 331288
rect 52420 331248 278688 331276
rect 52420 331236 52426 331248
rect 278682 331236 278688 331248
rect 278740 331236 278746 331288
rect 50982 329808 50988 329860
rect 51040 329848 51046 329860
rect 278682 329848 278688 329860
rect 51040 329820 278688 329848
rect 51040 329808 51046 329820
rect 278682 329808 278688 329820
rect 278740 329808 278746 329860
rect 522942 328516 522948 328568
rect 523000 328556 523006 328568
rect 529198 328556 529204 328568
rect 523000 328528 529204 328556
rect 523000 328516 523006 328528
rect 529198 328516 529204 328528
rect 529256 328516 529262 328568
rect 522942 328380 522948 328432
rect 523000 328420 523006 328432
rect 558178 328420 558184 328432
rect 523000 328392 558184 328420
rect 523000 328380 523006 328392
rect 558178 328380 558184 328392
rect 558236 328380 558242 328432
rect 49602 327088 49608 327140
rect 49660 327128 49666 327140
rect 278682 327128 278688 327140
rect 49660 327100 278688 327128
rect 49660 327088 49666 327100
rect 278682 327088 278688 327100
rect 278740 327088 278746 327140
rect 48222 325660 48228 325712
rect 48280 325700 48286 325712
rect 278038 325700 278044 325712
rect 48280 325672 278044 325700
rect 48280 325660 48286 325672
rect 278038 325660 278044 325672
rect 278096 325660 278102 325712
rect 522942 325592 522948 325644
rect 523000 325632 523006 325644
rect 540238 325632 540244 325644
rect 523000 325604 540244 325632
rect 523000 325592 523006 325604
rect 540238 325592 540244 325604
rect 540296 325592 540302 325644
rect 3510 324232 3516 324284
rect 3568 324272 3574 324284
rect 279694 324272 279700 324284
rect 3568 324244 279700 324272
rect 3568 324232 3574 324244
rect 279694 324232 279700 324244
rect 279752 324232 279758 324284
rect 522298 324096 522304 324148
rect 522356 324136 522362 324148
rect 525058 324136 525064 324148
rect 522356 324108 525064 324136
rect 522356 324096 522362 324108
rect 525058 324096 525064 324108
rect 525116 324096 525122 324148
rect 48130 322940 48136 322992
rect 48188 322980 48194 322992
rect 277670 322980 277676 322992
rect 48188 322952 277676 322980
rect 48188 322940 48194 322952
rect 277670 322940 277676 322952
rect 277728 322940 277734 322992
rect 46842 321580 46848 321632
rect 46900 321620 46906 321632
rect 278038 321620 278044 321632
rect 46900 321592 278044 321620
rect 46900 321580 46906 321592
rect 278038 321580 278044 321592
rect 278096 321580 278102 321632
rect 522666 321512 522672 321564
rect 522724 321552 522730 321564
rect 556798 321552 556804 321564
rect 522724 321524 556804 321552
rect 522724 321512 522730 321524
rect 556798 321512 556804 321524
rect 556856 321512 556862 321564
rect 522942 320084 522948 320136
rect 523000 320124 523006 320136
rect 538858 320124 538864 320136
rect 523000 320096 538864 320124
rect 523000 320084 523006 320096
rect 538858 320084 538864 320096
rect 538916 320084 538922 320136
rect 45462 318792 45468 318844
rect 45520 318832 45526 318844
rect 278682 318832 278688 318844
rect 45520 318804 278688 318832
rect 45520 318792 45526 318804
rect 278682 318792 278688 318804
rect 278740 318792 278746 318844
rect 44082 317432 44088 317484
rect 44140 317472 44146 317484
rect 278682 317472 278688 317484
rect 44140 317444 278688 317472
rect 44140 317432 44146 317444
rect 278682 317432 278688 317444
rect 278740 317432 278746 317484
rect 522298 316888 522304 316940
rect 522356 316928 522362 316940
rect 523678 316928 523684 316940
rect 522356 316900 523684 316928
rect 522356 316888 522362 316900
rect 523678 316888 523684 316900
rect 523736 316888 523742 316940
rect 42702 314644 42708 314696
rect 42760 314684 42766 314696
rect 278682 314684 278688 314696
rect 42760 314656 278688 314684
rect 42760 314644 42766 314656
rect 278682 314644 278688 314656
rect 278740 314644 278746 314696
rect 522942 314576 522948 314628
rect 523000 314616 523006 314628
rect 555418 314616 555424 314628
rect 523000 314588 555424 314616
rect 523000 314576 523006 314588
rect 555418 314576 555424 314588
rect 555476 314576 555482 314628
rect 41322 313284 41328 313336
rect 41380 313324 41386 313336
rect 278682 313324 278688 313336
rect 41380 313296 278688 313324
rect 41380 313284 41386 313296
rect 278682 313284 278688 313296
rect 278740 313284 278746 313336
rect 522942 313216 522948 313268
rect 523000 313256 523006 313268
rect 537478 313256 537484 313268
rect 523000 313228 537484 313256
rect 523000 313216 523006 313228
rect 537478 313216 537484 313228
rect 537536 313216 537542 313268
rect 39942 310496 39948 310548
rect 40000 310536 40006 310548
rect 278682 310536 278688 310548
rect 40000 310508 278688 310536
rect 40000 310496 40006 310508
rect 278682 310496 278688 310508
rect 278740 310496 278746 310548
rect 522298 310428 522304 310480
rect 522356 310468 522362 310480
rect 523770 310468 523776 310480
rect 522356 310440 523776 310468
rect 522356 310428 522362 310440
rect 523770 310428 523776 310440
rect 523828 310428 523834 310480
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 279602 309108 279608 309120
rect 3384 309080 279608 309108
rect 3384 309068 3390 309080
rect 279602 309068 279608 309080
rect 279660 309068 279666 309120
rect 522942 309068 522948 309120
rect 523000 309108 523006 309120
rect 554038 309108 554044 309120
rect 523000 309080 554044 309108
rect 523000 309068 523006 309080
rect 554038 309068 554044 309080
rect 554096 309068 554102 309120
rect 38562 307776 38568 307828
rect 38620 307816 38626 307828
rect 277854 307816 277860 307828
rect 38620 307788 277860 307816
rect 38620 307776 38626 307788
rect 277854 307776 277860 307788
rect 277912 307776 277918 307828
rect 38470 306348 38476 306400
rect 38528 306388 38534 306400
rect 278682 306388 278688 306400
rect 38528 306360 278688 306388
rect 38528 306348 38534 306360
rect 278682 306348 278688 306360
rect 278740 306348 278746 306400
rect 522942 306280 522948 306332
rect 523000 306320 523006 306332
rect 536098 306320 536104 306332
rect 523000 306292 536104 306320
rect 523000 306280 523006 306292
rect 536098 306280 536104 306292
rect 536156 306280 536162 306332
rect 522298 304784 522304 304836
rect 522356 304824 522362 304836
rect 523862 304824 523868 304836
rect 522356 304796 523868 304824
rect 522356 304784 522362 304796
rect 523862 304784 523868 304796
rect 523920 304784 523926 304836
rect 37182 303628 37188 303680
rect 37240 303668 37246 303680
rect 278682 303668 278688 303680
rect 37240 303640 278688 303668
rect 37240 303628 37246 303640
rect 278682 303628 278688 303640
rect 278740 303628 278746 303680
rect 35802 302200 35808 302252
rect 35860 302240 35866 302252
rect 278682 302240 278688 302252
rect 35860 302212 278688 302240
rect 35860 302200 35866 302212
rect 278682 302200 278688 302212
rect 278740 302200 278746 302252
rect 522942 302132 522948 302184
rect 523000 302172 523006 302184
rect 563698 302172 563704 302184
rect 523000 302144 563704 302172
rect 523000 302132 523006 302144
rect 563698 302132 563704 302144
rect 563756 302132 563762 302184
rect 522942 300772 522948 300824
rect 523000 300812 523006 300824
rect 549898 300812 549904 300824
rect 523000 300784 549904 300812
rect 523000 300772 523006 300784
rect 549898 300772 549904 300784
rect 549956 300772 549962 300824
rect 34422 299480 34428 299532
rect 34480 299520 34486 299532
rect 278682 299520 278688 299532
rect 34480 299492 278688 299520
rect 34480 299480 34486 299492
rect 278682 299480 278688 299492
rect 278740 299480 278746 299532
rect 33042 298120 33048 298172
rect 33100 298160 33106 298172
rect 278682 298160 278688 298172
rect 33100 298132 278688 298160
rect 33100 298120 33106 298132
rect 278682 298120 278688 298132
rect 278740 298120 278746 298172
rect 522942 298052 522948 298104
rect 523000 298092 523006 298104
rect 534718 298092 534724 298104
rect 523000 298064 534724 298092
rect 523000 298052 523006 298064
rect 534718 298052 534724 298064
rect 534776 298052 534782 298104
rect 522942 296624 522948 296676
rect 523000 296664 523006 296676
rect 580258 296664 580264 296676
rect 523000 296636 580264 296664
rect 523000 296624 523006 296636
rect 580258 296624 580264 296636
rect 580316 296624 580322 296676
rect 31662 295332 31668 295384
rect 31720 295372 31726 295384
rect 278682 295372 278688 295384
rect 31720 295344 278688 295372
rect 31720 295332 31726 295344
rect 278682 295332 278688 295344
rect 278740 295332 278746 295384
rect 3050 295264 3056 295316
rect 3108 295304 3114 295316
rect 279510 295304 279516 295316
rect 3108 295276 279516 295304
rect 3108 295264 3114 295276
rect 279510 295264 279516 295276
rect 279568 295264 279574 295316
rect 522482 294652 522488 294704
rect 522540 294692 522546 294704
rect 580718 294692 580724 294704
rect 522540 294664 580724 294692
rect 522540 294652 522546 294664
rect 580718 294652 580724 294664
rect 580776 294652 580782 294704
rect 522298 294584 522304 294636
rect 522356 294624 522362 294636
rect 579982 294624 579988 294636
rect 522356 294596 579988 294624
rect 522356 294584 522362 294596
rect 579982 294584 579988 294596
rect 580040 294584 580046 294636
rect 30282 293972 30288 294024
rect 30340 294012 30346 294024
rect 278682 294012 278688 294024
rect 30340 293984 278688 294012
rect 30340 293972 30346 293984
rect 278682 293972 278688 293984
rect 278740 293972 278746 294024
rect 522942 293904 522948 293956
rect 523000 293944 523006 293956
rect 547138 293944 547144 293956
rect 523000 293916 547144 293944
rect 523000 293904 523006 293916
rect 547138 293904 547144 293916
rect 547196 293904 547202 293956
rect 522574 292000 522580 292052
rect 522632 292040 522638 292052
rect 523954 292040 523960 292052
rect 522632 292012 523960 292040
rect 522632 292000 522638 292012
rect 523954 292000 523960 292012
rect 524012 292000 524018 292052
rect 30190 291184 30196 291236
rect 30248 291224 30254 291236
rect 278682 291224 278688 291236
rect 30248 291196 278688 291224
rect 30248 291184 30254 291196
rect 278682 291184 278688 291196
rect 278740 291184 278746 291236
rect 28902 289824 28908 289876
rect 28960 289864 28966 289876
rect 278682 289864 278688 289876
rect 28960 289836 278688 289864
rect 28960 289824 28966 289836
rect 278682 289824 278688 289836
rect 278740 289824 278746 289876
rect 522942 289756 522948 289808
rect 523000 289796 523006 289808
rect 580442 289796 580448 289808
rect 523000 289768 580448 289796
rect 523000 289756 523006 289768
rect 580442 289756 580448 289768
rect 580500 289756 580506 289808
rect 522574 288328 522580 288380
rect 522632 288368 522638 288380
rect 580350 288368 580356 288380
rect 522632 288340 580356 288368
rect 522632 288328 522638 288340
rect 580350 288328 580356 288340
rect 580408 288328 580414 288380
rect 27522 287036 27528 287088
rect 27580 287076 27586 287088
rect 278682 287076 278688 287088
rect 27580 287048 278688 287076
rect 27580 287036 27586 287048
rect 278682 287036 278688 287048
rect 278740 287036 278746 287088
rect 26142 285676 26148 285728
rect 26200 285716 26206 285728
rect 278682 285716 278688 285728
rect 26200 285688 278688 285716
rect 26200 285676 26206 285688
rect 278682 285676 278688 285688
rect 278740 285676 278746 285728
rect 522574 285608 522580 285660
rect 522632 285648 522638 285660
rect 580534 285648 580540 285660
rect 522632 285620 580540 285648
rect 522632 285608 522638 285620
rect 580534 285608 580540 285620
rect 580592 285608 580598 285660
rect 24762 282888 24768 282940
rect 24820 282928 24826 282940
rect 278682 282928 278688 282940
rect 24820 282900 278688 282928
rect 24820 282888 24826 282900
rect 278682 282888 278688 282900
rect 278740 282888 278746 282940
rect 522942 281460 522948 281512
rect 523000 281500 523006 281512
rect 580626 281500 580632 281512
rect 523000 281472 580632 281500
rect 523000 281460 523006 281472
rect 580626 281460 580632 281472
rect 580684 281460 580690 281512
rect 23382 280168 23388 280220
rect 23440 280208 23446 280220
rect 277854 280208 277860 280220
rect 23440 280180 277860 280208
rect 23440 280168 23446 280180
rect 277854 280168 277860 280180
rect 277912 280168 277918 280220
rect 3510 280100 3516 280152
rect 3568 280140 3574 280152
rect 279418 280140 279424 280152
rect 3568 280112 279424 280140
rect 3568 280100 3574 280112
rect 279418 280100 279424 280112
rect 279476 280100 279482 280152
rect 22002 278740 22008 278792
rect 22060 278780 22066 278792
rect 278682 278780 278688 278792
rect 22060 278752 278688 278780
rect 22060 278740 22066 278752
rect 278682 278740 278688 278752
rect 278740 278740 278746 278792
rect 21910 276020 21916 276072
rect 21968 276060 21974 276072
rect 278682 276060 278688 276072
rect 21968 276032 278688 276060
rect 21968 276020 21974 276032
rect 278682 276020 278688 276032
rect 278740 276020 278746 276072
rect 522942 275272 522948 275324
rect 523000 275312 523006 275324
rect 580166 275312 580172 275324
rect 523000 275284 580172 275312
rect 523000 275272 523006 275284
rect 580166 275272 580172 275284
rect 580224 275272 580230 275324
rect 20622 274660 20628 274712
rect 20680 274700 20686 274712
rect 278038 274700 278044 274712
rect 20680 274672 278044 274700
rect 20680 274660 20686 274672
rect 278038 274660 278044 274672
rect 278096 274660 278102 274712
rect 19242 271872 19248 271924
rect 19300 271912 19306 271924
rect 278682 271912 278688 271924
rect 19300 271884 278688 271912
rect 19300 271872 19306 271884
rect 278682 271872 278688 271884
rect 278740 271872 278746 271924
rect 17862 270512 17868 270564
rect 17920 270552 17926 270564
rect 278682 270552 278688 270564
rect 17920 270524 278688 270552
rect 17920 270512 17926 270524
rect 278682 270512 278688 270524
rect 278740 270512 278746 270564
rect 16482 267724 16488 267776
rect 16540 267764 16546 267776
rect 278682 267764 278688 267776
rect 16540 267736 278688 267764
rect 16540 267724 16546 267736
rect 278682 267724 278688 267736
rect 278740 267724 278746 267776
rect 15102 266364 15108 266416
rect 15160 266404 15166 266416
rect 278038 266404 278044 266416
rect 15160 266376 278044 266404
rect 15160 266364 15166 266376
rect 278038 266364 278044 266376
rect 278096 266364 278102 266416
rect 522482 265616 522488 265668
rect 522540 265656 522546 265668
rect 580166 265656 580172 265668
rect 522540 265628 580172 265656
rect 522540 265616 522546 265628
rect 580166 265616 580172 265628
rect 580224 265616 580230 265668
rect 522574 264936 522580 264988
rect 522632 264976 522638 264988
rect 523954 264976 523960 264988
rect 522632 264948 523960 264976
rect 522632 264936 522638 264948
rect 523954 264936 523960 264948
rect 524012 264936 524018 264988
rect 13722 263576 13728 263628
rect 13780 263616 13786 263628
rect 278682 263616 278688 263628
rect 13780 263588 278688 263616
rect 13780 263576 13786 263588
rect 278682 263576 278688 263588
rect 278740 263576 278746 263628
rect 13630 262216 13636 262268
rect 13688 262256 13694 262268
rect 278682 262256 278688 262268
rect 13688 262228 278688 262256
rect 13688 262216 13694 262228
rect 278682 262216 278688 262228
rect 278740 262216 278746 262268
rect 522574 260856 522580 260908
rect 522632 260896 522638 260908
rect 523862 260896 523868 260908
rect 522632 260868 523868 260896
rect 522632 260856 522638 260868
rect 523862 260856 523868 260868
rect 523920 260856 523926 260908
rect 12342 259428 12348 259480
rect 12400 259468 12406 259480
rect 278314 259468 278320 259480
rect 12400 259440 278320 259468
rect 12400 259428 12406 259440
rect 278314 259428 278320 259440
rect 278372 259428 278378 259480
rect 522574 259428 522580 259480
rect 522632 259468 522638 259480
rect 523770 259468 523776 259480
rect 522632 259440 523776 259468
rect 522632 259428 522638 259440
rect 523770 259428 523776 259440
rect 523828 259428 523834 259480
rect 10962 256708 10968 256760
rect 11020 256748 11026 256760
rect 277854 256748 277860 256760
rect 11020 256720 277860 256748
rect 11020 256708 11026 256720
rect 277854 256708 277860 256720
rect 277912 256708 277918 256760
rect 9582 255280 9588 255332
rect 9640 255320 9646 255332
rect 278682 255320 278688 255332
rect 9640 255292 278688 255320
rect 9640 255280 9646 255292
rect 278682 255280 278688 255292
rect 278740 255280 278746 255332
rect 8202 252560 8208 252612
rect 8260 252600 8266 252612
rect 277854 252600 277860 252612
rect 8260 252572 277860 252600
rect 8260 252560 8266 252572
rect 277854 252560 277860 252572
rect 277912 252560 277918 252612
rect 522298 252492 522304 252544
rect 522356 252532 522362 252544
rect 579798 252532 579804 252544
rect 522356 252504 579804 252532
rect 522356 252492 522362 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 6822 251200 6828 251252
rect 6880 251240 6886 251252
rect 278682 251240 278688 251252
rect 6880 251212 278688 251240
rect 6880 251200 6886 251212
rect 278682 251200 278688 251212
rect 278740 251200 278746 251252
rect 5442 248412 5448 248464
rect 5500 248452 5506 248464
rect 278682 248452 278688 248464
rect 5500 248424 278688 248452
rect 5500 248412 5506 248424
rect 278682 248412 278688 248424
rect 278740 248412 278746 248464
rect 522298 248412 522304 248464
rect 522356 248452 522362 248464
rect 531958 248452 531964 248464
rect 522356 248424 531964 248452
rect 522356 248412 522362 248424
rect 531958 248412 531964 248424
rect 532016 248412 532022 248464
rect 522298 247052 522304 247104
rect 522356 247092 522362 247104
rect 527818 247092 527824 247104
rect 522356 247064 527824 247092
rect 522356 247052 522362 247064
rect 527818 247052 527824 247064
rect 527876 247052 527882 247104
rect 522390 243176 522396 243228
rect 522448 243176 522454 243228
rect 522408 243012 522436 243176
rect 522316 242984 522436 243012
rect 2682 242904 2688 242956
rect 2740 242944 2746 242956
rect 277394 242944 277400 242956
rect 2740 242916 277400 242944
rect 2740 242904 2746 242916
rect 277394 242904 277400 242916
rect 277452 242904 277458 242956
rect 522316 242808 522344 242984
rect 522390 242904 522396 242956
rect 522448 242944 522454 242956
rect 529198 242944 529204 242956
rect 522448 242916 529204 242944
rect 522448 242904 522454 242916
rect 529198 242904 529204 242916
rect 529256 242904 529262 242956
rect 522390 242808 522396 242820
rect 522316 242780 522396 242808
rect 522390 242768 522396 242780
rect 522448 242768 522454 242820
rect 3510 240864 3516 240916
rect 3568 240904 3574 240916
rect 522390 240904 522396 240916
rect 3568 240876 522396 240904
rect 3568 240864 3574 240876
rect 522390 240864 522396 240876
rect 522448 240864 522454 240916
rect 3602 240796 3608 240848
rect 3660 240836 3666 240848
rect 519814 240836 519820 240848
rect 3660 240808 519820 240836
rect 3660 240796 3666 240808
rect 519814 240796 519820 240808
rect 519872 240796 519878 240848
rect 292500 240740 306420 240768
rect 280154 240660 280160 240712
rect 280212 240700 280218 240712
rect 280890 240700 280896 240712
rect 280212 240672 280896 240700
rect 280212 240660 280218 240672
rect 280890 240660 280896 240672
rect 280948 240700 280954 240712
rect 292500 240700 292528 240740
rect 306392 240712 306420 240740
rect 367020 240740 369716 240768
rect 280948 240672 292528 240700
rect 280948 240660 280954 240672
rect 306374 240660 306380 240712
rect 306432 240660 306438 240712
rect 315942 240660 315948 240712
rect 316000 240700 316006 240712
rect 316000 240672 316080 240700
rect 316000 240660 316006 240672
rect 316052 240644 316080 240672
rect 325602 240660 325608 240712
rect 325660 240700 325666 240712
rect 325660 240672 335308 240700
rect 325660 240660 325666 240672
rect 316034 240592 316040 240644
rect 316092 240592 316098 240644
rect 335280 240632 335308 240672
rect 340874 240660 340880 240712
rect 340932 240700 340938 240712
rect 350442 240700 350448 240712
rect 340932 240672 350448 240700
rect 340932 240660 340938 240672
rect 350442 240660 350448 240672
rect 350500 240660 350506 240712
rect 340782 240632 340788 240644
rect 335280 240604 340788 240632
rect 340782 240592 340788 240604
rect 340840 240592 340846 240644
rect 350626 240592 350632 240644
rect 350684 240632 350690 240644
rect 357434 240632 357440 240644
rect 350684 240604 357440 240632
rect 350684 240592 350690 240604
rect 357434 240592 357440 240604
rect 357492 240592 357498 240644
rect 360378 240592 360384 240644
rect 360436 240632 360442 240644
rect 367020 240632 367048 240740
rect 369688 240712 369716 240740
rect 369670 240660 369676 240712
rect 369728 240660 369734 240712
rect 360436 240604 367048 240632
rect 360436 240592 360442 240604
rect 306374 240456 306380 240508
rect 306432 240496 306438 240508
rect 315942 240496 315948 240508
rect 306432 240468 315948 240496
rect 306432 240456 306438 240468
rect 315942 240456 315948 240468
rect 316000 240456 316006 240508
rect 369670 240388 369676 240440
rect 369728 240428 369734 240440
rect 373258 240428 373264 240440
rect 369728 240400 373264 240428
rect 369728 240388 369734 240400
rect 373258 240388 373264 240400
rect 373316 240388 373322 240440
rect 1302 240116 1308 240168
rect 1360 240156 1366 240168
rect 278682 240156 278688 240168
rect 1360 240128 278688 240156
rect 1360 240116 1366 240128
rect 278682 240116 278688 240128
rect 278740 240116 278746 240168
rect 522390 240116 522396 240168
rect 522448 240156 522454 240168
rect 525058 240156 525064 240168
rect 522448 240128 525064 240156
rect 522448 240116 522454 240128
rect 525058 240116 525064 240128
rect 525116 240116 525122 240168
rect 333698 238688 333704 238740
rect 333756 238728 333762 238740
rect 344554 238728 344560 238740
rect 333756 238700 344560 238728
rect 333756 238688 333762 238700
rect 344554 238688 344560 238700
rect 344612 238688 344618 238740
rect 426342 238688 426348 238740
rect 426400 238728 426406 238740
rect 450538 238728 450544 238740
rect 426400 238700 450544 238728
rect 426400 238688 426406 238700
rect 450538 238688 450544 238700
rect 450596 238688 450602 238740
rect 459462 238688 459468 238740
rect 459520 238728 459526 238740
rect 473998 238728 474004 238740
rect 459520 238700 474004 238728
rect 459520 238688 459526 238700
rect 473998 238688 474004 238700
rect 474056 238688 474062 238740
rect 475562 238688 475568 238740
rect 475620 238728 475626 238740
rect 489914 238728 489920 238740
rect 475620 238700 489920 238728
rect 475620 238688 475626 238700
rect 489914 238688 489920 238700
rect 489972 238688 489978 238740
rect 332502 238620 332508 238672
rect 332560 238660 332566 238672
rect 346762 238660 346768 238672
rect 332560 238632 346768 238660
rect 332560 238620 332566 238632
rect 346762 238620 346768 238632
rect 346820 238620 346826 238672
rect 424410 238620 424416 238672
rect 424468 238660 424474 238672
rect 452010 238660 452016 238672
rect 424468 238632 452016 238660
rect 424468 238620 424474 238632
rect 452010 238620 452016 238632
rect 452068 238620 452074 238672
rect 463602 238620 463608 238672
rect 463660 238660 463666 238672
rect 492030 238660 492036 238672
rect 463660 238632 492036 238660
rect 463660 238620 463666 238632
rect 492030 238620 492036 238632
rect 492088 238620 492094 238672
rect 331122 238552 331128 238604
rect 331180 238592 331186 238604
rect 349154 238592 349160 238604
rect 331180 238564 349160 238592
rect 331180 238552 331186 238564
rect 349154 238552 349160 238564
rect 349212 238552 349218 238604
rect 422202 238552 422208 238604
rect 422260 238592 422266 238604
rect 453298 238592 453304 238604
rect 422260 238564 453304 238592
rect 422260 238552 422266 238564
rect 453298 238552 453304 238564
rect 453356 238552 453362 238604
rect 462222 238552 462228 238604
rect 462280 238592 462286 238604
rect 494238 238592 494244 238604
rect 462280 238564 494244 238592
rect 462280 238552 462286 238564
rect 494238 238552 494244 238564
rect 494296 238552 494302 238604
rect 329558 238484 329564 238536
rect 329616 238524 329622 238536
rect 351086 238524 351092 238536
rect 329616 238496 351092 238524
rect 329616 238484 329622 238496
rect 351086 238484 351092 238496
rect 351144 238484 351150 238536
rect 380434 238484 380440 238536
rect 380492 238524 380498 238536
rect 395154 238524 395160 238536
rect 380492 238496 395160 238524
rect 380492 238484 380498 238496
rect 395154 238484 395160 238496
rect 395212 238484 395218 238536
rect 417878 238484 417884 238536
rect 417936 238524 417942 238536
rect 456242 238524 456248 238536
rect 417936 238496 456248 238524
rect 417936 238484 417942 238496
rect 456242 238484 456248 238496
rect 456300 238484 456306 238536
rect 459462 238484 459468 238536
rect 459520 238524 459526 238536
rect 498654 238524 498660 238536
rect 459520 238496 498660 238524
rect 459520 238484 459526 238496
rect 498654 238484 498660 238496
rect 498712 238484 498718 238536
rect 294506 238416 294512 238468
rect 294564 238456 294570 238468
rect 295242 238456 295248 238468
rect 294564 238428 295248 238456
rect 294564 238416 294570 238428
rect 295242 238416 295248 238428
rect 295300 238416 295306 238468
rect 328362 238416 328368 238468
rect 328420 238456 328426 238468
rect 353294 238456 353300 238468
rect 328420 238428 353300 238456
rect 328420 238416 328426 238428
rect 353294 238416 353300 238428
rect 353352 238416 353358 238468
rect 380342 238416 380348 238468
rect 380400 238456 380406 238468
rect 397454 238456 397460 238468
rect 380400 238428 397460 238456
rect 380400 238416 380406 238428
rect 397454 238416 397460 238428
rect 397512 238416 397518 238468
rect 415302 238416 415308 238468
rect 415360 238456 415366 238468
rect 456058 238456 456064 238468
rect 415360 238428 456064 238456
rect 415360 238416 415366 238428
rect 456058 238416 456064 238428
rect 456116 238416 456122 238468
rect 456702 238416 456708 238468
rect 456760 238456 456766 238468
rect 503070 238456 503076 238468
rect 456760 238428 503076 238456
rect 456760 238416 456766 238428
rect 503070 238416 503076 238428
rect 503128 238416 503134 238468
rect 311802 238348 311808 238400
rect 311860 238388 311866 238400
rect 342898 238388 342904 238400
rect 311860 238360 342904 238388
rect 311860 238348 311866 238360
rect 342898 238348 342904 238360
rect 342956 238348 342962 238400
rect 380250 238348 380256 238400
rect 380308 238388 380314 238400
rect 399570 238388 399576 238400
rect 380308 238360 399576 238388
rect 380308 238348 380314 238360
rect 399570 238348 399576 238360
rect 399628 238348 399634 238400
rect 419994 238348 420000 238400
rect 420052 238388 420058 238400
rect 454678 238388 454684 238400
rect 420052 238360 454684 238388
rect 420052 238348 420058 238360
rect 454678 238348 454684 238360
rect 454736 238348 454742 238400
rect 455138 238348 455144 238400
rect 455196 238388 455202 238400
rect 507486 238388 507492 238400
rect 455196 238360 507492 238388
rect 455196 238348 455202 238360
rect 507486 238348 507492 238360
rect 507544 238348 507550 238400
rect 309962 238280 309968 238332
rect 310020 238320 310026 238332
rect 344278 238320 344284 238332
rect 310020 238292 344284 238320
rect 310020 238280 310026 238292
rect 344278 238280 344284 238292
rect 344336 238280 344342 238332
rect 389082 238280 389088 238332
rect 389140 238320 389146 238332
rect 451918 238320 451924 238332
rect 389140 238292 451924 238320
rect 389140 238280 389146 238292
rect 451918 238280 451924 238292
rect 451976 238280 451982 238332
rect 452562 238280 452568 238332
rect 452620 238320 452626 238332
rect 512086 238320 512092 238332
rect 452620 238292 512092 238320
rect 452620 238280 452626 238292
rect 512086 238280 512092 238292
rect 512144 238280 512150 238332
rect 305546 238212 305552 238264
rect 305604 238252 305610 238264
rect 342990 238252 342996 238264
rect 305604 238224 342996 238252
rect 305604 238212 305610 238224
rect 342990 238212 342996 238224
rect 343048 238212 343054 238264
rect 371142 238212 371148 238264
rect 371200 238252 371206 238264
rect 390738 238252 390744 238264
rect 371200 238224 390744 238252
rect 371200 238212 371206 238224
rect 390738 238212 390744 238224
rect 390796 238212 390802 238264
rect 395338 238212 395344 238264
rect 395396 238252 395402 238264
rect 406194 238252 406200 238264
rect 395396 238224 406200 238252
rect 395396 238212 395402 238224
rect 406194 238212 406200 238224
rect 406252 238212 406258 238264
rect 428826 238212 428832 238264
rect 428884 238252 428890 238264
rect 449158 238252 449164 238264
rect 428884 238224 449164 238252
rect 428884 238212 428890 238224
rect 449158 238212 449164 238224
rect 449216 238212 449222 238264
rect 449802 238212 449808 238264
rect 449860 238252 449866 238264
rect 516318 238252 516324 238264
rect 449860 238224 516324 238252
rect 449860 238212 449866 238224
rect 516318 238212 516324 238224
rect 516376 238212 516382 238264
rect 283466 238144 283472 238196
rect 283524 238184 283530 238196
rect 297818 238184 297824 238196
rect 283524 238156 297824 238184
rect 283524 238144 283530 238156
rect 297818 238144 297824 238156
rect 297876 238144 297882 238196
rect 303338 238144 303344 238196
rect 303396 238184 303402 238196
rect 341518 238184 341524 238196
rect 303396 238156 341524 238184
rect 303396 238144 303402 238156
rect 341518 238144 341524 238156
rect 341576 238144 341582 238196
rect 380526 238144 380532 238196
rect 380584 238184 380590 238196
rect 412818 238184 412824 238196
rect 380584 238156 412824 238184
rect 380584 238144 380590 238156
rect 412818 238144 412824 238156
rect 412876 238144 412882 238196
rect 431034 238144 431040 238196
rect 431092 238184 431098 238196
rect 447778 238184 447784 238196
rect 431092 238156 447784 238184
rect 431092 238144 431098 238156
rect 447778 238144 447784 238156
rect 447836 238144 447842 238196
rect 448422 238144 448428 238196
rect 448480 238184 448486 238196
rect 518526 238184 518532 238196
rect 448480 238156 518532 238184
rect 448480 238144 448486 238156
rect 518526 238144 518532 238156
rect 518584 238144 518590 238196
rect 281350 238076 281356 238128
rect 281408 238116 281414 238128
rect 297358 238116 297364 238128
rect 281408 238088 297364 238116
rect 281408 238076 281414 238088
rect 297358 238076 297364 238088
rect 297416 238076 297422 238128
rect 307662 238076 307668 238128
rect 307720 238116 307726 238128
rect 347038 238116 347044 238128
rect 307720 238088 347044 238116
rect 307720 238076 307726 238088
rect 347038 238076 347044 238088
rect 347096 238076 347102 238128
rect 380158 238076 380164 238128
rect 380216 238116 380222 238128
rect 403986 238116 403992 238128
rect 380216 238088 403992 238116
rect 380216 238076 380222 238088
rect 403986 238076 403992 238088
rect 404044 238076 404050 238128
rect 411162 238076 411168 238128
rect 411220 238116 411226 238128
rect 496354 238116 496360 238128
rect 411220 238088 496360 238116
rect 411220 238076 411226 238088
rect 496354 238076 496360 238088
rect 496412 238076 496418 238128
rect 285582 238008 285588 238060
rect 285640 238048 285646 238060
rect 345658 238048 345664 238060
rect 285640 238020 345664 238048
rect 285640 238008 285646 238020
rect 345658 238008 345664 238020
rect 345716 238008 345722 238060
rect 360562 238008 360568 238060
rect 360620 238048 360626 238060
rect 476758 238048 476764 238060
rect 360620 238020 476764 238048
rect 360620 238008 360626 238020
rect 476758 238008 476764 238020
rect 476816 238008 476822 238060
rect 461854 237940 461860 237992
rect 461912 237980 461918 237992
rect 474090 237980 474096 237992
rect 461912 237952 474096 237980
rect 461912 237940 461918 237952
rect 474090 237940 474096 237952
rect 474148 237940 474154 237992
rect 475470 237940 475476 237992
rect 475528 237980 475534 237992
rect 487614 237980 487620 237992
rect 475528 237952 487620 237980
rect 475528 237940 475534 237952
rect 487614 237940 487620 237952
rect 487672 237940 487678 237992
rect 464062 237872 464068 237924
rect 464120 237912 464126 237924
rect 475378 237912 475384 237924
rect 464120 237884 475384 237912
rect 464120 237872 464126 237884
rect 475378 237872 475384 237884
rect 475436 237872 475442 237924
rect 335170 237804 335176 237856
rect 335228 237844 335234 237856
rect 342346 237844 342352 237856
rect 335228 237816 342352 237844
rect 335228 237804 335234 237816
rect 342346 237804 342352 237816
rect 342404 237804 342410 237856
rect 470502 237804 470508 237856
rect 470560 237844 470566 237856
rect 473354 237844 473360 237856
rect 470560 237816 473360 237844
rect 470560 237804 470566 237816
rect 473354 237804 473360 237816
rect 473412 237804 473418 237856
rect 474274 237804 474280 237856
rect 474332 237844 474338 237856
rect 485774 237844 485780 237856
rect 474332 237816 485780 237844
rect 474332 237804 474338 237816
rect 485774 237804 485780 237816
rect 485832 237804 485838 237856
rect 466270 237736 466276 237788
rect 466328 237776 466334 237788
rect 475654 237776 475660 237788
rect 466328 237748 475660 237776
rect 466328 237736 466334 237748
rect 475654 237736 475660 237748
rect 475712 237736 475718 237788
rect 331950 237668 331956 237720
rect 332008 237708 332014 237720
rect 339586 237708 339592 237720
rect 332008 237680 339592 237708
rect 332008 237668 332014 237680
rect 339586 237668 339592 237680
rect 339644 237668 339650 237720
rect 474182 237668 474188 237720
rect 474240 237708 474246 237720
rect 483290 237708 483296 237720
rect 474240 237680 483296 237708
rect 474240 237668 474246 237680
rect 483290 237668 483296 237680
rect 483348 237668 483354 237720
rect 335262 237600 335268 237652
rect 335320 237640 335326 237652
rect 340138 237640 340144 237652
rect 335320 237612 340144 237640
rect 335320 237600 335326 237612
rect 340138 237600 340144 237612
rect 340196 237600 340202 237652
rect 468478 237600 468484 237652
rect 468536 237640 468542 237652
rect 474826 237640 474832 237652
rect 468536 237612 474832 237640
rect 468536 237600 468542 237612
rect 474826 237600 474832 237612
rect 474884 237600 474890 237652
rect 333882 237532 333888 237584
rect 333940 237572 333946 237584
rect 338206 237572 338212 237584
rect 333940 237544 338212 237572
rect 333940 237532 333946 237544
rect 338206 237532 338212 237544
rect 338264 237532 338270 237584
rect 337378 237504 337384 237516
rect 331416 237476 337384 237504
rect 287882 237396 287888 237448
rect 287940 237436 287946 237448
rect 288342 237436 288348 237448
rect 287940 237408 288348 237436
rect 287940 237396 287946 237408
rect 288342 237396 288348 237408
rect 288400 237396 288406 237448
rect 298922 237396 298928 237448
rect 298980 237436 298986 237448
rect 299382 237436 299388 237448
rect 298980 237408 299388 237436
rect 298980 237396 298986 237408
rect 299382 237396 299388 237408
rect 299440 237396 299446 237448
rect 316494 237396 316500 237448
rect 316552 237436 316558 237448
rect 317322 237436 317328 237448
rect 316552 237408 317328 237436
rect 316552 237396 316558 237408
rect 317322 237396 317328 237408
rect 317380 237396 317386 237448
rect 320910 237396 320916 237448
rect 320968 237436 320974 237448
rect 321462 237436 321468 237448
rect 320968 237408 321468 237436
rect 320968 237396 320974 237408
rect 321462 237396 321468 237408
rect 321520 237396 321526 237448
rect 327534 237396 327540 237448
rect 327592 237436 327598 237448
rect 328270 237436 328276 237448
rect 327592 237408 328276 237436
rect 327592 237396 327598 237408
rect 328270 237396 328276 237408
rect 328328 237396 328334 237448
rect 329742 237396 329748 237448
rect 329800 237436 329806 237448
rect 331416 237436 331444 237476
rect 337378 237464 337384 237476
rect 337436 237464 337442 237516
rect 367002 237464 367008 237516
rect 367060 237504 367066 237516
rect 371234 237504 371240 237516
rect 367060 237476 371240 237504
rect 367060 237464 367066 237476
rect 371234 237464 371240 237476
rect 371292 237464 371298 237516
rect 329800 237408 331444 237436
rect 329800 237396 329806 237408
rect 333698 237396 333704 237448
rect 333756 237436 333762 237448
rect 333882 237436 333888 237448
rect 333756 237408 333888 237436
rect 333756 237396 333762 237408
rect 333882 237396 333888 237408
rect 333940 237396 333946 237448
rect 336550 237396 336556 237448
rect 336608 237436 336614 237448
rect 338114 237436 338120 237448
rect 336608 237408 338120 237436
rect 336608 237396 336614 237408
rect 338114 237396 338120 237408
rect 338172 237396 338178 237448
rect 364978 237396 364984 237448
rect 365036 237436 365042 237448
rect 366358 237436 366364 237448
rect 365036 237408 366364 237436
rect 365036 237396 365042 237408
rect 366358 237396 366364 237408
rect 366416 237396 366422 237448
rect 366910 237396 366916 237448
rect 366968 237436 366974 237448
rect 368750 237436 368756 237448
rect 366968 237408 368756 237436
rect 366968 237396 366974 237408
rect 368750 237396 368756 237408
rect 368808 237396 368814 237448
rect 376018 237396 376024 237448
rect 376076 237436 376082 237448
rect 376662 237436 376668 237448
rect 376076 237408 376668 237436
rect 376076 237396 376082 237408
rect 376662 237396 376668 237408
rect 376720 237396 376726 237448
rect 382642 237396 382648 237448
rect 382700 237436 382706 237448
rect 383562 237436 383568 237448
rect 382700 237408 383568 237436
rect 382700 237396 382706 237408
rect 383562 237396 383568 237408
rect 383620 237396 383626 237448
rect 386966 237396 386972 237448
rect 387024 237436 387030 237448
rect 387702 237436 387708 237448
rect 387024 237408 387708 237436
rect 387024 237396 387030 237408
rect 387702 237396 387708 237408
rect 387760 237396 387766 237448
rect 391198 237396 391204 237448
rect 391256 237436 391262 237448
rect 392946 237436 392952 237448
rect 391256 237408 392952 237436
rect 391256 237396 391262 237408
rect 392946 237396 392952 237408
rect 393004 237396 393010 237448
rect 393958 237396 393964 237448
rect 394016 237436 394022 237448
rect 401778 237436 401784 237448
rect 394016 237408 401784 237436
rect 394016 237396 394022 237408
rect 401778 237396 401784 237408
rect 401836 237396 401842 237448
rect 453022 237396 453028 237448
rect 453080 237436 453086 237448
rect 453942 237436 453948 237448
rect 453080 237408 453948 237436
rect 453080 237396 453086 237408
rect 453942 237396 453948 237408
rect 454000 237396 454006 237448
rect 457438 237396 457444 237448
rect 457496 237436 457502 237448
rect 458082 237436 458088 237448
rect 457496 237408 458088 237436
rect 457496 237396 457502 237408
rect 458082 237396 458088 237408
rect 458140 237396 458146 237448
rect 471882 237396 471888 237448
rect 471940 237436 471946 237448
rect 474734 237436 474740 237448
rect 471940 237408 474740 237436
rect 471940 237396 471946 237408
rect 474734 237396 474740 237408
rect 474792 237396 474798 237448
rect 3510 237328 3516 237380
rect 3568 237368 3574 237380
rect 522114 237368 522120 237380
rect 3568 237340 522120 237368
rect 3568 237328 3574 237340
rect 522114 237328 522120 237340
rect 522172 237328 522178 237380
rect 329558 234540 329564 234592
rect 329616 234580 329622 234592
rect 329742 234580 329748 234592
rect 329616 234552 329748 234580
rect 329616 234540 329622 234552
rect 329742 234540 329748 234552
rect 329800 234540 329806 234592
rect 431954 232160 431960 232212
rect 432012 232200 432018 232212
rect 432690 232200 432696 232212
rect 432012 232172 432696 232200
rect 432012 232160 432018 232172
rect 432690 232160 432696 232172
rect 432748 232160 432754 232212
rect 336366 230460 336372 230512
rect 336424 230500 336430 230512
rect 336550 230500 336556 230512
rect 336424 230472 336556 230500
rect 336424 230460 336430 230472
rect 336550 230460 336556 230472
rect 336608 230460 336614 230512
rect 522942 229032 522948 229084
rect 523000 229072 523006 229084
rect 580166 229072 580172 229084
rect 523000 229044 580172 229072
rect 523000 229032 523006 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 522206 223564 522212 223576
rect 3200 223536 522212 223564
rect 3200 223524 3206 223536
rect 522206 223524 522212 223536
rect 522264 223524 522270 223576
rect 336366 222232 336372 222284
rect 336424 222272 336430 222284
rect 336642 222272 336648 222284
rect 336424 222244 336648 222272
rect 336424 222232 336430 222244
rect 336642 222232 336648 222244
rect 336700 222232 336706 222284
rect 329466 222164 329472 222216
rect 329524 222204 329530 222216
rect 329650 222204 329656 222216
rect 329524 222176 329656 222204
rect 329524 222164 329530 222176
rect 329650 222164 329656 222176
rect 329708 222164 329714 222216
rect 431770 222164 431776 222216
rect 431828 222204 431834 222216
rect 432046 222204 432052 222216
rect 431828 222176 432052 222204
rect 431828 222164 431834 222176
rect 432046 222164 432052 222176
rect 432104 222164 432110 222216
rect 522850 217948 522856 218000
rect 522908 217988 522914 218000
rect 580166 217988 580172 218000
rect 522908 217960 580172 217988
rect 522908 217948 522914 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 432046 215364 432052 215416
rect 432104 215364 432110 215416
rect 432064 215336 432092 215364
rect 432138 215336 432144 215348
rect 432064 215308 432144 215336
rect 432138 215296 432144 215308
rect 432196 215296 432202 215348
rect 3510 208292 3516 208344
rect 3568 208332 3574 208344
rect 522022 208332 522028 208344
rect 3568 208304 522028 208332
rect 3568 208292 3574 208304
rect 522022 208292 522028 208304
rect 522080 208292 522086 208344
rect 523954 205572 523960 205624
rect 524012 205612 524018 205624
rect 579798 205612 579804 205624
rect 524012 205584 579804 205612
rect 524012 205572 524018 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 470502 205232 470508 205284
rect 470560 205272 470566 205284
rect 476114 205272 476120 205284
rect 470560 205244 476120 205272
rect 470560 205232 470566 205244
rect 476114 205232 476120 205244
rect 476172 205232 476178 205284
rect 470410 205096 470416 205148
rect 470468 205136 470474 205148
rect 478874 205136 478880 205148
rect 470468 205108 478880 205136
rect 470468 205096 470474 205108
rect 478874 205096 478880 205108
rect 478932 205096 478938 205148
rect 469122 205028 469128 205080
rect 469180 205068 469186 205080
rect 480254 205068 480260 205080
rect 469180 205040 480260 205068
rect 469180 205028 469186 205040
rect 480254 205028 480260 205040
rect 480312 205028 480318 205080
rect 451182 204960 451188 205012
rect 451240 205000 451246 205012
rect 484394 205000 484400 205012
rect 451240 204972 484400 205000
rect 451240 204960 451246 204972
rect 484394 204960 484400 204972
rect 484452 204960 484458 205012
rect 373902 204892 373908 204944
rect 373960 204932 373966 204944
rect 490190 204932 490196 204944
rect 373960 204904 490196 204932
rect 373960 204892 373966 204904
rect 490190 204892 490196 204904
rect 490248 204892 490254 204944
rect 347774 204280 347780 204332
rect 347832 204320 347838 204332
rect 357342 204320 357348 204332
rect 347832 204292 357348 204320
rect 347832 204280 347838 204292
rect 357342 204280 357348 204292
rect 357400 204280 357406 204332
rect 389818 204280 389824 204332
rect 389876 204320 389882 204332
rect 394418 204320 394424 204332
rect 389876 204292 394424 204320
rect 389876 204280 389882 204292
rect 394418 204280 394424 204292
rect 394476 204280 394482 204332
rect 317322 204212 317328 204264
rect 317380 204252 317386 204264
rect 342806 204252 342812 204264
rect 317380 204224 342812 204252
rect 317380 204212 317386 204224
rect 342806 204212 342812 204224
rect 342864 204212 342870 204264
rect 342916 204224 344508 204252
rect 299382 204144 299388 204196
rect 299440 204184 299446 204196
rect 342916 204184 342944 204224
rect 299440 204156 342944 204184
rect 344480 204184 344508 204224
rect 347038 204212 347044 204264
rect 347096 204252 347102 204264
rect 351914 204252 351920 204264
rect 347096 204224 351920 204252
rect 347096 204212 347102 204224
rect 351914 204212 351920 204224
rect 351972 204212 351978 204264
rect 374638 204212 374644 204264
rect 374696 204252 374702 204264
rect 379514 204252 379520 204264
rect 374696 204224 379520 204252
rect 374696 204212 374702 204224
rect 379514 204212 379520 204224
rect 379572 204212 379578 204264
rect 416038 204212 416044 204264
rect 416096 204252 416102 204264
rect 427814 204252 427820 204264
rect 416096 204224 427820 204252
rect 416096 204212 416102 204224
rect 427814 204212 427820 204224
rect 427872 204212 427878 204264
rect 452010 204212 452016 204264
rect 452068 204252 452074 204264
rect 461486 204252 461492 204264
rect 452068 204224 461492 204252
rect 452068 204212 452074 204224
rect 461486 204212 461492 204224
rect 461544 204212 461550 204264
rect 464982 204212 464988 204264
rect 465040 204252 465046 204264
rect 475470 204252 475476 204264
rect 465040 204224 475476 204252
rect 465040 204212 465046 204224
rect 475470 204212 475476 204224
rect 475528 204212 475534 204264
rect 476758 204212 476764 204264
rect 476816 204252 476822 204264
rect 485774 204252 485780 204264
rect 476816 204224 485780 204252
rect 476816 204212 476822 204224
rect 485774 204212 485780 204224
rect 485832 204212 485838 204264
rect 357434 204184 357440 204196
rect 344480 204156 357440 204184
rect 299440 204144 299446 204156
rect 357434 204144 357440 204156
rect 357492 204144 357498 204196
rect 357986 204144 357992 204196
rect 358044 204184 358050 204196
rect 394510 204184 394516 204196
rect 358044 204156 394516 204184
rect 358044 204144 358050 204156
rect 394510 204144 394516 204156
rect 394568 204144 394574 204196
rect 394602 204144 394608 204196
rect 394660 204184 394666 204196
rect 412542 204184 412548 204196
rect 394660 204156 412548 204184
rect 394660 204144 394666 204156
rect 412542 204144 412548 204156
rect 412600 204144 412606 204196
rect 412634 204144 412640 204196
rect 412692 204184 412698 204196
rect 445754 204184 445760 204196
rect 412692 204156 445760 204184
rect 412692 204144 412698 204156
rect 445754 204144 445760 204156
rect 445812 204144 445818 204196
rect 450538 204144 450544 204196
rect 450596 204184 450602 204196
rect 450906 204184 450912 204196
rect 450596 204156 450912 204184
rect 450596 204144 450602 204156
rect 450906 204144 450912 204156
rect 450964 204184 450970 204196
rect 460658 204184 460664 204196
rect 450964 204156 460664 204184
rect 450964 204144 450970 204156
rect 460658 204144 460664 204156
rect 460716 204144 460722 204196
rect 466270 204144 466276 204196
rect 466328 204184 466334 204196
rect 474274 204184 474280 204196
rect 466328 204156 474280 204184
rect 466328 204144 466334 204156
rect 474274 204144 474280 204156
rect 474332 204144 474338 204196
rect 475378 204144 475384 204196
rect 475436 204184 475442 204196
rect 477494 204184 477500 204196
rect 475436 204156 477500 204184
rect 475436 204144 475442 204156
rect 477494 204144 477500 204156
rect 477552 204144 477558 204196
rect 330938 204076 330944 204128
rect 330996 204116 331002 204128
rect 337286 204116 337292 204128
rect 330996 204088 337292 204116
rect 330996 204076 331002 204088
rect 337286 204076 337292 204088
rect 337344 204076 337350 204128
rect 337378 204076 337384 204128
rect 337436 204116 337442 204128
rect 340966 204116 340972 204128
rect 337436 204088 340972 204116
rect 337436 204076 337442 204088
rect 340966 204076 340972 204088
rect 341024 204076 341030 204128
rect 342806 204076 342812 204128
rect 342864 204116 342870 204128
rect 347774 204116 347780 204128
rect 342864 204088 347780 204116
rect 342864 204076 342870 204088
rect 347774 204076 347780 204088
rect 347832 204076 347838 204128
rect 354030 204076 354036 204128
rect 354088 204116 354094 204128
rect 358630 204116 358636 204128
rect 354088 204088 358636 204116
rect 354088 204076 354094 204088
rect 358630 204076 358636 204088
rect 358688 204116 358694 204128
rect 364978 204116 364984 204128
rect 358688 204088 364984 204116
rect 358688 204076 358694 204088
rect 364978 204076 364984 204088
rect 365036 204076 365042 204128
rect 367094 204076 367100 204128
rect 367152 204116 367158 204128
rect 376570 204116 376576 204128
rect 367152 204088 376576 204116
rect 367152 204076 367158 204088
rect 376570 204076 376576 204088
rect 376628 204076 376634 204128
rect 379514 204076 379520 204128
rect 379572 204116 379578 204128
rect 389818 204116 389824 204128
rect 379572 204088 389824 204116
rect 379572 204076 379578 204088
rect 389818 204076 389824 204088
rect 389876 204076 389882 204128
rect 394418 204076 394424 204128
rect 394476 204116 394482 204128
rect 402882 204116 402888 204128
rect 394476 204088 402888 204116
rect 394476 204076 394482 204088
rect 402882 204076 402888 204088
rect 402940 204076 402946 204128
rect 402974 204076 402980 204128
rect 403032 204116 403038 204128
rect 416038 204116 416044 204128
rect 403032 204088 416044 204116
rect 403032 204076 403038 204088
rect 416038 204076 416044 204088
rect 416096 204076 416102 204128
rect 427906 204076 427912 204128
rect 427964 204116 427970 204128
rect 442994 204116 443000 204128
rect 427964 204088 443000 204116
rect 427964 204076 427970 204088
rect 442994 204076 443000 204088
rect 443052 204076 443058 204128
rect 449158 204076 449164 204128
rect 449216 204116 449222 204128
rect 459094 204116 459100 204128
rect 449216 204088 459100 204116
rect 449216 204076 449222 204088
rect 459094 204076 459100 204088
rect 459152 204076 459158 204128
rect 467282 204076 467288 204128
rect 467340 204116 467346 204128
rect 475746 204116 475752 204128
rect 467340 204088 475752 204116
rect 467340 204076 467346 204088
rect 475746 204076 475752 204088
rect 475804 204076 475810 204128
rect 475838 204076 475844 204128
rect 475896 204116 475902 204128
rect 483014 204116 483020 204128
rect 475896 204088 483020 204116
rect 475896 204076 475902 204088
rect 483014 204076 483020 204088
rect 483072 204076 483078 204128
rect 300762 204008 300768 204060
rect 300820 204048 300826 204060
rect 356054 204048 356060 204060
rect 300820 204020 356060 204048
rect 300820 204008 300826 204020
rect 356054 204008 356060 204020
rect 356112 204008 356118 204060
rect 360010 204008 360016 204060
rect 360068 204048 360074 204060
rect 441614 204048 441620 204060
rect 360068 204020 441620 204048
rect 360068 204008 360074 204020
rect 441614 204008 441620 204020
rect 441672 204008 441678 204060
rect 447778 204008 447784 204060
rect 447836 204048 447842 204060
rect 448422 204048 448428 204060
rect 447836 204020 448428 204048
rect 447836 204008 447842 204020
rect 448422 204008 448428 204020
rect 448480 204048 448486 204060
rect 457898 204048 457904 204060
rect 448480 204020 457904 204048
rect 448480 204008 448486 204020
rect 457898 204008 457904 204020
rect 457956 204008 457962 204060
rect 457990 204008 457996 204060
rect 458048 204048 458054 204060
rect 500954 204048 500960 204060
rect 458048 204020 500960 204048
rect 458048 204008 458054 204020
rect 500954 204008 500960 204020
rect 501012 204008 501018 204060
rect 314562 203940 314568 203992
rect 314620 203980 314626 203992
rect 349154 203980 349160 203992
rect 314620 203952 349160 203980
rect 314620 203940 314626 203952
rect 349154 203940 349160 203952
rect 349212 203940 349218 203992
rect 361298 203980 361304 203992
rect 356532 203952 361304 203980
rect 333790 203872 333796 203924
rect 333848 203912 333854 203924
rect 341702 203912 341708 203924
rect 333848 203884 341708 203912
rect 333848 203872 333854 203884
rect 341702 203872 341708 203884
rect 341760 203872 341766 203924
rect 349430 203912 349436 203924
rect 345124 203884 349436 203912
rect 318702 203804 318708 203856
rect 318760 203844 318766 203856
rect 335078 203844 335084 203856
rect 318760 203816 335084 203844
rect 318760 203804 318766 203816
rect 335078 203804 335084 203816
rect 335136 203804 335142 203856
rect 345014 203844 345020 203856
rect 335188 203816 345020 203844
rect 321462 203736 321468 203788
rect 321520 203776 321526 203788
rect 335188 203776 335216 203816
rect 345014 203804 345020 203816
rect 345072 203804 345078 203856
rect 321520 203748 335216 203776
rect 321520 203736 321526 203748
rect 335814 203736 335820 203788
rect 335872 203776 335878 203788
rect 335872 203748 337240 203776
rect 335872 203736 335878 203748
rect 322842 203668 322848 203720
rect 322900 203708 322906 203720
rect 335998 203708 336004 203720
rect 322900 203680 336004 203708
rect 322900 203668 322906 203680
rect 335998 203668 336004 203680
rect 336056 203668 336062 203720
rect 337212 203708 337240 203748
rect 337286 203736 337292 203788
rect 337344 203776 337350 203788
rect 340046 203776 340052 203788
rect 337344 203748 340052 203776
rect 337344 203736 337350 203748
rect 340046 203736 340052 203748
rect 340104 203776 340110 203788
rect 345124 203776 345152 203884
rect 349430 203872 349436 203884
rect 349488 203912 349494 203924
rect 354030 203912 354036 203924
rect 349488 203884 354036 203912
rect 349488 203872 349494 203884
rect 354030 203872 354036 203884
rect 354088 203872 354094 203924
rect 356532 203912 356560 203952
rect 361298 203940 361304 203952
rect 361356 203980 361362 203992
rect 438854 203980 438860 203992
rect 361356 203952 438860 203980
rect 361356 203940 361362 203952
rect 438854 203940 438860 203952
rect 438912 203940 438918 203992
rect 460842 203940 460848 203992
rect 460900 203980 460906 203992
rect 495434 203980 495440 203992
rect 460900 203952 495440 203980
rect 460900 203940 460906 203952
rect 495434 203940 495440 203952
rect 495492 203940 495498 203992
rect 354232 203884 356560 203912
rect 345566 203804 345572 203856
rect 345624 203844 345630 203856
rect 351638 203844 351644 203856
rect 345624 203816 351644 203844
rect 345624 203804 345630 203816
rect 351638 203804 351644 203816
rect 351696 203844 351702 203856
rect 354232 203844 354260 203884
rect 362862 203872 362868 203924
rect 362920 203912 362926 203924
rect 436094 203912 436100 203924
rect 362920 203884 436100 203912
rect 362920 203872 362926 203884
rect 436094 203872 436100 203884
rect 436152 203872 436158 203924
rect 453942 203872 453948 203924
rect 454000 203912 454006 203924
rect 483014 203912 483020 203924
rect 454000 203884 483020 203912
rect 454000 203872 454006 203884
rect 483014 203872 483020 203884
rect 483072 203872 483078 203924
rect 351696 203816 354260 203844
rect 351696 203804 351702 203816
rect 354582 203804 354588 203856
rect 354640 203844 354646 203856
rect 363414 203844 363420 203856
rect 354640 203816 363420 203844
rect 354640 203804 354646 203816
rect 363414 203804 363420 203816
rect 363472 203844 363478 203856
rect 434714 203844 434720 203856
rect 363472 203816 434720 203844
rect 363472 203804 363478 203816
rect 434714 203804 434720 203816
rect 434772 203804 434778 203856
rect 455230 203804 455236 203856
rect 455288 203844 455294 203856
rect 471054 203844 471060 203856
rect 455288 203816 471060 203844
rect 455288 203804 455294 203816
rect 471054 203804 471060 203816
rect 471112 203804 471118 203856
rect 474090 203804 474096 203856
rect 474148 203844 474154 203856
rect 477494 203844 477500 203856
rect 474148 203816 477500 203844
rect 474148 203804 474154 203816
rect 477494 203804 477500 203816
rect 477552 203804 477558 203856
rect 340104 203748 345152 203776
rect 340104 203736 340110 203748
rect 345658 203736 345664 203788
rect 345716 203776 345722 203788
rect 364334 203776 364340 203788
rect 345716 203748 364340 203776
rect 345716 203736 345722 203748
rect 364334 203736 364340 203748
rect 364392 203736 364398 203788
rect 432138 203776 432144 203788
rect 418172 203748 432144 203776
rect 337930 203708 337936 203720
rect 337212 203680 337936 203708
rect 337930 203668 337936 203680
rect 337988 203708 337994 203720
rect 340690 203708 340696 203720
rect 337988 203680 340696 203708
rect 337988 203668 337994 203680
rect 340690 203668 340696 203680
rect 340748 203668 340754 203720
rect 342254 203708 342260 203720
rect 340800 203680 342260 203708
rect 325602 203600 325608 203652
rect 325660 203640 325666 203652
rect 331214 203640 331220 203652
rect 325660 203612 331220 203640
rect 325660 203600 325666 203612
rect 331214 203600 331220 203612
rect 331272 203600 331278 203652
rect 340598 203600 340604 203652
rect 340656 203640 340662 203652
rect 340800 203640 340828 203680
rect 342254 203668 342260 203680
rect 342312 203668 342318 203720
rect 342806 203668 342812 203720
rect 342864 203708 342870 203720
rect 343634 203708 343640 203720
rect 342864 203680 343640 203708
rect 342864 203668 342870 203680
rect 343634 203668 343640 203680
rect 343692 203708 343698 203720
rect 353018 203708 353024 203720
rect 343692 203680 353024 203708
rect 343692 203668 343698 203680
rect 353018 203668 353024 203680
rect 353076 203708 353082 203720
rect 362862 203708 362868 203720
rect 353076 203680 362868 203708
rect 353076 203668 353082 203680
rect 362862 203668 362868 203680
rect 362920 203668 362926 203720
rect 408586 203708 408592 203720
rect 402992 203680 408592 203708
rect 340656 203612 340828 203640
rect 340656 203600 340662 203612
rect 341518 203600 341524 203652
rect 341576 203640 341582 203652
rect 354674 203640 354680 203652
rect 341576 203612 354680 203640
rect 341576 203600 341582 203612
rect 354674 203600 354680 203612
rect 354732 203600 354738 203652
rect 355594 203600 355600 203652
rect 355652 203640 355658 203652
rect 365070 203640 365076 203652
rect 355652 203612 365076 203640
rect 355652 203600 355658 203612
rect 365070 203600 365076 203612
rect 365128 203640 365134 203652
rect 369854 203640 369860 203652
rect 365128 203612 369860 203640
rect 365128 203600 365134 203612
rect 369854 203600 369860 203612
rect 369912 203600 369918 203652
rect 376294 203600 376300 203652
rect 376352 203640 376358 203652
rect 402992 203640 403020 203680
rect 408586 203668 408592 203680
rect 408644 203668 408650 203720
rect 408678 203668 408684 203720
rect 408736 203708 408742 203720
rect 408736 203680 417464 203708
rect 408736 203668 408742 203680
rect 376352 203612 385080 203640
rect 376352 203600 376358 203612
rect 328270 203532 328276 203584
rect 328328 203572 328334 203584
rect 342254 203572 342260 203584
rect 328328 203544 342260 203572
rect 328328 203532 328334 203544
rect 342254 203532 342260 203544
rect 342312 203532 342318 203584
rect 342714 203532 342720 203584
rect 342772 203572 342778 203584
rect 348418 203572 348424 203584
rect 342772 203544 348424 203572
rect 342772 203532 342778 203544
rect 348418 203532 348424 203544
rect 348476 203572 348482 203584
rect 357986 203572 357992 203584
rect 348476 203544 357992 203572
rect 348476 203532 348482 203544
rect 357986 203532 357992 203544
rect 358044 203532 358050 203584
rect 364978 203532 364984 203584
rect 365036 203572 365042 203584
rect 374638 203572 374644 203584
rect 365036 203544 374644 203572
rect 365036 203532 365042 203544
rect 374638 203532 374644 203544
rect 374696 203532 374702 203584
rect 385052 203572 385080 203612
rect 394620 203612 403020 203640
rect 417436 203640 417464 203680
rect 418172 203640 418200 203748
rect 432138 203736 432144 203748
rect 432196 203736 432202 203788
rect 458082 203736 458088 203788
rect 458140 203776 458146 203788
rect 470778 203776 470784 203788
rect 458140 203748 470784 203776
rect 458140 203736 458146 203748
rect 470778 203736 470784 203748
rect 470836 203736 470842 203788
rect 471330 203736 471336 203788
rect 471388 203776 471394 203788
rect 474366 203776 474372 203788
rect 471388 203748 474372 203776
rect 471388 203736 471394 203748
rect 474366 203736 474372 203748
rect 474424 203736 474430 203788
rect 474458 203736 474464 203788
rect 474516 203776 474522 203788
rect 475838 203776 475844 203788
rect 474516 203748 475844 203776
rect 474516 203736 474522 203748
rect 475838 203736 475844 203748
rect 475896 203736 475902 203788
rect 463510 203668 463516 203720
rect 463568 203708 463574 203720
rect 470502 203708 470508 203720
rect 463568 203680 470508 203708
rect 463568 203668 463574 203680
rect 470502 203668 470508 203680
rect 470560 203668 470566 203720
rect 473906 203708 473912 203720
rect 470612 203680 473912 203708
rect 417436 203612 418200 203640
rect 394620 203572 394648 203612
rect 456702 203600 456708 203652
rect 456760 203640 456766 203652
rect 464706 203640 464712 203652
rect 456760 203612 464712 203640
rect 456760 203600 456766 203612
rect 464706 203600 464712 203612
rect 464764 203640 464770 203652
rect 470612 203640 470640 203680
rect 473906 203668 473912 203680
rect 473964 203668 473970 203720
rect 473998 203668 474004 203720
rect 474056 203708 474062 203720
rect 478874 203708 478880 203720
rect 474056 203680 478880 203708
rect 474056 203668 474062 203680
rect 478874 203668 478880 203680
rect 478932 203668 478938 203720
rect 464764 203612 470640 203640
rect 464764 203600 464770 203612
rect 470778 203600 470784 203652
rect 470836 203640 470842 203652
rect 480622 203640 480628 203652
rect 470836 203612 480628 203640
rect 470836 203600 470842 203612
rect 480622 203600 480628 203612
rect 480680 203600 480686 203652
rect 385052 203544 394648 203572
rect 456058 203532 456064 203584
rect 456116 203572 456122 203584
rect 465902 203572 465908 203584
rect 456116 203544 465908 203572
rect 456116 203532 456122 203544
rect 465902 203532 465908 203544
rect 465960 203572 465966 203584
rect 467282 203572 467288 203584
rect 465960 203544 467288 203572
rect 465960 203532 465966 203544
rect 467282 203532 467288 203544
rect 467340 203532 467346 203584
rect 470410 203572 470416 203584
rect 467392 203544 470416 203572
rect 335078 203464 335084 203516
rect 335136 203504 335142 203516
rect 346394 203504 346400 203516
rect 335136 203476 346400 203504
rect 335136 203464 335142 203476
rect 346394 203464 346400 203476
rect 346452 203464 346458 203516
rect 369854 203464 369860 203516
rect 369912 203504 369918 203516
rect 376294 203504 376300 203516
rect 369912 203476 376300 203504
rect 369912 203464 369918 203476
rect 376294 203464 376300 203476
rect 376352 203464 376358 203516
rect 461486 203464 461492 203516
rect 461544 203504 461550 203516
rect 467392 203504 467420 203544
rect 470410 203532 470416 203544
rect 470468 203532 470474 203584
rect 470686 203532 470692 203584
rect 470744 203572 470750 203584
rect 475562 203572 475568 203584
rect 470744 203544 475568 203572
rect 470744 203532 470750 203544
rect 475562 203532 475568 203544
rect 475620 203532 475626 203584
rect 475746 203532 475752 203584
rect 475804 203572 475810 203584
rect 484394 203572 484400 203584
rect 475804 203544 484400 203572
rect 475804 203532 475810 203544
rect 484394 203532 484400 203544
rect 484452 203532 484458 203584
rect 472894 203504 472900 203516
rect 461544 203476 467420 203504
rect 467484 203476 470548 203504
rect 461544 203464 461550 203476
rect 329742 203396 329748 203448
rect 329800 203436 329806 203448
rect 329800 203408 335952 203436
rect 329800 203396 329806 203408
rect 328270 203328 328276 203380
rect 328328 203368 328334 203380
rect 335814 203368 335820 203380
rect 328328 203340 335820 203368
rect 328328 203328 328334 203340
rect 335814 203328 335820 203340
rect 335872 203328 335878 203380
rect 335924 203368 335952 203408
rect 335998 203396 336004 203448
rect 336056 203436 336062 203448
rect 343634 203436 343640 203448
rect 336056 203408 343640 203436
rect 336056 203396 336062 203408
rect 343634 203396 343640 203408
rect 343692 203396 343698 203448
rect 344186 203396 344192 203448
rect 344244 203436 344250 203448
rect 347038 203436 347044 203448
rect 344244 203408 347044 203436
rect 344244 203396 344250 203408
rect 347038 203396 347044 203408
rect 347096 203436 347102 203448
rect 356422 203436 356428 203448
rect 347096 203408 356428 203436
rect 347096 203396 347102 203408
rect 356422 203396 356428 203408
rect 356480 203436 356486 203448
rect 447134 203436 447140 203448
rect 356480 203408 447140 203436
rect 356480 203396 356486 203408
rect 447134 203396 447140 203408
rect 447192 203396 447198 203448
rect 463050 203396 463056 203448
rect 463108 203436 463114 203448
rect 467484 203436 467512 203476
rect 463108 203408 467512 203436
rect 470520 203436 470548 203476
rect 470704 203476 472900 203504
rect 470704 203436 470732 203476
rect 472894 203464 472900 203476
rect 472952 203504 472958 203516
rect 472952 203476 479196 203504
rect 472952 203464 472958 203476
rect 470520 203408 470732 203436
rect 463108 203396 463114 203408
rect 471790 203396 471796 203448
rect 471848 203436 471854 203448
rect 479168 203436 479196 203476
rect 481634 203436 481640 203448
rect 471848 203408 479104 203436
rect 479168 203408 481640 203436
rect 471848 203396 471854 203408
rect 339218 203368 339224 203380
rect 335924 203340 339224 203368
rect 339218 203328 339224 203340
rect 339276 203368 339282 203380
rect 342714 203368 342720 203380
rect 339276 203340 342720 203368
rect 339276 203328 339282 203340
rect 342714 203328 342720 203340
rect 342772 203328 342778 203380
rect 342824 203340 349292 203368
rect 332410 203260 332416 203312
rect 332468 203300 332474 203312
rect 341334 203300 341340 203312
rect 332468 203272 341340 203300
rect 332468 203260 332474 203272
rect 341334 203260 341340 203272
rect 341392 203300 341398 203312
rect 342824 203300 342852 203340
rect 341392 203272 342852 203300
rect 341392 203260 341398 203272
rect 342898 203260 342904 203312
rect 342956 203300 342962 203312
rect 349154 203300 349160 203312
rect 342956 203272 349160 203300
rect 342956 203260 342962 203272
rect 349154 203260 349160 203272
rect 349212 203260 349218 203312
rect 349264 203300 349292 203340
rect 460658 203328 460664 203380
rect 460716 203368 460722 203380
rect 467558 203368 467564 203380
rect 460716 203340 467564 203368
rect 460716 203328 460722 203340
rect 467558 203328 467564 203340
rect 467616 203328 467622 203380
rect 467668 203340 474320 203368
rect 351178 203300 351184 203312
rect 349264 203272 351184 203300
rect 351178 203260 351184 203272
rect 351236 203260 351242 203312
rect 366358 203260 366364 203312
rect 366416 203300 366422 203312
rect 368474 203300 368480 203312
rect 366416 203272 368480 203300
rect 366416 203260 366422 203272
rect 368474 203260 368480 203272
rect 368532 203260 368538 203312
rect 457898 203260 457904 203312
rect 457956 203300 457962 203312
rect 467190 203300 467196 203312
rect 457956 203272 467196 203300
rect 457956 203260 457962 203272
rect 467190 203260 467196 203272
rect 467248 203300 467254 203312
rect 467668 203300 467696 203340
rect 467248 203272 467696 203300
rect 467248 203260 467254 203272
rect 467742 203260 467748 203312
rect 467800 203300 467806 203312
rect 474182 203300 474188 203312
rect 467800 203272 474188 203300
rect 467800 203260 467806 203272
rect 474182 203260 474188 203272
rect 474240 203260 474246 203312
rect 474292 203300 474320 203340
rect 474366 203328 474372 203380
rect 474424 203368 474430 203380
rect 478966 203368 478972 203380
rect 474424 203340 478972 203368
rect 474424 203328 474430 203340
rect 478966 203328 478972 203340
rect 479024 203328 479030 203380
rect 479076 203368 479104 203408
rect 481634 203396 481640 203408
rect 481692 203396 481698 203448
rect 480530 203368 480536 203380
rect 479076 203340 480536 203368
rect 480530 203328 480536 203340
rect 480588 203328 480594 203380
rect 476114 203300 476120 203312
rect 474292 203272 476120 203300
rect 476114 203260 476120 203272
rect 476172 203260 476178 203312
rect 331214 203192 331220 203244
rect 331272 203232 331278 203244
rect 331272 203204 331352 203232
rect 331272 203192 331278 203204
rect 331324 203164 331352 203204
rect 336550 203192 336556 203244
rect 336608 203232 336614 203244
rect 345934 203232 345940 203244
rect 336608 203204 345940 203232
rect 336608 203192 336614 203204
rect 345934 203192 345940 203204
rect 345992 203232 345998 203244
rect 355594 203232 355600 203244
rect 345992 203204 355600 203232
rect 345992 203192 345998 203204
rect 355594 203192 355600 203204
rect 355652 203192 355658 203244
rect 459094 203192 459100 203244
rect 459152 203232 459158 203244
rect 468478 203232 468484 203244
rect 459152 203204 468484 203232
rect 459152 203192 459158 203204
rect 468478 203192 468484 203204
rect 468536 203232 468542 203244
rect 477494 203232 477500 203244
rect 468536 203204 477500 203232
rect 468536 203192 468542 203204
rect 477494 203192 477500 203204
rect 477552 203192 477558 203244
rect 340598 203164 340604 203176
rect 331324 203136 340604 203164
rect 340598 203124 340604 203136
rect 340656 203124 340662 203176
rect 340782 203124 340788 203176
rect 340840 203164 340846 203176
rect 344186 203164 344192 203176
rect 340840 203136 344192 203164
rect 340840 203124 340846 203136
rect 344186 203124 344192 203136
rect 344244 203124 344250 203176
rect 344278 203124 344284 203176
rect 344336 203164 344342 203176
rect 351086 203164 351092 203176
rect 344336 203136 351092 203164
rect 344336 203124 344342 203136
rect 351086 203124 351092 203136
rect 351144 203124 351150 203176
rect 351178 203124 351184 203176
rect 351236 203164 351242 203176
rect 360010 203164 360016 203176
rect 351236 203136 360016 203164
rect 351236 203124 351242 203136
rect 360010 203124 360016 203136
rect 360068 203124 360074 203176
rect 453298 203124 453304 203176
rect 453356 203164 453362 203176
rect 462406 203164 462412 203176
rect 453356 203136 462412 203164
rect 453356 203124 453362 203136
rect 462406 203124 462412 203136
rect 462464 203164 462470 203176
rect 471054 203164 471060 203176
rect 462464 203136 471060 203164
rect 462464 203124 462470 203136
rect 471054 203124 471060 203136
rect 471112 203124 471118 203176
rect 471146 203124 471152 203176
rect 471204 203164 471210 203176
rect 481634 203164 481640 203176
rect 471204 203136 481640 203164
rect 471204 203124 471210 203136
rect 481634 203124 481640 203136
rect 481692 203124 481698 203176
rect 335262 203056 335268 203108
rect 335320 203096 335326 203108
rect 342806 203096 342812 203108
rect 335320 203068 342812 203096
rect 335320 203056 335326 203068
rect 342806 203056 342812 203068
rect 342864 203056 342870 203108
rect 342898 203056 342904 203108
rect 342956 203096 342962 203108
rect 344922 203096 344928 203108
rect 342956 203068 344928 203096
rect 342956 203056 342962 203068
rect 344922 203056 344928 203068
rect 344980 203096 344986 203108
rect 354582 203096 354588 203108
rect 344980 203068 354588 203096
rect 344980 203056 344986 203068
rect 354582 203056 354588 203068
rect 354640 203056 354646 203108
rect 450998 203056 451004 203108
rect 451056 203096 451062 203108
rect 513374 203096 513380 203108
rect 451056 203068 513380 203096
rect 451056 203056 451062 203068
rect 513374 203056 513380 203068
rect 513432 203056 513438 203108
rect 296622 202988 296628 203040
rect 296680 203028 296686 203040
rect 357434 203028 357440 203040
rect 296680 203000 357440 203028
rect 296680 202988 296686 203000
rect 357434 202988 357440 203000
rect 357492 202988 357498 203040
rect 453942 202988 453948 203040
rect 454000 203028 454006 203040
rect 509234 203028 509240 203040
rect 454000 203000 509240 203028
rect 454000 202988 454006 203000
rect 509234 202988 509240 203000
rect 509292 202988 509298 203040
rect 336642 202920 336648 202972
rect 336700 202960 336706 202972
rect 342898 202960 342904 202972
rect 336700 202932 342904 202960
rect 336700 202920 336706 202932
rect 342898 202920 342904 202932
rect 342956 202920 342962 202972
rect 342990 202920 342996 202972
rect 343048 202960 343054 202972
rect 353294 202960 353300 202972
rect 343048 202932 353300 202960
rect 343048 202920 343054 202932
rect 353294 202920 353300 202932
rect 353352 202920 353358 202972
rect 455322 202920 455328 202972
rect 455380 202960 455386 202972
rect 505094 202960 505100 202972
rect 455380 202932 505100 202960
rect 455380 202920 455386 202932
rect 505094 202920 505100 202932
rect 505152 202920 505158 202972
rect 295242 202852 295248 202904
rect 295300 202892 295306 202904
rect 358814 202892 358820 202904
rect 295300 202864 358820 202892
rect 295300 202852 295306 202864
rect 358814 202852 358820 202864
rect 358872 202852 358878 202904
rect 454678 202852 454684 202904
rect 454736 202892 454742 202904
rect 463050 202892 463056 202904
rect 454736 202864 463056 202892
rect 454736 202852 454742 202864
rect 463050 202852 463056 202864
rect 463108 202852 463114 202904
rect 469490 202852 469496 202904
rect 469548 202892 469554 202904
rect 477494 202892 477500 202904
rect 469548 202864 477500 202892
rect 469548 202852 469554 202864
rect 477494 202852 477500 202864
rect 477552 202852 477558 202904
rect 297358 202784 297364 202836
rect 297416 202824 297422 202836
rect 297910 202824 297916 202836
rect 297416 202796 297916 202824
rect 297416 202784 297422 202796
rect 297910 202784 297916 202796
rect 297968 202784 297974 202836
rect 408494 201560 408500 201612
rect 408552 201600 408558 201612
rect 409138 201600 409144 201612
rect 408552 201572 409144 201600
rect 408552 201560 408558 201572
rect 409138 201560 409144 201572
rect 409196 201600 409202 201612
rect 500310 201600 500316 201612
rect 409196 201572 500316 201600
rect 409196 201560 409202 201572
rect 500310 201560 500316 201572
rect 500368 201560 500374 201612
rect 297910 201492 297916 201544
rect 297968 201532 297974 201544
rect 417418 201532 417424 201544
rect 297968 201504 417424 201532
rect 297968 201492 297974 201504
rect 417418 201492 417424 201504
rect 417476 201492 417482 201544
rect 451918 201424 451924 201476
rect 451976 201464 451982 201476
rect 499666 201464 499672 201476
rect 451976 201436 499672 201464
rect 451976 201424 451982 201436
rect 499666 201424 499672 201436
rect 499724 201424 499730 201476
rect 387702 201356 387708 201408
rect 387760 201396 387766 201408
rect 500218 201396 500224 201408
rect 387760 201368 500224 201396
rect 387760 201356 387766 201368
rect 500218 201356 500224 201368
rect 500276 201356 500282 201408
rect 384942 201288 384948 201340
rect 385000 201328 385006 201340
rect 499850 201328 499856 201340
rect 385000 201300 499856 201328
rect 385000 201288 385006 201300
rect 499850 201288 499856 201300
rect 499908 201288 499914 201340
rect 383562 201220 383568 201272
rect 383620 201260 383626 201272
rect 499758 201260 499764 201272
rect 383620 201232 499764 201260
rect 383620 201220 383626 201232
rect 499758 201220 499764 201232
rect 499816 201220 499822 201272
rect 380802 201152 380808 201204
rect 380860 201192 380866 201204
rect 499942 201192 499948 201204
rect 380860 201164 499948 201192
rect 380860 201152 380866 201164
rect 499942 201152 499948 201164
rect 500000 201152 500006 201204
rect 378042 201084 378048 201136
rect 378100 201124 378106 201136
rect 500034 201124 500040 201136
rect 378100 201096 500040 201124
rect 378100 201084 378106 201096
rect 500034 201084 500040 201096
rect 500092 201084 500098 201136
rect 376662 201016 376668 201068
rect 376720 201056 376726 201068
rect 500126 201056 500132 201068
rect 376720 201028 500132 201056
rect 376720 201016 376726 201028
rect 500126 201016 500132 201028
rect 500184 201016 500190 201068
rect 2958 200948 2964 201000
rect 3016 200988 3022 201000
rect 521838 200988 521844 201000
rect 3016 200960 521844 200988
rect 3016 200948 3022 200960
rect 521838 200948 521844 200960
rect 521896 200948 521902 201000
rect 3786 200880 3792 200932
rect 3844 200920 3850 200932
rect 521746 200920 521752 200932
rect 3844 200892 521752 200920
rect 3844 200880 3850 200892
rect 521746 200880 521752 200892
rect 521804 200880 521810 200932
rect 3602 200812 3608 200864
rect 3660 200852 3666 200864
rect 521654 200852 521660 200864
rect 3660 200824 521660 200852
rect 3660 200812 3666 200824
rect 521654 200812 521660 200824
rect 521712 200812 521718 200864
rect 3878 200744 3884 200796
rect 3936 200784 3942 200796
rect 521930 200784 521936 200796
rect 3936 200756 521936 200784
rect 3936 200744 3942 200756
rect 521930 200744 521936 200756
rect 521988 200744 521994 200796
rect 379790 183472 379796 183524
rect 379848 183512 379854 183524
rect 409138 183512 409144 183524
rect 379848 183484 409144 183512
rect 379848 183472 379854 183484
rect 409138 183472 409144 183484
rect 409196 183472 409202 183524
rect 523862 182112 523868 182164
rect 523920 182152 523926 182164
rect 580166 182152 580172 182164
rect 523920 182124 580172 182152
rect 523920 182112 523926 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 522758 171028 522764 171080
rect 522816 171068 522822 171080
rect 580166 171068 580172 171080
rect 522816 171040 580172 171068
rect 522816 171028 522822 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 523770 158652 523776 158704
rect 523828 158692 523834 158704
rect 579798 158692 579804 158704
rect 523828 158664 579804 158692
rect 523828 158652 523834 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 522666 135192 522672 135244
rect 522724 135232 522730 135244
rect 580166 135232 580172 135244
rect 522724 135204 580172 135232
rect 522724 135192 522730 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 379974 124108 379980 124160
rect 380032 124148 380038 124160
rect 391198 124148 391204 124160
rect 380032 124120 391204 124148
rect 380032 124108 380038 124120
rect 391198 124108 391204 124120
rect 391256 124108 391262 124160
rect 522574 124108 522580 124160
rect 522632 124148 522638 124160
rect 580166 124148 580172 124160
rect 522632 124120 580172 124148
rect 522632 124108 522638 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 380066 118600 380072 118652
rect 380124 118640 380130 118652
rect 393958 118640 393964 118652
rect 380124 118612 393964 118640
rect 380124 118600 380130 118612
rect 393958 118600 393964 118612
rect 394016 118600 394022 118652
rect 379974 115880 379980 115932
rect 380032 115920 380038 115932
rect 395338 115920 395344 115932
rect 380032 115892 395344 115920
rect 380032 115880 380038 115892
rect 395338 115880 395344 115892
rect 395396 115880 395402 115932
rect 523678 111732 523684 111784
rect 523736 111772 523742 111784
rect 579798 111772 579804 111784
rect 523736 111744 579804 111772
rect 523736 111732 523742 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 300762 110916 300768 110968
rect 300820 110956 300826 110968
rect 416774 110956 416780 110968
rect 300820 110928 416780 110956
rect 300820 110916 300826 110928
rect 416774 110916 416780 110928
rect 416832 110916 416838 110968
rect 297910 108944 297916 108996
rect 297968 108984 297974 108996
rect 303614 108984 303620 108996
rect 297968 108956 303620 108984
rect 297968 108944 297974 108956
rect 303614 108944 303620 108956
rect 303672 108984 303678 108996
rect 305638 108984 305644 108996
rect 303672 108956 305644 108984
rect 303672 108944 303678 108956
rect 305638 108944 305644 108956
rect 305696 108984 305702 108996
rect 307754 108984 307760 108996
rect 305696 108956 307760 108984
rect 305696 108944 305702 108956
rect 307754 108944 307760 108956
rect 307812 108944 307818 108996
rect 418062 108944 418068 108996
rect 418120 108984 418126 108996
rect 424226 108984 424232 108996
rect 418120 108956 424232 108984
rect 418120 108944 418126 108956
rect 424226 108944 424232 108956
rect 424284 108984 424290 108996
rect 427814 108984 427820 108996
rect 424284 108956 427820 108984
rect 424284 108944 424290 108956
rect 427814 108944 427820 108956
rect 427872 108944 427878 108996
rect 531958 88272 531964 88324
rect 532016 88312 532022 88324
rect 580166 88312 580172 88324
rect 532016 88284 580172 88312
rect 532016 88272 532022 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 522482 77188 522488 77240
rect 522540 77228 522546 77240
rect 580166 77228 580172 77240
rect 522540 77200 580172 77228
rect 522540 77188 522546 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 527818 64812 527824 64864
rect 527876 64852 527882 64864
rect 579798 64852 579804 64864
rect 527876 64824 579804 64852
rect 527876 64812 527882 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 529198 41352 529204 41404
rect 529256 41392 529262 41404
rect 580166 41392 580172 41404
rect 529256 41364 580172 41392
rect 529256 41352 529262 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 522298 30268 522304 30320
rect 522356 30308 522362 30320
rect 580166 30308 580172 30320
rect 522356 30280 580172 30308
rect 522356 30268 522362 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 525058 17892 525064 17944
rect 525116 17932 525122 17944
rect 579798 17932 579804 17944
rect 525116 17904 579804 17932
rect 525116 17892 525122 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 522114 8276 522120 8288
rect 3476 8248 522120 8276
rect 3476 8236 3482 8248
rect 522114 8236 522120 8248
rect 522172 8236 522178 8288
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 8202 3584 8208 3596
rect 7708 3556 8208 3584
rect 7708 3544 7714 3556
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 9582 3584 9588 3596
rect 8904 3556 9588 3584
rect 8904 3544 8910 3556
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 10962 3584 10968 3596
rect 10100 3556 10968 3584
rect 10100 3544 10106 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 12342 3584 12348 3596
rect 11296 3556 12348 3584
rect 11296 3544 11302 3556
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 13630 3584 13636 3596
rect 12492 3556 13636 3584
rect 12492 3544 12498 3556
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 16482 3584 16488 3596
rect 16080 3556 16488 3584
rect 16080 3544 16086 3556
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17862 3584 17868 3596
rect 17276 3556 17868 3584
rect 17276 3544 17282 3556
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 19242 3584 19248 3596
rect 18380 3556 19248 3584
rect 18380 3544 18386 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 20622 3584 20628 3596
rect 19576 3556 20628 3584
rect 19576 3544 19582 3556
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 21910 3584 21916 3596
rect 20772 3556 21916 3584
rect 20772 3544 20778 3556
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 24762 3584 24768 3596
rect 24360 3556 24768 3584
rect 24360 3544 24366 3556
rect 24762 3544 24768 3556
rect 24820 3544 24826 3596
rect 25498 3544 25504 3596
rect 25556 3584 25562 3596
rect 26142 3584 26148 3596
rect 25556 3556 26148 3584
rect 25556 3544 25562 3556
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 26694 3544 26700 3596
rect 26752 3584 26758 3596
rect 27522 3584 27528 3596
rect 26752 3556 27528 3584
rect 26752 3544 26758 3556
rect 27522 3544 27528 3556
rect 27580 3544 27586 3596
rect 27890 3544 27896 3596
rect 27948 3584 27954 3596
rect 28902 3584 28908 3596
rect 27948 3556 28908 3584
rect 27948 3544 27954 3556
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 29086 3544 29092 3596
rect 29144 3584 29150 3596
rect 30190 3584 30196 3596
rect 29144 3556 30196 3584
rect 29144 3544 29150 3556
rect 30190 3544 30196 3556
rect 30248 3544 30254 3596
rect 33870 3544 33876 3596
rect 33928 3584 33934 3596
rect 34422 3584 34428 3596
rect 33928 3556 34428 3584
rect 33928 3544 33934 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 34974 3544 34980 3596
rect 35032 3584 35038 3596
rect 35802 3584 35808 3596
rect 35032 3556 35808 3584
rect 35032 3544 35038 3556
rect 35802 3544 35808 3556
rect 35860 3544 35866 3596
rect 36170 3544 36176 3596
rect 36228 3584 36234 3596
rect 37182 3584 37188 3596
rect 36228 3556 37188 3584
rect 36228 3544 36234 3556
rect 37182 3544 37188 3556
rect 37240 3544 37246 3596
rect 37366 3544 37372 3596
rect 37424 3584 37430 3596
rect 38470 3584 38476 3596
rect 37424 3556 38476 3584
rect 37424 3544 37430 3556
rect 38470 3544 38476 3556
rect 38528 3544 38534 3596
rect 42150 3544 42156 3596
rect 42208 3584 42214 3596
rect 42702 3584 42708 3596
rect 42208 3556 42708 3584
rect 42208 3544 42214 3556
rect 42702 3544 42708 3556
rect 42760 3544 42766 3596
rect 43346 3544 43352 3596
rect 43404 3584 43410 3596
rect 44082 3584 44088 3596
rect 43404 3556 44088 3584
rect 43404 3544 43410 3556
rect 44082 3544 44088 3556
rect 44140 3544 44146 3596
rect 44542 3544 44548 3596
rect 44600 3584 44606 3596
rect 45462 3584 45468 3596
rect 44600 3556 45468 3584
rect 44600 3544 44606 3556
rect 45462 3544 45468 3556
rect 45520 3544 45526 3596
rect 45738 3544 45744 3596
rect 45796 3584 45802 3596
rect 46842 3584 46848 3596
rect 45796 3556 46848 3584
rect 45796 3544 45802 3556
rect 46842 3544 46848 3556
rect 46900 3544 46906 3596
rect 46934 3544 46940 3596
rect 46992 3584 46998 3596
rect 48130 3584 48136 3596
rect 46992 3556 48136 3584
rect 46992 3544 46998 3556
rect 48130 3544 48136 3556
rect 48188 3544 48194 3596
rect 50522 3544 50528 3596
rect 50580 3584 50586 3596
rect 50982 3584 50988 3596
rect 50580 3556 50988 3584
rect 50580 3544 50586 3556
rect 50982 3544 50988 3556
rect 51040 3544 51046 3596
rect 51626 3544 51632 3596
rect 51684 3584 51690 3596
rect 52362 3584 52368 3596
rect 51684 3556 52368 3584
rect 51684 3544 51690 3556
rect 52362 3544 52368 3556
rect 52420 3544 52426 3596
rect 52822 3544 52828 3596
rect 52880 3584 52886 3596
rect 53742 3584 53748 3596
rect 52880 3556 53748 3584
rect 52880 3544 52886 3556
rect 53742 3544 53748 3556
rect 53800 3544 53806 3596
rect 54018 3544 54024 3596
rect 54076 3584 54082 3596
rect 55122 3584 55128 3596
rect 54076 3556 55128 3584
rect 54076 3544 54082 3556
rect 55122 3544 55128 3556
rect 55180 3544 55186 3596
rect 55214 3544 55220 3596
rect 55272 3584 55278 3596
rect 56410 3584 56416 3596
rect 55272 3556 56416 3584
rect 55272 3544 55278 3556
rect 56410 3544 56416 3556
rect 56468 3544 56474 3596
rect 58802 3544 58808 3596
rect 58860 3584 58866 3596
rect 59262 3584 59268 3596
rect 58860 3556 59268 3584
rect 58860 3544 58866 3556
rect 59262 3544 59268 3556
rect 59320 3544 59326 3596
rect 59998 3544 60004 3596
rect 60056 3584 60062 3596
rect 60642 3584 60648 3596
rect 60056 3556 60648 3584
rect 60056 3544 60062 3556
rect 60642 3544 60648 3556
rect 60700 3544 60706 3596
rect 61194 3544 61200 3596
rect 61252 3584 61258 3596
rect 62022 3584 62028 3596
rect 61252 3556 62028 3584
rect 61252 3544 61258 3556
rect 62022 3544 62028 3556
rect 62080 3544 62086 3596
rect 63586 3544 63592 3596
rect 63644 3584 63650 3596
rect 64690 3584 64696 3596
rect 63644 3556 64696 3584
rect 63644 3544 63650 3556
rect 64690 3544 64696 3556
rect 64748 3544 64754 3596
rect 68278 3544 68284 3596
rect 68336 3584 68342 3596
rect 68922 3584 68928 3596
rect 68336 3556 68928 3584
rect 68336 3544 68342 3556
rect 68922 3544 68928 3556
rect 68980 3544 68986 3596
rect 69474 3544 69480 3596
rect 69532 3584 69538 3596
rect 70302 3584 70308 3596
rect 69532 3556 70308 3584
rect 69532 3544 69538 3556
rect 70302 3544 70308 3556
rect 70360 3544 70366 3596
rect 70670 3544 70676 3596
rect 70728 3584 70734 3596
rect 71682 3584 71688 3596
rect 70728 3556 71688 3584
rect 70728 3544 70734 3556
rect 71682 3544 71688 3556
rect 71740 3544 71746 3596
rect 71866 3544 71872 3596
rect 71924 3584 71930 3596
rect 72970 3584 72976 3596
rect 71924 3556 72976 3584
rect 71924 3544 71930 3556
rect 72970 3544 72976 3556
rect 73028 3544 73034 3596
rect 76650 3544 76656 3596
rect 76708 3584 76714 3596
rect 77202 3584 77208 3596
rect 76708 3556 77208 3584
rect 76708 3544 76714 3556
rect 77202 3544 77208 3556
rect 77260 3544 77266 3596
rect 77846 3544 77852 3596
rect 77904 3584 77910 3596
rect 78582 3584 78588 3596
rect 77904 3556 78588 3584
rect 77904 3544 77910 3556
rect 78582 3544 78588 3556
rect 78640 3544 78646 3596
rect 79042 3544 79048 3596
rect 79100 3584 79106 3596
rect 79962 3584 79968 3596
rect 79100 3556 79968 3584
rect 79100 3544 79106 3556
rect 79962 3544 79968 3556
rect 80020 3544 80026 3596
rect 80238 3544 80244 3596
rect 80296 3584 80302 3596
rect 81342 3584 81348 3596
rect 80296 3556 81348 3584
rect 80296 3544 80302 3556
rect 81342 3544 81348 3556
rect 81400 3544 81406 3596
rect 81434 3544 81440 3596
rect 81492 3584 81498 3596
rect 82630 3584 82636 3596
rect 81492 3556 82636 3584
rect 81492 3544 81498 3556
rect 82630 3544 82636 3556
rect 82688 3544 82694 3596
rect 84930 3544 84936 3596
rect 84988 3584 84994 3596
rect 85482 3584 85488 3596
rect 84988 3556 85488 3584
rect 84988 3544 84994 3556
rect 85482 3544 85488 3556
rect 85540 3544 85546 3596
rect 86126 3544 86132 3596
rect 86184 3584 86190 3596
rect 86862 3584 86868 3596
rect 86184 3556 86868 3584
rect 86184 3544 86190 3556
rect 86862 3544 86868 3556
rect 86920 3544 86926 3596
rect 87322 3544 87328 3596
rect 87380 3584 87386 3596
rect 88242 3584 88248 3596
rect 87380 3556 88248 3584
rect 87380 3544 87386 3556
rect 88242 3544 88248 3556
rect 88300 3544 88306 3596
rect 88518 3544 88524 3596
rect 88576 3584 88582 3596
rect 89622 3584 89628 3596
rect 88576 3556 89628 3584
rect 88576 3544 88582 3556
rect 89622 3544 89628 3556
rect 89680 3544 89686 3596
rect 89714 3544 89720 3596
rect 89772 3584 89778 3596
rect 90910 3584 90916 3596
rect 89772 3556 90916 3584
rect 89772 3544 89778 3556
rect 90910 3544 90916 3556
rect 90968 3544 90974 3596
rect 93302 3544 93308 3596
rect 93360 3584 93366 3596
rect 93762 3584 93768 3596
rect 93360 3556 93768 3584
rect 93360 3544 93366 3556
rect 93762 3544 93768 3556
rect 93820 3544 93826 3596
rect 94498 3544 94504 3596
rect 94556 3584 94562 3596
rect 95142 3584 95148 3596
rect 94556 3556 95148 3584
rect 94556 3544 94562 3556
rect 95142 3544 95148 3556
rect 95200 3544 95206 3596
rect 95694 3544 95700 3596
rect 95752 3584 95758 3596
rect 96522 3584 96528 3596
rect 95752 3556 96528 3584
rect 95752 3544 95758 3556
rect 96522 3544 96528 3556
rect 96580 3544 96586 3596
rect 96890 3544 96896 3596
rect 96948 3584 96954 3596
rect 97902 3584 97908 3596
rect 96948 3556 97908 3584
rect 96948 3544 96954 3556
rect 97902 3544 97908 3556
rect 97960 3544 97966 3596
rect 98086 3544 98092 3596
rect 98144 3584 98150 3596
rect 99190 3584 99196 3596
rect 98144 3556 99196 3584
rect 98144 3544 98150 3556
rect 99190 3544 99196 3556
rect 99248 3544 99254 3596
rect 102778 3544 102784 3596
rect 102836 3584 102842 3596
rect 103422 3584 103428 3596
rect 102836 3556 103428 3584
rect 102836 3544 102842 3556
rect 103422 3544 103428 3556
rect 103480 3544 103486 3596
rect 103974 3544 103980 3596
rect 104032 3584 104038 3596
rect 104802 3584 104808 3596
rect 104032 3556 104808 3584
rect 104032 3544 104038 3556
rect 104802 3544 104808 3556
rect 104860 3544 104866 3596
rect 105170 3544 105176 3596
rect 105228 3584 105234 3596
rect 106182 3584 106188 3596
rect 105228 3556 106188 3584
rect 105228 3544 105234 3556
rect 106182 3544 106188 3556
rect 106240 3544 106246 3596
rect 106366 3544 106372 3596
rect 106424 3584 106430 3596
rect 107470 3584 107476 3596
rect 106424 3556 107476 3584
rect 106424 3544 106430 3556
rect 107470 3544 107476 3556
rect 107528 3544 107534 3596
rect 111150 3544 111156 3596
rect 111208 3584 111214 3596
rect 111702 3584 111708 3596
rect 111208 3556 111708 3584
rect 111208 3544 111214 3556
rect 111702 3544 111708 3556
rect 111760 3544 111766 3596
rect 112346 3544 112352 3596
rect 112404 3584 112410 3596
rect 113082 3584 113088 3596
rect 112404 3556 113088 3584
rect 112404 3544 112410 3556
rect 113082 3544 113088 3556
rect 113140 3544 113146 3596
rect 113542 3544 113548 3596
rect 113600 3584 113606 3596
rect 114462 3584 114468 3596
rect 113600 3556 114468 3584
rect 113600 3544 113606 3556
rect 114462 3544 114468 3556
rect 114520 3544 114526 3596
rect 114738 3544 114744 3596
rect 114796 3584 114802 3596
rect 115842 3584 115848 3596
rect 114796 3556 115848 3584
rect 114796 3544 114802 3556
rect 115842 3544 115848 3556
rect 115900 3544 115906 3596
rect 115934 3544 115940 3596
rect 115992 3584 115998 3596
rect 117130 3584 117136 3596
rect 115992 3556 117136 3584
rect 115992 3544 115998 3556
rect 117130 3544 117136 3556
rect 117188 3544 117194 3596
rect 119430 3544 119436 3596
rect 119488 3584 119494 3596
rect 119982 3584 119988 3596
rect 119488 3556 119988 3584
rect 119488 3544 119494 3556
rect 119982 3544 119988 3556
rect 120040 3544 120046 3596
rect 120626 3544 120632 3596
rect 120684 3584 120690 3596
rect 121362 3584 121368 3596
rect 120684 3556 121368 3584
rect 120684 3544 120690 3556
rect 121362 3544 121368 3556
rect 121420 3544 121426 3596
rect 121822 3544 121828 3596
rect 121880 3584 121886 3596
rect 122742 3584 122748 3596
rect 121880 3556 122748 3584
rect 121880 3544 121886 3556
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 123018 3544 123024 3596
rect 123076 3584 123082 3596
rect 124122 3584 124128 3596
rect 123076 3556 124128 3584
rect 123076 3544 123082 3556
rect 124122 3544 124128 3556
rect 124180 3544 124186 3596
rect 124214 3544 124220 3596
rect 124272 3584 124278 3596
rect 125410 3584 125416 3596
rect 124272 3556 125416 3584
rect 124272 3544 124278 3556
rect 125410 3544 125416 3556
rect 125468 3544 125474 3596
rect 127802 3544 127808 3596
rect 127860 3584 127866 3596
rect 128262 3584 128268 3596
rect 127860 3556 128268 3584
rect 127860 3544 127866 3556
rect 128262 3544 128268 3556
rect 128320 3544 128326 3596
rect 128998 3544 129004 3596
rect 129056 3584 129062 3596
rect 129642 3584 129648 3596
rect 129056 3556 129648 3584
rect 129056 3544 129062 3556
rect 129642 3544 129648 3556
rect 129700 3544 129706 3596
rect 130194 3544 130200 3596
rect 130252 3584 130258 3596
rect 131022 3584 131028 3596
rect 130252 3556 131028 3584
rect 130252 3544 130258 3556
rect 131022 3544 131028 3556
rect 131080 3544 131086 3596
rect 131390 3544 131396 3596
rect 131448 3584 131454 3596
rect 132402 3584 132408 3596
rect 131448 3556 132408 3584
rect 131448 3544 131454 3556
rect 132402 3544 132408 3556
rect 132460 3544 132466 3596
rect 132586 3544 132592 3596
rect 132644 3584 132650 3596
rect 133782 3584 133788 3596
rect 132644 3556 133788 3584
rect 132644 3544 132650 3556
rect 133782 3544 133788 3556
rect 133840 3544 133846 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 278130 3516 278136 3528
rect 2924 3488 278136 3516
rect 2924 3476 2930 3488
rect 278130 3476 278136 3488
rect 278188 3476 278194 3528
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 278038 3448 278044 3460
rect 4120 3420 278044 3448
rect 4120 3408 4126 3420
rect 278038 3408 278044 3420
rect 278096 3408 278102 3460
rect 101582 3272 101588 3324
rect 101640 3312 101646 3324
rect 102042 3312 102048 3324
rect 101640 3284 102048 3312
rect 101640 3272 101646 3284
rect 102042 3272 102048 3284
rect 102100 3272 102106 3324
rect 62390 3136 62396 3188
rect 62448 3176 62454 3188
rect 63402 3176 63408 3188
rect 62448 3148 63408 3176
rect 62448 3136 62454 3148
rect 63402 3136 63408 3148
rect 63460 3136 63466 3188
rect 142062 2796 142068 2848
rect 142120 2836 142126 2848
rect 145650 2836 145656 2848
rect 142120 2808 145656 2836
rect 142120 2796 142126 2808
rect 145650 2796 145656 2808
rect 145708 2836 145714 2848
rect 149238 2836 149244 2848
rect 145708 2808 149244 2836
rect 145708 2796 145714 2808
rect 149238 2796 149244 2808
rect 149296 2836 149302 2848
rect 152734 2836 152740 2848
rect 149296 2808 152740 2836
rect 149296 2796 149302 2808
rect 152734 2796 152740 2808
rect 152792 2836 152798 2848
rect 156322 2836 156328 2848
rect 152792 2808 156328 2836
rect 152792 2796 152798 2808
rect 156322 2796 156328 2808
rect 156380 2836 156386 2848
rect 159910 2836 159916 2848
rect 156380 2808 159916 2836
rect 156380 2796 156386 2808
rect 159910 2796 159916 2808
rect 159968 2836 159974 2848
rect 163498 2836 163504 2848
rect 159968 2808 163504 2836
rect 159968 2796 159974 2808
rect 163498 2796 163504 2808
rect 163556 2836 163562 2848
rect 167086 2836 167092 2848
rect 163556 2808 167092 2836
rect 163556 2796 163562 2808
rect 167086 2796 167092 2808
rect 167144 2836 167150 2848
rect 170582 2836 170588 2848
rect 167144 2808 170588 2836
rect 167144 2796 167150 2808
rect 170582 2796 170588 2808
rect 170640 2836 170646 2848
rect 174170 2836 174176 2848
rect 170640 2808 174176 2836
rect 170640 2796 170646 2808
rect 174170 2796 174176 2808
rect 174228 2836 174234 2848
rect 177758 2836 177764 2848
rect 174228 2808 177764 2836
rect 174228 2796 174234 2808
rect 177758 2796 177764 2808
rect 177816 2836 177822 2848
rect 181346 2836 181352 2848
rect 177816 2808 181352 2836
rect 177816 2796 177822 2808
rect 181346 2796 181352 2808
rect 181404 2836 181410 2848
rect 184842 2836 184848 2848
rect 181404 2808 184848 2836
rect 181404 2796 181410 2808
rect 184842 2796 184848 2808
rect 184900 2836 184906 2848
rect 188430 2836 188436 2848
rect 184900 2808 188436 2836
rect 184900 2796 184906 2808
rect 188430 2796 188436 2808
rect 188488 2836 188494 2848
rect 192018 2836 192024 2848
rect 188488 2808 192024 2836
rect 188488 2796 188494 2808
rect 192018 2796 192024 2808
rect 192076 2836 192082 2848
rect 195606 2836 195612 2848
rect 192076 2808 195612 2836
rect 192076 2796 192082 2808
rect 195606 2796 195612 2808
rect 195664 2836 195670 2848
rect 199194 2836 199200 2848
rect 195664 2808 199200 2836
rect 195664 2796 195670 2808
rect 199194 2796 199200 2808
rect 199252 2836 199258 2848
rect 202690 2836 202696 2848
rect 199252 2808 202696 2836
rect 199252 2796 199258 2808
rect 202690 2796 202696 2808
rect 202748 2836 202754 2848
rect 206278 2836 206284 2848
rect 202748 2808 206284 2836
rect 202748 2796 202754 2808
rect 206278 2796 206284 2808
rect 206336 2836 206342 2848
rect 209866 2836 209872 2848
rect 206336 2808 209872 2836
rect 206336 2796 206342 2808
rect 209866 2796 209872 2808
rect 209924 2836 209930 2848
rect 213454 2836 213460 2848
rect 209924 2808 213460 2836
rect 209924 2796 209930 2808
rect 213454 2796 213460 2808
rect 213512 2836 213518 2848
rect 217042 2836 217048 2848
rect 213512 2808 217048 2836
rect 213512 2796 213518 2808
rect 217042 2796 217048 2808
rect 217100 2836 217106 2848
rect 220538 2836 220544 2848
rect 217100 2808 220544 2836
rect 217100 2796 217106 2808
rect 220538 2796 220544 2808
rect 220596 2836 220602 2848
rect 224126 2836 224132 2848
rect 220596 2808 224132 2836
rect 220596 2796 220602 2808
rect 224126 2796 224132 2808
rect 224184 2836 224190 2848
rect 227714 2836 227720 2848
rect 224184 2808 227720 2836
rect 224184 2796 224190 2808
rect 227714 2796 227720 2808
rect 227772 2836 227778 2848
rect 231302 2836 231308 2848
rect 227772 2808 231308 2836
rect 227772 2796 227778 2808
rect 231302 2796 231308 2808
rect 231360 2836 231366 2848
rect 234798 2836 234804 2848
rect 231360 2808 234804 2836
rect 231360 2796 231366 2808
rect 234798 2796 234804 2808
rect 234856 2836 234862 2848
rect 238386 2836 238392 2848
rect 234856 2808 238392 2836
rect 234856 2796 234862 2808
rect 238386 2796 238392 2808
rect 238444 2836 238450 2848
rect 241974 2836 241980 2848
rect 238444 2808 241980 2836
rect 238444 2796 238450 2808
rect 241974 2796 241980 2808
rect 242032 2836 242038 2848
rect 245562 2836 245568 2848
rect 242032 2808 245568 2836
rect 242032 2796 242038 2808
rect 245562 2796 245568 2808
rect 245620 2836 245626 2848
rect 249150 2836 249156 2848
rect 245620 2808 249156 2836
rect 245620 2796 245626 2808
rect 249150 2796 249156 2808
rect 249208 2836 249214 2848
rect 252646 2836 252652 2848
rect 249208 2808 252652 2836
rect 249208 2796 249214 2808
rect 252646 2796 252652 2808
rect 252704 2836 252710 2848
rect 256234 2836 256240 2848
rect 252704 2808 256240 2836
rect 252704 2796 252710 2808
rect 256234 2796 256240 2808
rect 256292 2836 256298 2848
rect 259822 2836 259828 2848
rect 256292 2808 259828 2836
rect 256292 2796 256298 2808
rect 259822 2796 259828 2808
rect 259880 2836 259886 2848
rect 263410 2836 263416 2848
rect 259880 2808 263416 2836
rect 259880 2796 259886 2808
rect 263410 2796 263416 2808
rect 263468 2836 263474 2848
rect 266998 2836 267004 2848
rect 263468 2808 267004 2836
rect 263468 2796 263474 2808
rect 266998 2796 267004 2808
rect 267056 2836 267062 2848
rect 270494 2836 270500 2848
rect 267056 2808 270500 2836
rect 267056 2796 267062 2808
rect 270494 2796 270500 2808
rect 270552 2836 270558 2848
rect 274082 2836 274088 2848
rect 270552 2808 274088 2836
rect 270552 2796 270558 2808
rect 274082 2796 274088 2808
rect 274140 2836 274146 2848
rect 277670 2836 277676 2848
rect 274140 2808 277676 2836
rect 274140 2796 274146 2808
rect 277670 2796 277676 2808
rect 277728 2836 277734 2848
rect 281258 2836 281264 2848
rect 277728 2808 281264 2836
rect 277728 2796 277734 2808
rect 281258 2796 281264 2808
rect 281316 2836 281322 2848
rect 284754 2836 284760 2848
rect 281316 2808 284760 2836
rect 281316 2796 281322 2808
rect 284754 2796 284760 2808
rect 284812 2836 284818 2848
rect 288342 2836 288348 2848
rect 284812 2808 288348 2836
rect 284812 2796 284818 2808
rect 288342 2796 288348 2808
rect 288400 2836 288406 2848
rect 291930 2836 291936 2848
rect 288400 2808 291936 2836
rect 288400 2796 288406 2808
rect 291930 2796 291936 2808
rect 291988 2836 291994 2848
rect 295518 2836 295524 2848
rect 291988 2808 295524 2836
rect 291988 2796 291994 2808
rect 295518 2796 295524 2808
rect 295576 2836 295582 2848
rect 299106 2836 299112 2848
rect 295576 2808 299112 2836
rect 295576 2796 295582 2808
rect 299106 2796 299112 2808
rect 299164 2836 299170 2848
rect 302602 2836 302608 2848
rect 299164 2808 302608 2836
rect 299164 2796 299170 2808
rect 302602 2796 302608 2808
rect 302660 2836 302666 2848
rect 305638 2836 305644 2848
rect 302660 2808 305644 2836
rect 302660 2796 302666 2808
rect 305638 2796 305644 2808
rect 305696 2836 305702 2848
rect 306190 2836 306196 2848
rect 305696 2808 306196 2836
rect 305696 2796 305702 2808
rect 306190 2796 306196 2808
rect 306248 2836 306254 2848
rect 309778 2836 309784 2848
rect 306248 2808 309784 2836
rect 306248 2796 306254 2808
rect 309778 2796 309784 2808
rect 309836 2836 309842 2848
rect 313366 2836 313372 2848
rect 309836 2808 313372 2836
rect 309836 2796 309842 2808
rect 313366 2796 313372 2808
rect 313424 2836 313430 2848
rect 316954 2836 316960 2848
rect 313424 2808 316960 2836
rect 313424 2796 313430 2808
rect 316954 2796 316960 2808
rect 317012 2836 317018 2848
rect 320450 2836 320456 2848
rect 317012 2808 320456 2836
rect 317012 2796 317018 2808
rect 320450 2796 320456 2808
rect 320508 2836 320514 2848
rect 324038 2836 324044 2848
rect 320508 2808 324044 2836
rect 320508 2796 320514 2808
rect 324038 2796 324044 2808
rect 324096 2836 324102 2848
rect 327626 2836 327632 2848
rect 324096 2808 327632 2836
rect 324096 2796 324102 2808
rect 327626 2796 327632 2808
rect 327684 2836 327690 2848
rect 331214 2836 331220 2848
rect 327684 2808 331220 2836
rect 327684 2796 327690 2808
rect 331214 2796 331220 2808
rect 331272 2836 331278 2848
rect 334710 2836 334716 2848
rect 331272 2808 334716 2836
rect 331272 2796 331278 2808
rect 334710 2796 334716 2808
rect 334768 2836 334774 2848
rect 338298 2836 338304 2848
rect 334768 2808 338304 2836
rect 334768 2796 334774 2808
rect 338298 2796 338304 2808
rect 338356 2836 338362 2848
rect 341886 2836 341892 2848
rect 338356 2808 341892 2836
rect 338356 2796 338362 2808
rect 341886 2796 341892 2808
rect 341944 2836 341950 2848
rect 345474 2836 345480 2848
rect 341944 2808 345480 2836
rect 341944 2796 341950 2808
rect 345474 2796 345480 2808
rect 345532 2836 345538 2848
rect 349062 2836 349068 2848
rect 345532 2808 349068 2836
rect 345532 2796 345538 2808
rect 349062 2796 349068 2808
rect 349120 2836 349126 2848
rect 352558 2836 352564 2848
rect 349120 2808 352564 2836
rect 349120 2796 349126 2808
rect 352558 2796 352564 2808
rect 352616 2836 352622 2848
rect 356146 2836 356152 2848
rect 352616 2808 356152 2836
rect 352616 2796 352622 2808
rect 356146 2796 356152 2808
rect 356204 2836 356210 2848
rect 359734 2836 359740 2848
rect 356204 2808 359740 2836
rect 356204 2796 356210 2808
rect 359734 2796 359740 2808
rect 359792 2836 359798 2848
rect 363322 2836 363328 2848
rect 359792 2808 363328 2836
rect 359792 2796 359798 2808
rect 363322 2796 363328 2808
rect 363380 2836 363386 2848
rect 366910 2836 366916 2848
rect 363380 2808 366916 2836
rect 363380 2796 363386 2808
rect 366910 2796 366916 2808
rect 366968 2836 366974 2848
rect 370406 2836 370412 2848
rect 366968 2808 370412 2836
rect 366968 2796 366974 2808
rect 370406 2796 370412 2808
rect 370464 2836 370470 2848
rect 373994 2836 374000 2848
rect 370464 2808 374000 2836
rect 370464 2796 370470 2808
rect 373994 2796 374000 2808
rect 374052 2836 374058 2848
rect 377582 2836 377588 2848
rect 374052 2808 377588 2836
rect 374052 2796 374058 2808
rect 377582 2796 377588 2808
rect 377640 2836 377646 2848
rect 381170 2836 381176 2848
rect 377640 2808 381176 2836
rect 377640 2796 377646 2808
rect 381170 2796 381176 2808
rect 381228 2836 381234 2848
rect 384666 2836 384672 2848
rect 381228 2808 384672 2836
rect 381228 2796 381234 2808
rect 384666 2796 384672 2808
rect 384724 2836 384730 2848
rect 388254 2836 388260 2848
rect 384724 2808 388260 2836
rect 384724 2796 384730 2808
rect 388254 2796 388260 2808
rect 388312 2836 388318 2848
rect 391842 2836 391848 2848
rect 388312 2808 391848 2836
rect 388312 2796 388318 2808
rect 391842 2796 391848 2808
rect 391900 2836 391906 2848
rect 395430 2836 395436 2848
rect 391900 2808 395436 2836
rect 391900 2796 391906 2808
rect 395430 2796 395436 2808
rect 395488 2836 395494 2848
rect 399018 2836 399024 2848
rect 395488 2808 399024 2836
rect 395488 2796 395494 2808
rect 399018 2796 399024 2808
rect 399076 2836 399082 2848
rect 402514 2836 402520 2848
rect 399076 2808 402520 2836
rect 399076 2796 399082 2808
rect 402514 2796 402520 2808
rect 402572 2836 402578 2848
rect 406102 2836 406108 2848
rect 402572 2808 406108 2836
rect 402572 2796 402578 2808
rect 406102 2796 406108 2808
rect 406160 2836 406166 2848
rect 409690 2836 409696 2848
rect 406160 2808 409696 2836
rect 406160 2796 406166 2808
rect 409690 2796 409696 2808
rect 409748 2836 409754 2848
rect 413278 2836 413284 2848
rect 409748 2808 413284 2836
rect 409748 2796 409754 2808
rect 413278 2796 413284 2808
rect 413336 2836 413342 2848
rect 416866 2836 416872 2848
rect 413336 2808 416872 2836
rect 413336 2796 413342 2808
rect 416866 2796 416872 2808
rect 416924 2836 416930 2848
rect 420362 2836 420368 2848
rect 416924 2808 420368 2836
rect 416924 2796 416930 2808
rect 420362 2796 420368 2808
rect 420420 2836 420426 2848
rect 423950 2836 423956 2848
rect 420420 2808 423956 2836
rect 420420 2796 420426 2808
rect 423950 2796 423956 2808
rect 424008 2836 424014 2848
rect 427538 2836 427544 2848
rect 424008 2808 427544 2836
rect 424008 2796 424014 2808
rect 427538 2796 427544 2808
rect 427596 2836 427602 2848
rect 431126 2836 431132 2848
rect 427596 2808 431132 2836
rect 427596 2796 427602 2808
rect 431126 2796 431132 2808
rect 431184 2836 431190 2848
rect 434622 2836 434628 2848
rect 431184 2808 434628 2836
rect 431184 2796 431190 2808
rect 434622 2796 434628 2808
rect 434680 2836 434686 2848
rect 438210 2836 438216 2848
rect 434680 2808 438216 2836
rect 434680 2796 434686 2808
rect 438210 2796 438216 2808
rect 438268 2836 438274 2848
rect 441798 2836 441804 2848
rect 438268 2808 441804 2836
rect 438268 2796 438274 2808
rect 441798 2796 441804 2808
rect 441856 2836 441862 2848
rect 445386 2836 445392 2848
rect 441856 2808 445392 2836
rect 441856 2796 441862 2808
rect 445386 2796 445392 2808
rect 445444 2836 445450 2848
rect 448974 2836 448980 2848
rect 445444 2808 448980 2836
rect 445444 2796 445450 2808
rect 448974 2796 448980 2808
rect 449032 2836 449038 2848
rect 452470 2836 452476 2848
rect 449032 2808 452476 2836
rect 449032 2796 449038 2808
rect 452470 2796 452476 2808
rect 452528 2836 452534 2848
rect 456058 2836 456064 2848
rect 452528 2808 456064 2836
rect 452528 2796 452534 2808
rect 456058 2796 456064 2808
rect 456116 2836 456122 2848
rect 459646 2836 459652 2848
rect 456116 2808 459652 2836
rect 456116 2796 456122 2808
rect 459646 2796 459652 2808
rect 459704 2836 459710 2848
rect 463234 2836 463240 2848
rect 459704 2808 463240 2836
rect 459704 2796 459710 2808
rect 463234 2796 463240 2808
rect 463292 2836 463298 2848
rect 466822 2836 466828 2848
rect 463292 2808 466828 2836
rect 463292 2796 463298 2808
rect 466822 2796 466828 2808
rect 466880 2836 466886 2848
rect 470318 2836 470324 2848
rect 466880 2808 470324 2836
rect 466880 2796 466886 2808
rect 470318 2796 470324 2808
rect 470376 2836 470382 2848
rect 473906 2836 473912 2848
rect 470376 2808 473912 2836
rect 470376 2796 470382 2808
rect 473906 2796 473912 2808
rect 473964 2836 473970 2848
rect 477494 2836 477500 2848
rect 473964 2808 477500 2836
rect 473964 2796 473970 2808
rect 477494 2796 477500 2808
rect 477552 2836 477558 2848
rect 481082 2836 481088 2848
rect 477552 2808 481088 2836
rect 477552 2796 477558 2808
rect 481082 2796 481088 2808
rect 481140 2836 481146 2848
rect 484578 2836 484584 2848
rect 481140 2808 484584 2836
rect 481140 2796 481146 2808
rect 484578 2796 484584 2808
rect 484636 2836 484642 2848
rect 488166 2836 488172 2848
rect 484636 2808 488172 2836
rect 484636 2796 484642 2808
rect 488166 2796 488172 2808
rect 488224 2836 488230 2848
rect 491754 2836 491760 2848
rect 488224 2808 491760 2836
rect 488224 2796 488230 2808
rect 491754 2796 491760 2808
rect 491812 2836 491818 2848
rect 495342 2836 495348 2848
rect 491812 2808 495348 2836
rect 491812 2796 491818 2808
rect 495342 2796 495348 2808
rect 495400 2836 495406 2848
rect 498930 2836 498936 2848
rect 495400 2808 498936 2836
rect 495400 2796 495406 2808
rect 498930 2796 498936 2808
rect 498988 2836 498994 2848
rect 502426 2836 502432 2848
rect 498988 2808 502432 2836
rect 498988 2796 498994 2808
rect 502426 2796 502432 2808
rect 502484 2836 502490 2848
rect 506014 2836 506020 2848
rect 502484 2808 506020 2836
rect 502484 2796 502490 2808
rect 506014 2796 506020 2808
rect 506072 2836 506078 2848
rect 509602 2836 509608 2848
rect 506072 2808 509608 2836
rect 506072 2796 506078 2808
rect 509602 2796 509608 2808
rect 509660 2836 509666 2848
rect 513190 2836 513196 2848
rect 509660 2808 513196 2836
rect 509660 2796 509666 2808
rect 513190 2796 513196 2808
rect 513248 2836 513254 2848
rect 516778 2836 516784 2848
rect 513248 2808 516784 2836
rect 513248 2796 513254 2808
rect 516778 2796 516784 2808
rect 516836 2836 516842 2848
rect 520274 2836 520280 2848
rect 516836 2808 520280 2836
rect 516836 2796 516842 2808
rect 520274 2796 520280 2808
rect 520332 2836 520338 2848
rect 523862 2836 523868 2848
rect 520332 2808 523868 2836
rect 520332 2796 520338 2808
rect 523862 2796 523868 2808
rect 523920 2836 523926 2848
rect 527450 2836 527456 2848
rect 523920 2808 527456 2836
rect 523920 2796 523926 2808
rect 527450 2796 527456 2808
rect 527508 2836 527514 2848
rect 531038 2836 531044 2848
rect 527508 2808 531044 2836
rect 527508 2796 527514 2808
rect 531038 2796 531044 2808
rect 531096 2836 531102 2848
rect 534534 2836 534540 2848
rect 531096 2808 534540 2836
rect 531096 2796 531102 2808
rect 534534 2796 534540 2808
rect 534592 2836 534598 2848
rect 538122 2836 538128 2848
rect 534592 2808 538128 2836
rect 534592 2796 534598 2808
rect 538122 2796 538128 2808
rect 538180 2836 538186 2848
rect 541710 2836 541716 2848
rect 538180 2808 541716 2836
rect 538180 2796 538186 2808
rect 541710 2796 541716 2808
rect 541768 2836 541774 2848
rect 545298 2836 545304 2848
rect 541768 2808 545304 2836
rect 541768 2796 541774 2808
rect 545298 2796 545304 2808
rect 545356 2836 545362 2848
rect 548886 2836 548892 2848
rect 545356 2808 548892 2836
rect 545356 2796 545362 2808
rect 548886 2796 548892 2808
rect 548944 2836 548950 2848
rect 552382 2836 552388 2848
rect 548944 2808 552388 2836
rect 548944 2796 548950 2808
rect 552382 2796 552388 2808
rect 552440 2836 552446 2848
rect 555970 2836 555976 2848
rect 552440 2808 555976 2836
rect 552440 2796 552446 2808
rect 555970 2796 555976 2808
rect 556028 2836 556034 2848
rect 559558 2836 559564 2848
rect 556028 2808 559564 2836
rect 556028 2796 556034 2808
rect 559558 2796 559564 2808
rect 559616 2836 559622 2848
rect 563146 2836 563152 2848
rect 559616 2808 563152 2836
rect 559616 2796 559622 2808
rect 563146 2796 563152 2808
rect 563204 2836 563210 2848
rect 566734 2836 566740 2848
rect 563204 2808 566740 2836
rect 563204 2796 563210 2808
rect 566734 2796 566740 2808
rect 566792 2836 566798 2848
rect 570230 2836 570236 2848
rect 566792 2808 570236 2836
rect 566792 2796 566798 2808
rect 570230 2796 570236 2808
rect 570288 2836 570294 2848
rect 573818 2836 573824 2848
rect 570288 2808 573824 2836
rect 570288 2796 570294 2808
rect 573818 2796 573824 2808
rect 573876 2836 573882 2848
rect 577406 2836 577412 2848
rect 573876 2808 577412 2836
rect 573876 2796 573882 2808
rect 577406 2796 577412 2808
rect 577464 2836 577470 2848
rect 580994 2836 581000 2848
rect 577464 2808 581000 2836
rect 577464 2796 577470 2808
rect 580994 2796 581000 2808
rect 581052 2796 581058 2848
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 5442 592 5448 604
rect 5316 564 5448 592
rect 5316 552 5322 564
rect 5442 552 5448 564
rect 5500 552 5506 604
rect 138474 552 138480 604
rect 138532 592 138538 604
rect 142062 592 142068 604
rect 138532 564 142068 592
rect 138532 552 138538 564
rect 142062 552 142068 564
rect 142120 552 142126 604
<< via1 >>
rect 170312 700884 170364 700936
rect 171048 700884 171100 700936
rect 478512 700816 478564 700868
rect 519084 700816 519136 700868
rect 413652 700748 413704 700800
rect 519176 700748 519228 700800
rect 348792 700680 348844 700732
rect 520280 700680 520332 700732
rect 283840 700612 283892 700664
rect 520372 700612 520424 700664
rect 267648 700544 267700 700596
rect 519268 700544 519320 700596
rect 218980 700476 219032 700528
rect 519452 700476 519504 700528
rect 202788 700408 202840 700460
rect 519360 700408 519412 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 154120 700340 154172 700392
rect 520464 700340 520516 700392
rect 137836 700272 137888 700324
rect 519544 700272 519596 700324
rect 531964 700272 532016 700324
rect 559656 700272 559708 700324
rect 462320 700068 462372 700120
rect 463608 700068 463660 700120
rect 397460 699932 397512 699984
rect 398748 699932 398800 699984
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300584 699660 300636 699712
rect 364984 699660 365036 699712
rect 365628 699660 365680 699712
rect 429844 699660 429896 699712
rect 430488 699660 430540 699712
rect 494796 699660 494848 699712
rect 495348 699660 495400 699712
rect 542728 698232 542780 698284
rect 543556 698232 543608 698284
rect 545764 696940 545816 696992
rect 580172 696940 580224 696992
rect 542544 694084 542596 694136
rect 542728 694084 542780 694136
rect 560944 685856 560996 685908
rect 580172 685856 580224 685908
rect 542452 684496 542504 684548
rect 542544 684496 542596 684548
rect 529204 673480 529256 673532
rect 580172 673480 580224 673532
rect 542544 666544 542596 666596
rect 542820 666544 542872 666596
rect 542544 661716 542596 661768
rect 542820 661716 542872 661768
rect 542544 656888 542596 656940
rect 542636 656888 542688 656940
rect 540244 650020 540296 650072
rect 580172 650020 580224 650072
rect 542544 647232 542596 647284
rect 542636 647232 542688 647284
rect 542544 640364 542596 640416
rect 542636 640364 542688 640416
rect 558184 638936 558236 638988
rect 580172 638936 580224 638988
rect 542452 630640 542504 630692
rect 542636 630640 542688 630692
rect 525064 626560 525116 626612
rect 580172 626560 580224 626612
rect 488540 613368 488592 613420
rect 493968 613368 494020 613420
rect 373632 612756 373684 612808
rect 379612 612756 379664 612808
rect 488540 612756 488592 612808
rect 493968 612756 494020 612808
rect 499580 612756 499632 612808
rect 542452 611328 542504 611380
rect 542636 611328 542688 611380
rect 495348 610852 495400 610904
rect 520556 610852 520608 610904
rect 463608 610784 463660 610836
rect 519636 610784 519688 610836
rect 430488 610716 430540 610768
rect 520648 610716 520700 610768
rect 365628 610648 365680 610700
rect 520740 610648 520792 610700
rect 332508 610580 332560 610632
rect 519728 610580 519780 610632
rect 379980 610376 380032 610428
rect 496452 610376 496504 610428
rect 3424 610308 3476 610360
rect 520832 610308 520884 610360
rect 542452 608540 542504 608592
rect 542544 608540 542596 608592
rect 389088 605820 389140 605872
rect 416780 605820 416832 605872
rect 387708 604460 387760 604512
rect 416780 604460 416832 604512
rect 384948 603100 385000 603152
rect 416780 603100 416832 603152
rect 538864 603100 538916 603152
rect 580172 603100 580224 603152
rect 383568 601672 383620 601724
rect 416780 601672 416832 601724
rect 542452 601672 542504 601724
rect 542728 601672 542780 601724
rect 380808 600312 380860 600364
rect 416780 600312 416832 600364
rect 378048 598952 378100 599004
rect 416780 598952 416832 599004
rect 542544 598884 542596 598936
rect 542728 598884 542780 598936
rect 410524 597524 410576 597576
rect 416780 597524 416832 597576
rect 556804 592016 556856 592068
rect 580172 592016 580224 592068
rect 542544 589296 542596 589348
rect 542820 589296 542872 589348
rect 542820 582428 542872 582480
rect 542728 582292 542780 582344
rect 523684 579640 523736 579692
rect 580172 579640 580224 579692
rect 542452 563116 542504 563168
rect 542452 562980 542504 563032
rect 537484 556180 537536 556232
rect 580172 556180 580224 556232
rect 542360 553392 542412 553444
rect 542452 553324 542504 553376
rect 542360 550604 542412 550656
rect 542452 550604 542504 550656
rect 555424 545096 555476 545148
rect 580172 545096 580224 545148
rect 542360 543736 542412 543788
rect 542452 543600 542504 543652
rect 411168 539588 411220 539640
rect 416780 539588 416832 539640
rect 379520 538228 379572 538280
rect 379796 538228 379848 538280
rect 409144 538228 409196 538280
rect 416780 538228 416832 538280
rect 379520 536052 379572 536104
rect 379796 536052 379848 536104
rect 542452 534012 542504 534064
rect 542636 534012 542688 534064
rect 523776 532720 523828 532772
rect 580172 532720 580224 532772
rect 542636 524424 542688 524476
rect 542728 524356 542780 524408
rect 408500 521568 408552 521620
rect 409144 521568 409196 521620
rect 297272 520888 297324 520940
rect 408500 520888 408552 520940
rect 379612 519528 379664 519580
rect 379796 519528 379848 519580
rect 318708 518848 318760 518900
rect 327172 518848 327224 518900
rect 317328 518780 317380 518832
rect 325424 518780 325476 518832
rect 331220 518780 331272 518832
rect 340512 518780 340564 518832
rect 369860 518780 369912 518832
rect 379428 518780 379480 518832
rect 379520 518780 379572 518832
rect 388996 518780 389048 518832
rect 393320 518780 393372 518832
rect 402888 518780 402940 518832
rect 451280 518780 451332 518832
rect 459560 518780 459612 518832
rect 307576 518712 307628 518764
rect 324320 518712 324372 518764
rect 326436 518712 326488 518764
rect 335544 518712 335596 518764
rect 345480 518712 345532 518764
rect 441620 518712 441672 518764
rect 443184 518712 443236 518764
rect 452568 518712 452620 518764
rect 460940 518712 460992 518764
rect 314568 518644 314620 518696
rect 323124 518644 323176 518696
rect 332324 518644 332376 518696
rect 320088 518576 320140 518628
rect 328920 518576 328972 518628
rect 337200 518644 337252 518696
rect 346492 518644 346544 518696
rect 443000 518644 443052 518696
rect 453672 518644 453724 518696
rect 462320 518644 462372 518696
rect 317328 518508 317380 518560
rect 326436 518508 326488 518560
rect 327172 518508 327224 518560
rect 336648 518508 336700 518560
rect 341616 518576 341668 518628
rect 342168 518576 342220 518628
rect 347780 518576 347832 518628
rect 348608 518576 348660 518628
rect 350540 518576 350592 518628
rect 357440 518576 357492 518628
rect 362224 518576 362276 518628
rect 379428 518576 379480 518628
rect 379520 518576 379572 518628
rect 402888 518576 402940 518628
rect 432512 518576 432564 518628
rect 446588 518576 446640 518628
rect 456064 518576 456116 518628
rect 465080 518576 465132 518628
rect 338120 518508 338172 518560
rect 347688 518508 347740 518560
rect 445760 518508 445812 518560
rect 447416 518508 447468 518560
rect 456892 518508 456944 518560
rect 315948 518440 316000 518492
rect 324412 518440 324464 518492
rect 292488 518372 292540 518424
rect 316040 518372 316092 518424
rect 325424 518440 325476 518492
rect 334164 518440 334216 518492
rect 335176 518440 335228 518492
rect 362224 518440 362276 518492
rect 369860 518440 369912 518492
rect 388996 518440 389048 518492
rect 393320 518440 393372 518492
rect 448796 518440 448848 518492
rect 458272 518440 458324 518492
rect 466552 518440 466604 518492
rect 333428 518372 333480 518424
rect 342996 518372 343048 518424
rect 343548 518372 343600 518424
rect 350540 518372 350592 518424
rect 357440 518372 357492 518424
rect 373908 518372 373960 518424
rect 426440 518372 426492 518424
rect 445392 518372 445444 518424
rect 455328 518372 455380 518424
rect 456892 518372 456944 518424
rect 466460 518372 466512 518424
rect 295248 518304 295300 518356
rect 317420 518304 317472 518356
rect 321100 518304 321152 518356
rect 330116 518304 330168 518356
rect 339960 518304 340012 518356
rect 347780 518304 347832 518356
rect 362868 518304 362920 518356
rect 430580 518304 430632 518356
rect 432512 518304 432564 518356
rect 447140 518304 447192 518356
rect 449900 518304 449952 518356
rect 459560 518304 459612 518356
rect 467840 518304 467892 518356
rect 313188 518236 313240 518288
rect 321744 518236 321796 518288
rect 331220 518236 331272 518288
rect 335176 518236 335228 518288
rect 344192 518236 344244 518288
rect 344928 518236 344980 518288
rect 361488 518236 361540 518288
rect 429292 518236 429344 518288
rect 432604 518236 432656 518288
rect 442080 518236 442132 518288
rect 303620 518168 303672 518220
rect 423680 518168 423732 518220
rect 444288 518236 444340 518288
rect 453672 518236 453724 518288
rect 455328 518236 455380 518288
rect 463700 518236 463752 518288
rect 451280 518168 451332 518220
rect 306288 518100 306340 518152
rect 322940 518100 322992 518152
rect 358728 518100 358780 518152
rect 429200 518100 429252 518152
rect 303528 518032 303580 518084
rect 321836 518032 321888 518084
rect 355968 518032 356020 518084
rect 425612 518032 425664 518084
rect 435916 518032 435968 518084
rect 444288 518032 444340 518084
rect 299388 517964 299440 518016
rect 318800 517964 318852 518016
rect 296628 517896 296680 517948
rect 317512 517896 317564 517948
rect 285588 517828 285640 517880
rect 312084 517828 312136 517880
rect 314568 517828 314620 517880
rect 327080 517964 327132 518016
rect 340512 517964 340564 518016
rect 431960 517964 432012 518016
rect 300676 517760 300728 517812
rect 320180 517760 320232 517812
rect 321468 517760 321520 517812
rect 331220 517896 331272 517948
rect 343548 517896 343600 517948
rect 436100 517896 436152 517948
rect 436744 517896 436796 517948
rect 437296 517896 437348 517948
rect 446588 517896 446640 517948
rect 280896 517692 280948 517744
rect 303620 517692 303672 517744
rect 310428 517692 310480 517744
rect 288348 517624 288400 517676
rect 313280 517624 313332 517676
rect 322848 517692 322900 517744
rect 332600 517828 332652 517880
rect 433892 517828 433944 517880
rect 443184 517828 443236 517880
rect 438124 517760 438176 517812
rect 447416 517760 447468 517812
rect 328368 517692 328420 517744
rect 333980 517692 334032 517744
rect 440884 517692 440936 517744
rect 449900 517692 449952 517744
rect 324320 517624 324372 517676
rect 326344 517624 326396 517676
rect 329840 517624 329892 517676
rect 330484 517624 330536 517676
rect 335728 517624 335780 517676
rect 344928 517624 344980 517676
rect 438860 517624 438912 517676
rect 439504 517624 439556 517676
rect 448796 517624 448848 517676
rect 289728 517556 289780 517608
rect 314660 517556 314712 517608
rect 317328 517556 317380 517608
rect 311808 517488 311860 517540
rect 325700 517488 325752 517540
rect 327724 517556 327776 517608
rect 332600 517556 332652 517608
rect 333888 517556 333940 517608
rect 338120 517556 338172 517608
rect 342168 517556 342220 517608
rect 434720 517556 434772 517608
rect 436652 517556 436704 517608
rect 436928 517556 436980 517608
rect 445392 517556 445444 517608
rect 328460 517488 328512 517540
rect 333244 517488 333296 517540
rect 336740 517488 336792 517540
rect 337384 517488 337436 517540
rect 339500 517488 339552 517540
rect 379612 514020 379664 514072
rect 379796 514020 379848 514072
rect 542544 511980 542596 512032
rect 542820 511980 542872 512032
rect 433800 511912 433852 511964
rect 433892 511912 433944 511964
rect 3332 509260 3384 509312
rect 520004 509260 520056 509312
rect 536104 509260 536156 509312
rect 580172 509260 580224 509312
rect 433800 502324 433852 502376
rect 434076 502324 434128 502376
rect 542636 502324 542688 502376
rect 542820 502324 542872 502376
rect 379612 499536 379664 499588
rect 379796 499536 379848 499588
rect 554044 498176 554096 498228
rect 580172 498176 580224 498228
rect 3424 495456 3476 495508
rect 521292 495456 521344 495508
rect 379612 494708 379664 494760
rect 379796 494708 379848 494760
rect 433616 492600 433668 492652
rect 433892 492600 433944 492652
rect 542544 492600 542596 492652
rect 542636 492600 542688 492652
rect 523868 485800 523920 485852
rect 580172 485800 580224 485852
rect 542544 485732 542596 485784
rect 542636 485732 542688 485784
rect 297824 482944 297876 482996
rect 299572 482944 299624 482996
rect 307668 482944 307720 482996
rect 297456 482876 297508 482928
rect 428832 482944 428884 482996
rect 439504 482944 439556 482996
rect 455328 482944 455380 482996
rect 492036 482944 492088 482996
rect 283472 482808 283524 482860
rect 379704 482808 379756 482860
rect 390744 482876 390796 482928
rect 426164 482876 426216 482928
rect 438124 482876 438176 482928
rect 453856 482876 453908 482928
rect 489920 482876 489972 482928
rect 387616 482808 387668 482860
rect 433248 482808 433300 482860
rect 450268 482808 450320 482860
rect 458088 482808 458140 482860
rect 496452 482808 496504 482860
rect 297548 482740 297600 482792
rect 387340 482740 387392 482792
rect 434628 482740 434680 482792
rect 452660 482740 452712 482792
rect 456708 482740 456760 482792
rect 494244 482740 494296 482792
rect 281356 482672 281408 482724
rect 379796 482672 379848 482724
rect 382648 482672 382700 482724
rect 383568 482672 383620 482724
rect 386972 482672 387024 482724
rect 387708 482672 387760 482724
rect 436008 482672 436060 482724
rect 454592 482672 454644 482724
rect 459468 482672 459520 482724
rect 498660 482672 498712 482724
rect 297640 482604 297692 482656
rect 397460 482604 397512 482656
rect 437388 482604 437440 482656
rect 456892 482604 456944 482656
rect 460848 482604 460900 482656
rect 500960 482604 501012 482656
rect 287888 482536 287940 482588
rect 288348 482536 288400 482588
rect 294512 482536 294564 482588
rect 295248 482536 295300 482588
rect 298928 482536 298980 482588
rect 299388 482536 299440 482588
rect 297732 482468 297784 482520
rect 399576 482536 399628 482588
rect 424416 482536 424468 482588
rect 436744 482536 436796 482588
rect 438676 482536 438728 482588
rect 459008 482536 459060 482588
rect 460756 482536 460808 482588
rect 503076 482536 503128 482588
rect 299572 482468 299624 482520
rect 401784 482468 401836 482520
rect 420000 482468 420052 482520
rect 435364 482468 435416 482520
rect 438768 482468 438820 482520
rect 461216 482468 461268 482520
rect 462228 482468 462280 482520
rect 505284 482468 505336 482520
rect 297916 482400 297968 482452
rect 403992 482400 404044 482452
rect 422208 482400 422260 482452
rect 436928 482400 436980 482452
rect 440148 482400 440200 482452
rect 463700 482400 463752 482452
rect 464988 482400 465040 482452
rect 509700 482400 509752 482452
rect 298008 482332 298060 482384
rect 406200 482332 406252 482384
rect 417792 482332 417844 482384
rect 433800 482332 433852 482384
rect 441528 482332 441580 482384
rect 465632 482332 465684 482384
rect 466368 482332 466420 482384
rect 512000 482332 512052 482384
rect 297364 482264 297416 482316
rect 412824 482264 412876 482316
rect 415216 482264 415268 482316
rect 432604 482264 432656 482316
rect 442908 482264 442960 482316
rect 467840 482264 467892 482316
rect 469128 482264 469180 482316
rect 516324 482264 516376 482316
rect 305552 482196 305604 482248
rect 306288 482196 306340 482248
rect 309968 482196 310020 482248
rect 310428 482196 310480 482248
rect 311716 482196 311768 482248
rect 371240 482196 371292 482248
rect 376024 482196 376076 482248
rect 410524 482196 410576 482248
rect 431040 482196 431092 482248
rect 440884 482196 440936 482248
rect 453948 482196 454000 482248
rect 487620 482196 487672 482248
rect 310244 482128 310296 482180
rect 368756 482128 368808 482180
rect 387616 482128 387668 482180
rect 392952 482128 393004 482180
rect 452568 482128 452620 482180
rect 485780 482128 485832 482180
rect 310336 482060 310388 482112
rect 366548 482060 366600 482112
rect 451188 482060 451240 482112
rect 483296 482060 483348 482112
rect 309048 481992 309100 482044
rect 364340 481992 364392 482044
rect 448428 481992 448480 482044
rect 478880 481992 478932 482044
rect 316500 481924 316552 481976
rect 317328 481924 317380 481976
rect 320916 481924 320968 481976
rect 321468 481924 321520 481976
rect 327540 481924 327592 481976
rect 328368 481924 328420 481976
rect 329748 481924 329800 481976
rect 330484 481924 330536 481976
rect 331956 481924 332008 481976
rect 333244 481924 333296 481976
rect 336372 481924 336424 481976
rect 337384 481924 337436 481976
rect 338580 481924 338632 481976
rect 339408 481924 339460 481976
rect 346308 481924 346360 481976
rect 346768 481924 346820 481976
rect 348424 481924 348476 481976
rect 349160 481924 349212 481976
rect 349252 481924 349304 481976
rect 351092 481924 351144 481976
rect 358268 481924 358320 481976
rect 358728 481924 358780 481976
rect 449808 481924 449860 481976
rect 481088 481924 481140 481976
rect 325332 481856 325384 481908
rect 327724 481856 327776 481908
rect 360568 481856 360620 481908
rect 361488 481856 361540 481908
rect 445576 481856 445628 481908
rect 474740 481856 474792 481908
rect 318708 481788 318760 481840
rect 326344 481788 326396 481840
rect 348976 481788 349028 481840
rect 353300 481788 353352 481840
rect 447048 481788 447100 481840
rect 476672 481788 476724 481840
rect 445668 481720 445720 481772
rect 472256 481720 472308 481772
rect 444288 481652 444340 481704
rect 470048 481652 470100 481704
rect 2964 480224 3016 480276
rect 520188 480224 520240 480276
rect 387340 480088 387392 480140
rect 395482 480088 395534 480140
rect 367192 479816 367244 479868
rect 369952 479816 370004 479868
rect 398748 479816 398800 479868
rect 520096 479816 520148 479868
rect 300584 479748 300636 479800
rect 520924 479748 520976 479800
rect 235908 479680 235960 479732
rect 521016 479680 521068 479732
rect 171048 479612 171100 479664
rect 521108 479612 521160 479664
rect 106188 479544 106240 479596
rect 521200 479544 521252 479596
rect 3608 479476 3660 479528
rect 521384 479476 521436 479528
rect 50988 479408 51040 479460
rect 57796 479408 57848 479460
rect 128268 479408 128320 479460
rect 135168 479408 135220 479460
rect 278872 479408 278924 479460
rect 283564 479408 283616 479460
rect 466368 479408 466420 479460
rect 473268 479408 473320 479460
rect 147588 479340 147640 479392
rect 154488 479340 154540 479392
rect 166908 479340 166960 479392
rect 173808 479340 173860 479392
rect 186228 479340 186280 479392
rect 193128 479340 193180 479392
rect 205548 479340 205600 479392
rect 212448 479340 212500 479392
rect 224868 479340 224920 479392
rect 231768 479340 231820 479392
rect 244188 479340 244240 479392
rect 251088 479340 251140 479392
rect 485688 479340 485740 479392
rect 492588 479340 492640 479392
rect 57980 479272 58032 479324
rect 61844 479272 61896 479324
rect 309140 479272 309192 479324
rect 316776 479272 316828 479324
rect 279700 479136 279752 479188
rect 519912 479136 519964 479188
rect 279608 479068 279660 479120
rect 521568 479068 521620 479120
rect 279976 479000 280028 479052
rect 523132 479000 523184 479052
rect 135168 478932 135220 478984
rect 277400 478932 277452 478984
rect 279884 478932 279936 478984
rect 523040 478932 523092 478984
rect 3424 478864 3476 478916
rect 519820 478864 519872 478916
rect 520096 478728 520148 478780
rect 519912 478660 519964 478712
rect 279148 478524 279200 478576
rect 520188 478524 520240 478576
rect 280068 478456 280120 478508
rect 521476 478456 521528 478508
rect 279792 478388 279844 478440
rect 522672 478388 522724 478440
rect 279516 478320 279568 478372
rect 522856 478320 522908 478372
rect 3792 478252 3844 478304
rect 522488 478252 522540 478304
rect 3516 478184 3568 478236
rect 522304 478184 522356 478236
rect 3700 478116 3752 478168
rect 522580 478116 522632 478168
rect 279240 478048 279292 478100
rect 522764 478048 522816 478100
rect 279424 477980 279476 478032
rect 522396 477980 522448 478032
rect 279332 477912 279384 477964
rect 524420 477912 524472 477964
rect 133788 476076 133840 476128
rect 277400 476076 277452 476128
rect 542452 476076 542504 476128
rect 542636 476076 542688 476128
rect 132408 473356 132460 473408
rect 278688 473356 278740 473408
rect 542544 473288 542596 473340
rect 542636 473288 542688 473340
rect 131028 471996 131080 472048
rect 278688 471996 278740 472048
rect 129648 469208 129700 469260
rect 277860 469208 277912 469260
rect 128268 467848 128320 467900
rect 278688 467848 278740 467900
rect 542636 466420 542688 466472
rect 542544 466352 542596 466404
rect 126888 465060 126940 465112
rect 278688 465060 278740 465112
rect 125508 463700 125560 463752
rect 278688 463700 278740 463752
rect 549904 462340 549956 462392
rect 580172 462340 580224 462392
rect 125416 460912 125468 460964
rect 278688 460912 278740 460964
rect 124128 459552 124180 459604
rect 278688 459552 278740 459604
rect 122748 456764 122800 456816
rect 278688 456764 278740 456816
rect 121368 455404 121420 455456
rect 278688 455404 278740 455456
rect 119988 452616 120040 452668
rect 278688 452616 278740 452668
rect 3516 452548 3568 452600
rect 279148 452548 279200 452600
rect 118608 451256 118660 451308
rect 278688 451256 278740 451308
rect 563704 451256 563756 451308
rect 580172 451256 580224 451308
rect 117228 448536 117280 448588
rect 278688 448536 278740 448588
rect 542360 447108 542412 447160
rect 542452 447040 542504 447092
rect 117136 445748 117188 445800
rect 278688 445748 278740 445800
rect 115848 444388 115900 444440
rect 278688 444388 278740 444440
rect 542176 444320 542228 444372
rect 542452 444320 542504 444372
rect 114468 441600 114520 441652
rect 277860 441600 277912 441652
rect 113088 440240 113140 440292
rect 278688 440240 278740 440292
rect 534724 438880 534776 438932
rect 580172 438880 580224 438932
rect 3516 438812 3568 438864
rect 279240 438812 279292 438864
rect 522212 437588 522264 437640
rect 111708 437452 111760 437504
rect 278688 437452 278740 437504
rect 519820 437452 519872 437504
rect 522212 437452 522264 437504
rect 522948 437452 523000 437504
rect 110328 436092 110380 436144
rect 278044 436092 278096 436144
rect 108948 433304 109000 433356
rect 278688 433304 278740 433356
rect 107568 431944 107620 431996
rect 278688 431944 278740 431996
rect 107476 429156 107528 429208
rect 277676 429156 277728 429208
rect 106188 427796 106240 427848
rect 278688 427796 278740 427848
rect 542360 427796 542412 427848
rect 542452 427728 542504 427780
rect 104808 425076 104860 425128
rect 278688 425076 278740 425128
rect 3240 425008 3292 425060
rect 279332 425008 279384 425060
rect 542176 425008 542228 425060
rect 542452 425008 542504 425060
rect 103428 423648 103480 423700
rect 278688 423648 278740 423700
rect 102048 420928 102100 420980
rect 278688 420928 278740 420980
rect 522672 420044 522724 420096
rect 524420 420044 524472 420096
rect 100668 418140 100720 418192
rect 278688 418140 278740 418192
rect 99288 416780 99340 416832
rect 278688 416780 278740 416832
rect 547144 415420 547196 415472
rect 580172 415420 580224 415472
rect 99196 413992 99248 414044
rect 277860 413992 277912 414044
rect 97908 412632 97960 412684
rect 278688 412632 278740 412684
rect 96528 409844 96580 409896
rect 278688 409844 278740 409896
rect 95148 408484 95200 408536
rect 278688 408484 278740 408536
rect 542360 408484 542412 408536
rect 542452 408348 542504 408400
rect 93768 405696 93820 405748
rect 278688 405696 278740 405748
rect 92388 404336 92440 404388
rect 278688 404336 278740 404388
rect 542084 404268 542136 404320
rect 542452 404268 542504 404320
rect 91008 401616 91060 401668
rect 278412 401616 278464 401668
rect 90916 400188 90968 400240
rect 278688 400188 278740 400240
rect 89628 397468 89680 397520
rect 278688 397468 278740 397520
rect 88248 396040 88300 396092
rect 278688 396040 278740 396092
rect 3148 395972 3200 396024
rect 280068 395972 280120 396024
rect 86868 393320 86920 393372
rect 278688 393320 278740 393372
rect 542176 393252 542228 393304
rect 542360 393252 542412 393304
rect 523960 391960 524012 392012
rect 579896 391960 579948 392012
rect 85488 390532 85540 390584
rect 278320 390532 278372 390584
rect 84108 389172 84160 389224
rect 278688 389172 278740 389224
rect 82728 386384 82780 386436
rect 277860 386384 277912 386436
rect 82636 385024 82688 385076
rect 277676 385024 277728 385076
rect 542176 383664 542228 383716
rect 542452 383664 542504 383716
rect 81348 382236 81400 382288
rect 278688 382236 278740 382288
rect 79968 380876 80020 380928
rect 278044 380876 278096 380928
rect 3516 380808 3568 380860
rect 279976 380808 280028 380860
rect 542452 379448 542504 379500
rect 542636 379448 542688 379500
rect 78588 378156 78640 378208
rect 278688 378156 278740 378208
rect 77208 376728 77260 376780
rect 278688 376728 278740 376780
rect 75828 374008 75880 374060
rect 278412 374008 278464 374060
rect 74448 372580 74500 372632
rect 278044 372580 278096 372632
rect 73068 369860 73120 369912
rect 278320 369860 278372 369912
rect 72976 368500 73028 368552
rect 278688 368500 278740 368552
rect 3516 367004 3568 367056
rect 279884 367004 279936 367056
rect 542452 367004 542504 367056
rect 542728 367004 542780 367056
rect 71688 365712 71740 365764
rect 278688 365712 278740 365764
rect 70308 362924 70360 362976
rect 277860 362924 277912 362976
rect 68928 361564 68980 361616
rect 278688 361564 278740 361616
rect 67548 358776 67600 358828
rect 277860 358776 277912 358828
rect 66168 357416 66220 357468
rect 278688 357416 278740 357468
rect 542452 357416 542504 357468
rect 542544 357416 542596 357468
rect 64788 354696 64840 354748
rect 278688 354696 278740 354748
rect 64696 353268 64748 353320
rect 278044 353268 278096 353320
rect 63408 350548 63460 350600
rect 278688 350548 278740 350600
rect 542544 350548 542596 350600
rect 542728 350480 542780 350532
rect 62028 349120 62080 349172
rect 278688 349120 278740 349172
rect 60648 346400 60700 346452
rect 278688 346400 278740 346452
rect 59268 345040 59320 345092
rect 278688 345040 278740 345092
rect 57888 342252 57940 342304
rect 278320 342252 278372 342304
rect 56508 340892 56560 340944
rect 278688 340892 278740 340944
rect 522948 340824 523000 340876
rect 542728 340824 542780 340876
rect 56416 338104 56468 338156
rect 278688 338104 278740 338156
rect 3516 338036 3568 338088
rect 279792 338036 279844 338088
rect 522948 337900 523000 337952
rect 527180 337900 527232 337952
rect 522580 336676 522632 336728
rect 531964 336676 532016 336728
rect 55128 335316 55180 335368
rect 277860 335316 277912 335368
rect 53748 333956 53800 334008
rect 278688 333956 278740 334008
rect 522948 333888 523000 333940
rect 560944 333888 560996 333940
rect 522580 332528 522632 332580
rect 545764 332528 545816 332580
rect 52368 331236 52420 331288
rect 278688 331236 278740 331288
rect 50988 329808 51040 329860
rect 278688 329808 278740 329860
rect 522948 328516 523000 328568
rect 529204 328516 529256 328568
rect 522948 328380 523000 328432
rect 558184 328380 558236 328432
rect 49608 327088 49660 327140
rect 278688 327088 278740 327140
rect 48228 325660 48280 325712
rect 278044 325660 278096 325712
rect 522948 325592 523000 325644
rect 540244 325592 540296 325644
rect 3516 324232 3568 324284
rect 279700 324232 279752 324284
rect 522304 324096 522356 324148
rect 525064 324096 525116 324148
rect 48136 322940 48188 322992
rect 277676 322940 277728 322992
rect 46848 321580 46900 321632
rect 278044 321580 278096 321632
rect 522672 321512 522724 321564
rect 556804 321512 556856 321564
rect 522948 320084 523000 320136
rect 538864 320084 538916 320136
rect 45468 318792 45520 318844
rect 278688 318792 278740 318844
rect 44088 317432 44140 317484
rect 278688 317432 278740 317484
rect 522304 316888 522356 316940
rect 523684 316888 523736 316940
rect 42708 314644 42760 314696
rect 278688 314644 278740 314696
rect 522948 314576 523000 314628
rect 555424 314576 555476 314628
rect 41328 313284 41380 313336
rect 278688 313284 278740 313336
rect 522948 313216 523000 313268
rect 537484 313216 537536 313268
rect 39948 310496 40000 310548
rect 278688 310496 278740 310548
rect 522304 310428 522356 310480
rect 523776 310428 523828 310480
rect 3332 309068 3384 309120
rect 279608 309068 279660 309120
rect 522948 309068 523000 309120
rect 554044 309068 554096 309120
rect 38568 307776 38620 307828
rect 277860 307776 277912 307828
rect 38476 306348 38528 306400
rect 278688 306348 278740 306400
rect 522948 306280 523000 306332
rect 536104 306280 536156 306332
rect 522304 304784 522356 304836
rect 523868 304784 523920 304836
rect 37188 303628 37240 303680
rect 278688 303628 278740 303680
rect 35808 302200 35860 302252
rect 278688 302200 278740 302252
rect 522948 302132 523000 302184
rect 563704 302132 563756 302184
rect 522948 300772 523000 300824
rect 549904 300772 549956 300824
rect 34428 299480 34480 299532
rect 278688 299480 278740 299532
rect 33048 298120 33100 298172
rect 278688 298120 278740 298172
rect 522948 298052 523000 298104
rect 534724 298052 534776 298104
rect 522948 296624 523000 296676
rect 580264 296624 580316 296676
rect 31668 295332 31720 295384
rect 278688 295332 278740 295384
rect 3056 295264 3108 295316
rect 279516 295264 279568 295316
rect 522488 294652 522540 294704
rect 580724 294652 580776 294704
rect 522304 294584 522356 294636
rect 579988 294584 580040 294636
rect 30288 293972 30340 294024
rect 278688 293972 278740 294024
rect 522948 293904 523000 293956
rect 547144 293904 547196 293956
rect 522580 292000 522632 292052
rect 523960 292000 524012 292052
rect 30196 291184 30248 291236
rect 278688 291184 278740 291236
rect 28908 289824 28960 289876
rect 278688 289824 278740 289876
rect 522948 289756 523000 289808
rect 580448 289756 580500 289808
rect 522580 288328 522632 288380
rect 580356 288328 580408 288380
rect 27528 287036 27580 287088
rect 278688 287036 278740 287088
rect 26148 285676 26200 285728
rect 278688 285676 278740 285728
rect 522580 285608 522632 285660
rect 580540 285608 580592 285660
rect 24768 282888 24820 282940
rect 278688 282888 278740 282940
rect 522948 281460 523000 281512
rect 580632 281460 580684 281512
rect 23388 280168 23440 280220
rect 277860 280168 277912 280220
rect 3516 280100 3568 280152
rect 279424 280100 279476 280152
rect 22008 278740 22060 278792
rect 278688 278740 278740 278792
rect 21916 276020 21968 276072
rect 278688 276020 278740 276072
rect 522948 275272 523000 275324
rect 580172 275272 580224 275324
rect 20628 274660 20680 274712
rect 278044 274660 278096 274712
rect 19248 271872 19300 271924
rect 278688 271872 278740 271924
rect 17868 270512 17920 270564
rect 278688 270512 278740 270564
rect 16488 267724 16540 267776
rect 278688 267724 278740 267776
rect 15108 266364 15160 266416
rect 278044 266364 278096 266416
rect 522488 265616 522540 265668
rect 580172 265616 580224 265668
rect 522580 264936 522632 264988
rect 523960 264936 524012 264988
rect 13728 263576 13780 263628
rect 278688 263576 278740 263628
rect 13636 262216 13688 262268
rect 278688 262216 278740 262268
rect 522580 260856 522632 260908
rect 523868 260856 523920 260908
rect 12348 259428 12400 259480
rect 278320 259428 278372 259480
rect 522580 259428 522632 259480
rect 523776 259428 523828 259480
rect 10968 256708 11020 256760
rect 277860 256708 277912 256760
rect 9588 255280 9640 255332
rect 278688 255280 278740 255332
rect 8208 252560 8260 252612
rect 277860 252560 277912 252612
rect 522304 252492 522356 252544
rect 579804 252492 579856 252544
rect 6828 251200 6880 251252
rect 278688 251200 278740 251252
rect 5448 248412 5500 248464
rect 278688 248412 278740 248464
rect 522304 248412 522356 248464
rect 531964 248412 532016 248464
rect 522304 247052 522356 247104
rect 527824 247052 527876 247104
rect 522396 243176 522448 243228
rect 2688 242904 2740 242956
rect 277400 242904 277452 242956
rect 522396 242904 522448 242956
rect 529204 242904 529256 242956
rect 522396 242768 522448 242820
rect 3516 240864 3568 240916
rect 522396 240864 522448 240916
rect 3608 240796 3660 240848
rect 519820 240796 519872 240848
rect 280160 240660 280212 240712
rect 280896 240660 280948 240712
rect 306380 240660 306432 240712
rect 315948 240660 316000 240712
rect 325608 240660 325660 240712
rect 316040 240592 316092 240644
rect 340880 240660 340932 240712
rect 350448 240660 350500 240712
rect 340788 240592 340840 240644
rect 350632 240592 350684 240644
rect 357440 240592 357492 240644
rect 360384 240592 360436 240644
rect 369676 240660 369728 240712
rect 306380 240456 306432 240508
rect 315948 240456 316000 240508
rect 369676 240388 369728 240440
rect 373264 240388 373316 240440
rect 1308 240116 1360 240168
rect 278688 240116 278740 240168
rect 522396 240116 522448 240168
rect 525064 240116 525116 240168
rect 333704 238688 333756 238740
rect 344560 238688 344612 238740
rect 426348 238688 426400 238740
rect 450544 238688 450596 238740
rect 459468 238688 459520 238740
rect 474004 238688 474056 238740
rect 475568 238688 475620 238740
rect 489920 238688 489972 238740
rect 332508 238620 332560 238672
rect 346768 238620 346820 238672
rect 424416 238620 424468 238672
rect 452016 238620 452068 238672
rect 463608 238620 463660 238672
rect 492036 238620 492088 238672
rect 331128 238552 331180 238604
rect 349160 238552 349212 238604
rect 422208 238552 422260 238604
rect 453304 238552 453356 238604
rect 462228 238552 462280 238604
rect 494244 238552 494296 238604
rect 329564 238484 329616 238536
rect 351092 238484 351144 238536
rect 380440 238484 380492 238536
rect 395160 238484 395212 238536
rect 417884 238484 417936 238536
rect 456248 238484 456300 238536
rect 459468 238484 459520 238536
rect 498660 238484 498712 238536
rect 294512 238416 294564 238468
rect 295248 238416 295300 238468
rect 328368 238416 328420 238468
rect 353300 238416 353352 238468
rect 380348 238416 380400 238468
rect 397460 238416 397512 238468
rect 415308 238416 415360 238468
rect 456064 238416 456116 238468
rect 456708 238416 456760 238468
rect 503076 238416 503128 238468
rect 311808 238348 311860 238400
rect 342904 238348 342956 238400
rect 380256 238348 380308 238400
rect 399576 238348 399628 238400
rect 420000 238348 420052 238400
rect 454684 238348 454736 238400
rect 455144 238348 455196 238400
rect 507492 238348 507544 238400
rect 309968 238280 310020 238332
rect 344284 238280 344336 238332
rect 389088 238280 389140 238332
rect 451924 238280 451976 238332
rect 452568 238280 452620 238332
rect 512092 238280 512144 238332
rect 305552 238212 305604 238264
rect 342996 238212 343048 238264
rect 371148 238212 371200 238264
rect 390744 238212 390796 238264
rect 395344 238212 395396 238264
rect 406200 238212 406252 238264
rect 428832 238212 428884 238264
rect 449164 238212 449216 238264
rect 449808 238212 449860 238264
rect 516324 238212 516376 238264
rect 283472 238144 283524 238196
rect 297824 238144 297876 238196
rect 303344 238144 303396 238196
rect 341524 238144 341576 238196
rect 380532 238144 380584 238196
rect 412824 238144 412876 238196
rect 431040 238144 431092 238196
rect 447784 238144 447836 238196
rect 448428 238144 448480 238196
rect 518532 238144 518584 238196
rect 281356 238076 281408 238128
rect 297364 238076 297416 238128
rect 307668 238076 307720 238128
rect 347044 238076 347096 238128
rect 380164 238076 380216 238128
rect 403992 238076 404044 238128
rect 411168 238076 411220 238128
rect 496360 238076 496412 238128
rect 285588 238008 285640 238060
rect 345664 238008 345716 238060
rect 360568 238008 360620 238060
rect 476764 238008 476816 238060
rect 461860 237940 461912 237992
rect 474096 237940 474148 237992
rect 475476 237940 475528 237992
rect 487620 237940 487672 237992
rect 464068 237872 464120 237924
rect 475384 237872 475436 237924
rect 335176 237804 335228 237856
rect 342352 237804 342404 237856
rect 470508 237804 470560 237856
rect 473360 237804 473412 237856
rect 474280 237804 474332 237856
rect 485780 237804 485832 237856
rect 466276 237736 466328 237788
rect 475660 237736 475712 237788
rect 331956 237668 332008 237720
rect 339592 237668 339644 237720
rect 474188 237668 474240 237720
rect 483296 237668 483348 237720
rect 335268 237600 335320 237652
rect 340144 237600 340196 237652
rect 468484 237600 468536 237652
rect 474832 237600 474884 237652
rect 333888 237532 333940 237584
rect 338212 237532 338264 237584
rect 287888 237396 287940 237448
rect 288348 237396 288400 237448
rect 298928 237396 298980 237448
rect 299388 237396 299440 237448
rect 316500 237396 316552 237448
rect 317328 237396 317380 237448
rect 320916 237396 320968 237448
rect 321468 237396 321520 237448
rect 327540 237396 327592 237448
rect 328276 237396 328328 237448
rect 329748 237396 329800 237448
rect 337384 237464 337436 237516
rect 367008 237464 367060 237516
rect 371240 237464 371292 237516
rect 333704 237396 333756 237448
rect 333888 237396 333940 237448
rect 336556 237396 336608 237448
rect 338120 237396 338172 237448
rect 364984 237396 365036 237448
rect 366364 237396 366416 237448
rect 366916 237396 366968 237448
rect 368756 237396 368808 237448
rect 376024 237396 376076 237448
rect 376668 237396 376720 237448
rect 382648 237396 382700 237448
rect 383568 237396 383620 237448
rect 386972 237396 387024 237448
rect 387708 237396 387760 237448
rect 391204 237396 391256 237448
rect 392952 237396 393004 237448
rect 393964 237396 394016 237448
rect 401784 237396 401836 237448
rect 453028 237396 453080 237448
rect 453948 237396 454000 237448
rect 457444 237396 457496 237448
rect 458088 237396 458140 237448
rect 471888 237396 471940 237448
rect 474740 237396 474792 237448
rect 3516 237328 3568 237380
rect 522120 237328 522172 237380
rect 329564 234540 329616 234592
rect 329748 234540 329800 234592
rect 431960 232160 432012 232212
rect 432696 232160 432748 232212
rect 336372 230460 336424 230512
rect 336556 230460 336608 230512
rect 522948 229032 523000 229084
rect 580172 229032 580224 229084
rect 3148 223524 3200 223576
rect 522212 223524 522264 223576
rect 336372 222232 336424 222284
rect 336648 222232 336700 222284
rect 329472 222164 329524 222216
rect 329656 222164 329708 222216
rect 431776 222164 431828 222216
rect 432052 222164 432104 222216
rect 522856 217948 522908 218000
rect 580172 217948 580224 218000
rect 432052 215364 432104 215416
rect 432144 215296 432196 215348
rect 3516 208292 3568 208344
rect 522028 208292 522080 208344
rect 523960 205572 524012 205624
rect 579804 205572 579856 205624
rect 470508 205232 470560 205284
rect 476120 205232 476172 205284
rect 470416 205096 470468 205148
rect 478880 205096 478932 205148
rect 469128 205028 469180 205080
rect 480260 205028 480312 205080
rect 451188 204960 451240 205012
rect 484400 204960 484452 205012
rect 373908 204892 373960 204944
rect 490196 204892 490248 204944
rect 347780 204280 347832 204332
rect 357348 204280 357400 204332
rect 389824 204280 389876 204332
rect 394424 204280 394476 204332
rect 317328 204212 317380 204264
rect 342812 204212 342864 204264
rect 299388 204144 299440 204196
rect 347044 204212 347096 204264
rect 351920 204212 351972 204264
rect 374644 204212 374696 204264
rect 379520 204212 379572 204264
rect 416044 204212 416096 204264
rect 427820 204212 427872 204264
rect 452016 204212 452068 204264
rect 461492 204212 461544 204264
rect 464988 204212 465040 204264
rect 475476 204212 475528 204264
rect 476764 204212 476816 204264
rect 485780 204212 485832 204264
rect 357440 204144 357492 204196
rect 357992 204144 358044 204196
rect 394516 204144 394568 204196
rect 394608 204144 394660 204196
rect 412548 204144 412600 204196
rect 412640 204144 412692 204196
rect 445760 204144 445812 204196
rect 450544 204144 450596 204196
rect 450912 204144 450964 204196
rect 460664 204144 460716 204196
rect 466276 204144 466328 204196
rect 474280 204144 474332 204196
rect 475384 204144 475436 204196
rect 477500 204144 477552 204196
rect 330944 204076 330996 204128
rect 337292 204076 337344 204128
rect 337384 204076 337436 204128
rect 340972 204076 341024 204128
rect 342812 204076 342864 204128
rect 347780 204076 347832 204128
rect 354036 204076 354088 204128
rect 358636 204076 358688 204128
rect 364984 204076 365036 204128
rect 367100 204076 367152 204128
rect 376576 204076 376628 204128
rect 379520 204076 379572 204128
rect 389824 204076 389876 204128
rect 394424 204076 394476 204128
rect 402888 204076 402940 204128
rect 402980 204076 403032 204128
rect 416044 204076 416096 204128
rect 427912 204076 427964 204128
rect 443000 204076 443052 204128
rect 449164 204076 449216 204128
rect 459100 204076 459152 204128
rect 467288 204076 467340 204128
rect 475752 204076 475804 204128
rect 475844 204076 475896 204128
rect 483020 204076 483072 204128
rect 300768 204008 300820 204060
rect 356060 204008 356112 204060
rect 360016 204008 360068 204060
rect 441620 204008 441672 204060
rect 447784 204008 447836 204060
rect 448428 204008 448480 204060
rect 457904 204008 457956 204060
rect 457996 204008 458048 204060
rect 500960 204008 501012 204060
rect 314568 203940 314620 203992
rect 349160 203940 349212 203992
rect 333796 203872 333848 203924
rect 341708 203872 341760 203924
rect 318708 203804 318760 203856
rect 335084 203804 335136 203856
rect 321468 203736 321520 203788
rect 345020 203804 345072 203856
rect 335820 203736 335872 203788
rect 322848 203668 322900 203720
rect 336004 203668 336056 203720
rect 337292 203736 337344 203788
rect 340052 203736 340104 203788
rect 349436 203872 349488 203924
rect 354036 203872 354088 203924
rect 361304 203940 361356 203992
rect 438860 203940 438912 203992
rect 460848 203940 460900 203992
rect 495440 203940 495492 203992
rect 345572 203804 345624 203856
rect 351644 203804 351696 203856
rect 362868 203872 362920 203924
rect 436100 203872 436152 203924
rect 453948 203872 454000 203924
rect 483020 203872 483072 203924
rect 354588 203804 354640 203856
rect 363420 203804 363472 203856
rect 434720 203804 434772 203856
rect 455236 203804 455288 203856
rect 471060 203804 471112 203856
rect 474096 203804 474148 203856
rect 477500 203804 477552 203856
rect 345664 203736 345716 203788
rect 364340 203736 364392 203788
rect 337936 203668 337988 203720
rect 340696 203668 340748 203720
rect 325608 203600 325660 203652
rect 331220 203600 331272 203652
rect 340604 203600 340656 203652
rect 342260 203668 342312 203720
rect 342812 203668 342864 203720
rect 343640 203668 343692 203720
rect 353024 203668 353076 203720
rect 362868 203668 362920 203720
rect 341524 203600 341576 203652
rect 354680 203600 354732 203652
rect 355600 203600 355652 203652
rect 365076 203600 365128 203652
rect 369860 203600 369912 203652
rect 376300 203600 376352 203652
rect 408592 203668 408644 203720
rect 408684 203668 408736 203720
rect 328276 203532 328328 203584
rect 342260 203532 342312 203584
rect 342720 203532 342772 203584
rect 348424 203532 348476 203584
rect 357992 203532 358044 203584
rect 364984 203532 365036 203584
rect 374644 203532 374696 203584
rect 432144 203736 432196 203788
rect 458088 203736 458140 203788
rect 470784 203736 470836 203788
rect 471336 203736 471388 203788
rect 474372 203736 474424 203788
rect 474464 203736 474516 203788
rect 475844 203736 475896 203788
rect 463516 203668 463568 203720
rect 470508 203668 470560 203720
rect 456708 203600 456760 203652
rect 464712 203600 464764 203652
rect 473912 203668 473964 203720
rect 474004 203668 474056 203720
rect 478880 203668 478932 203720
rect 470784 203600 470836 203652
rect 480628 203600 480680 203652
rect 456064 203532 456116 203584
rect 465908 203532 465960 203584
rect 467288 203532 467340 203584
rect 335084 203464 335136 203516
rect 346400 203464 346452 203516
rect 369860 203464 369912 203516
rect 376300 203464 376352 203516
rect 461492 203464 461544 203516
rect 470416 203532 470468 203584
rect 470692 203532 470744 203584
rect 475568 203532 475620 203584
rect 475752 203532 475804 203584
rect 484400 203532 484452 203584
rect 329748 203396 329800 203448
rect 328276 203328 328328 203380
rect 335820 203328 335872 203380
rect 336004 203396 336056 203448
rect 343640 203396 343692 203448
rect 344192 203396 344244 203448
rect 347044 203396 347096 203448
rect 356428 203396 356480 203448
rect 447140 203396 447192 203448
rect 463056 203396 463108 203448
rect 472900 203464 472952 203516
rect 471796 203396 471848 203448
rect 339224 203328 339276 203380
rect 342720 203328 342772 203380
rect 332416 203260 332468 203312
rect 341340 203260 341392 203312
rect 342904 203260 342956 203312
rect 349160 203260 349212 203312
rect 460664 203328 460716 203380
rect 467564 203328 467616 203380
rect 351184 203260 351236 203312
rect 366364 203260 366416 203312
rect 368480 203260 368532 203312
rect 457904 203260 457956 203312
rect 467196 203260 467248 203312
rect 467748 203260 467800 203312
rect 474188 203260 474240 203312
rect 474372 203328 474424 203380
rect 478972 203328 479024 203380
rect 481640 203396 481692 203448
rect 480536 203328 480588 203380
rect 476120 203260 476172 203312
rect 331220 203192 331272 203244
rect 336556 203192 336608 203244
rect 345940 203192 345992 203244
rect 355600 203192 355652 203244
rect 459100 203192 459152 203244
rect 468484 203192 468536 203244
rect 477500 203192 477552 203244
rect 340604 203124 340656 203176
rect 340788 203124 340840 203176
rect 344192 203124 344244 203176
rect 344284 203124 344336 203176
rect 351092 203124 351144 203176
rect 351184 203124 351236 203176
rect 360016 203124 360068 203176
rect 453304 203124 453356 203176
rect 462412 203124 462464 203176
rect 471060 203124 471112 203176
rect 471152 203124 471204 203176
rect 481640 203124 481692 203176
rect 335268 203056 335320 203108
rect 342812 203056 342864 203108
rect 342904 203056 342956 203108
rect 344928 203056 344980 203108
rect 354588 203056 354640 203108
rect 451004 203056 451056 203108
rect 513380 203056 513432 203108
rect 296628 202988 296680 203040
rect 357440 202988 357492 203040
rect 453948 202988 454000 203040
rect 509240 202988 509292 203040
rect 336648 202920 336700 202972
rect 342904 202920 342956 202972
rect 342996 202920 343048 202972
rect 353300 202920 353352 202972
rect 455328 202920 455380 202972
rect 505100 202920 505152 202972
rect 295248 202852 295300 202904
rect 358820 202852 358872 202904
rect 454684 202852 454736 202904
rect 463056 202852 463108 202904
rect 469496 202852 469548 202904
rect 477500 202852 477552 202904
rect 297364 202784 297416 202836
rect 297916 202784 297968 202836
rect 408500 201560 408552 201612
rect 409144 201560 409196 201612
rect 500316 201560 500368 201612
rect 297916 201492 297968 201544
rect 417424 201492 417476 201544
rect 451924 201424 451976 201476
rect 499672 201424 499724 201476
rect 387708 201356 387760 201408
rect 500224 201356 500276 201408
rect 384948 201288 385000 201340
rect 499856 201288 499908 201340
rect 383568 201220 383620 201272
rect 499764 201220 499816 201272
rect 380808 201152 380860 201204
rect 499948 201152 500000 201204
rect 378048 201084 378100 201136
rect 500040 201084 500092 201136
rect 376668 201016 376720 201068
rect 500132 201016 500184 201068
rect 2964 200948 3016 201000
rect 521844 200948 521896 201000
rect 3792 200880 3844 200932
rect 521752 200880 521804 200932
rect 3608 200812 3660 200864
rect 521660 200812 521712 200864
rect 3884 200744 3936 200796
rect 521936 200744 521988 200796
rect 379796 183472 379848 183524
rect 409144 183472 409196 183524
rect 523868 182112 523920 182164
rect 580172 182112 580224 182164
rect 522764 171028 522816 171080
rect 580172 171028 580224 171080
rect 523776 158652 523828 158704
rect 579804 158652 579856 158704
rect 522672 135192 522724 135244
rect 580172 135192 580224 135244
rect 379980 124108 380032 124160
rect 391204 124108 391256 124160
rect 522580 124108 522632 124160
rect 580172 124108 580224 124160
rect 380072 118600 380124 118652
rect 393964 118600 394016 118652
rect 379980 115880 380032 115932
rect 395344 115880 395396 115932
rect 523684 111732 523736 111784
rect 579804 111732 579856 111784
rect 300768 110916 300820 110968
rect 416780 110916 416832 110968
rect 297916 108944 297968 108996
rect 303620 108944 303672 108996
rect 305644 108944 305696 108996
rect 307760 108944 307812 108996
rect 418068 108944 418120 108996
rect 424232 108944 424284 108996
rect 427820 108944 427872 108996
rect 531964 88272 532016 88324
rect 580172 88272 580224 88324
rect 522488 77188 522540 77240
rect 580172 77188 580224 77240
rect 527824 64812 527876 64864
rect 579804 64812 579856 64864
rect 529204 41352 529256 41404
rect 580172 41352 580224 41404
rect 522304 30268 522356 30320
rect 580172 30268 580224 30320
rect 525064 17892 525116 17944
rect 579804 17892 579856 17944
rect 3424 8236 3476 8288
rect 522120 8236 522172 8288
rect 7656 3544 7708 3596
rect 8208 3544 8260 3596
rect 8852 3544 8904 3596
rect 9588 3544 9640 3596
rect 10048 3544 10100 3596
rect 10968 3544 11020 3596
rect 11244 3544 11296 3596
rect 12348 3544 12400 3596
rect 12440 3544 12492 3596
rect 13636 3544 13688 3596
rect 16028 3544 16080 3596
rect 16488 3544 16540 3596
rect 17224 3544 17276 3596
rect 17868 3544 17920 3596
rect 18328 3544 18380 3596
rect 19248 3544 19300 3596
rect 19524 3544 19576 3596
rect 20628 3544 20680 3596
rect 20720 3544 20772 3596
rect 21916 3544 21968 3596
rect 24308 3544 24360 3596
rect 24768 3544 24820 3596
rect 25504 3544 25556 3596
rect 26148 3544 26200 3596
rect 26700 3544 26752 3596
rect 27528 3544 27580 3596
rect 27896 3544 27948 3596
rect 28908 3544 28960 3596
rect 29092 3544 29144 3596
rect 30196 3544 30248 3596
rect 33876 3544 33928 3596
rect 34428 3544 34480 3596
rect 34980 3544 35032 3596
rect 35808 3544 35860 3596
rect 36176 3544 36228 3596
rect 37188 3544 37240 3596
rect 37372 3544 37424 3596
rect 38476 3544 38528 3596
rect 42156 3544 42208 3596
rect 42708 3544 42760 3596
rect 43352 3544 43404 3596
rect 44088 3544 44140 3596
rect 44548 3544 44600 3596
rect 45468 3544 45520 3596
rect 45744 3544 45796 3596
rect 46848 3544 46900 3596
rect 46940 3544 46992 3596
rect 48136 3544 48188 3596
rect 50528 3544 50580 3596
rect 50988 3544 51040 3596
rect 51632 3544 51684 3596
rect 52368 3544 52420 3596
rect 52828 3544 52880 3596
rect 53748 3544 53800 3596
rect 54024 3544 54076 3596
rect 55128 3544 55180 3596
rect 55220 3544 55272 3596
rect 56416 3544 56468 3596
rect 58808 3544 58860 3596
rect 59268 3544 59320 3596
rect 60004 3544 60056 3596
rect 60648 3544 60700 3596
rect 61200 3544 61252 3596
rect 62028 3544 62080 3596
rect 63592 3544 63644 3596
rect 64696 3544 64748 3596
rect 68284 3544 68336 3596
rect 68928 3544 68980 3596
rect 69480 3544 69532 3596
rect 70308 3544 70360 3596
rect 70676 3544 70728 3596
rect 71688 3544 71740 3596
rect 71872 3544 71924 3596
rect 72976 3544 73028 3596
rect 76656 3544 76708 3596
rect 77208 3544 77260 3596
rect 77852 3544 77904 3596
rect 78588 3544 78640 3596
rect 79048 3544 79100 3596
rect 79968 3544 80020 3596
rect 80244 3544 80296 3596
rect 81348 3544 81400 3596
rect 81440 3544 81492 3596
rect 82636 3544 82688 3596
rect 84936 3544 84988 3596
rect 85488 3544 85540 3596
rect 86132 3544 86184 3596
rect 86868 3544 86920 3596
rect 87328 3544 87380 3596
rect 88248 3544 88300 3596
rect 88524 3544 88576 3596
rect 89628 3544 89680 3596
rect 89720 3544 89772 3596
rect 90916 3544 90968 3596
rect 93308 3544 93360 3596
rect 93768 3544 93820 3596
rect 94504 3544 94556 3596
rect 95148 3544 95200 3596
rect 95700 3544 95752 3596
rect 96528 3544 96580 3596
rect 96896 3544 96948 3596
rect 97908 3544 97960 3596
rect 98092 3544 98144 3596
rect 99196 3544 99248 3596
rect 102784 3544 102836 3596
rect 103428 3544 103480 3596
rect 103980 3544 104032 3596
rect 104808 3544 104860 3596
rect 105176 3544 105228 3596
rect 106188 3544 106240 3596
rect 106372 3544 106424 3596
rect 107476 3544 107528 3596
rect 111156 3544 111208 3596
rect 111708 3544 111760 3596
rect 112352 3544 112404 3596
rect 113088 3544 113140 3596
rect 113548 3544 113600 3596
rect 114468 3544 114520 3596
rect 114744 3544 114796 3596
rect 115848 3544 115900 3596
rect 115940 3544 115992 3596
rect 117136 3544 117188 3596
rect 119436 3544 119488 3596
rect 119988 3544 120040 3596
rect 120632 3544 120684 3596
rect 121368 3544 121420 3596
rect 121828 3544 121880 3596
rect 122748 3544 122800 3596
rect 123024 3544 123076 3596
rect 124128 3544 124180 3596
rect 124220 3544 124272 3596
rect 125416 3544 125468 3596
rect 127808 3544 127860 3596
rect 128268 3544 128320 3596
rect 129004 3544 129056 3596
rect 129648 3544 129700 3596
rect 130200 3544 130252 3596
rect 131028 3544 131080 3596
rect 131396 3544 131448 3596
rect 132408 3544 132460 3596
rect 132592 3544 132644 3596
rect 133788 3544 133840 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 2872 3476 2924 3528
rect 278136 3476 278188 3528
rect 4068 3408 4120 3460
rect 278044 3408 278096 3460
rect 101588 3272 101640 3324
rect 102048 3272 102100 3324
rect 62396 3136 62448 3188
rect 63408 3136 63460 3188
rect 142068 2796 142120 2848
rect 145656 2796 145708 2848
rect 149244 2796 149296 2848
rect 152740 2796 152792 2848
rect 156328 2796 156380 2848
rect 159916 2796 159968 2848
rect 163504 2796 163556 2848
rect 167092 2796 167144 2848
rect 170588 2796 170640 2848
rect 174176 2796 174228 2848
rect 177764 2796 177816 2848
rect 181352 2796 181404 2848
rect 184848 2796 184900 2848
rect 188436 2796 188488 2848
rect 192024 2796 192076 2848
rect 195612 2796 195664 2848
rect 199200 2796 199252 2848
rect 202696 2796 202748 2848
rect 206284 2796 206336 2848
rect 209872 2796 209924 2848
rect 213460 2796 213512 2848
rect 217048 2796 217100 2848
rect 220544 2796 220596 2848
rect 224132 2796 224184 2848
rect 227720 2796 227772 2848
rect 231308 2796 231360 2848
rect 234804 2796 234856 2848
rect 238392 2796 238444 2848
rect 241980 2796 242032 2848
rect 245568 2796 245620 2848
rect 249156 2796 249208 2848
rect 252652 2796 252704 2848
rect 256240 2796 256292 2848
rect 259828 2796 259880 2848
rect 263416 2796 263468 2848
rect 267004 2796 267056 2848
rect 270500 2796 270552 2848
rect 274088 2796 274140 2848
rect 277676 2796 277728 2848
rect 281264 2796 281316 2848
rect 284760 2796 284812 2848
rect 288348 2796 288400 2848
rect 291936 2796 291988 2848
rect 295524 2796 295576 2848
rect 299112 2796 299164 2848
rect 302608 2796 302660 2848
rect 305644 2796 305696 2848
rect 306196 2796 306248 2848
rect 309784 2796 309836 2848
rect 313372 2796 313424 2848
rect 316960 2796 317012 2848
rect 320456 2796 320508 2848
rect 324044 2796 324096 2848
rect 327632 2796 327684 2848
rect 331220 2796 331272 2848
rect 334716 2796 334768 2848
rect 338304 2796 338356 2848
rect 341892 2796 341944 2848
rect 345480 2796 345532 2848
rect 349068 2796 349120 2848
rect 352564 2796 352616 2848
rect 356152 2796 356204 2848
rect 359740 2796 359792 2848
rect 363328 2796 363380 2848
rect 366916 2796 366968 2848
rect 370412 2796 370464 2848
rect 374000 2796 374052 2848
rect 377588 2796 377640 2848
rect 381176 2796 381228 2848
rect 384672 2796 384724 2848
rect 388260 2796 388312 2848
rect 391848 2796 391900 2848
rect 395436 2796 395488 2848
rect 399024 2796 399076 2848
rect 402520 2796 402572 2848
rect 406108 2796 406160 2848
rect 409696 2796 409748 2848
rect 413284 2796 413336 2848
rect 416872 2796 416924 2848
rect 420368 2796 420420 2848
rect 423956 2796 424008 2848
rect 427544 2796 427596 2848
rect 431132 2796 431184 2848
rect 434628 2796 434680 2848
rect 438216 2796 438268 2848
rect 441804 2796 441856 2848
rect 445392 2796 445444 2848
rect 448980 2796 449032 2848
rect 452476 2796 452528 2848
rect 456064 2796 456116 2848
rect 459652 2796 459704 2848
rect 463240 2796 463292 2848
rect 466828 2796 466880 2848
rect 470324 2796 470376 2848
rect 473912 2796 473964 2848
rect 477500 2796 477552 2848
rect 481088 2796 481140 2848
rect 484584 2796 484636 2848
rect 488172 2796 488224 2848
rect 491760 2796 491812 2848
rect 495348 2796 495400 2848
rect 498936 2796 498988 2848
rect 502432 2796 502484 2848
rect 506020 2796 506072 2848
rect 509608 2796 509660 2848
rect 513196 2796 513248 2848
rect 516784 2796 516836 2848
rect 520280 2796 520332 2848
rect 523868 2796 523920 2848
rect 527456 2796 527508 2848
rect 531044 2796 531096 2848
rect 534540 2796 534592 2848
rect 538128 2796 538180 2848
rect 541716 2796 541768 2848
rect 545304 2796 545356 2848
rect 548892 2796 548944 2848
rect 552388 2796 552440 2848
rect 555976 2796 556028 2848
rect 559564 2796 559616 2848
rect 563152 2796 563204 2848
rect 566740 2796 566792 2848
rect 570236 2796 570288 2848
rect 573824 2796 573876 2848
rect 577412 2796 577464 2848
rect 581000 2796 581052 2848
rect 5264 552 5316 604
rect 5448 552 5500 604
rect 138480 552 138532 604
rect 142068 552 142120 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 24320 700505 24348 703520
rect 24306 700496 24362 700505
rect 24306 700431 24362 700440
rect 40512 700398 40540 703520
rect 72988 700641 73016 703520
rect 89180 700777 89208 703520
rect 89166 700768 89222 700777
rect 89166 700703 89222 700712
rect 72974 700632 73030 700641
rect 72974 700567 73030 700576
rect 40500 700392 40552 700398
rect 8114 700360 8170 700369
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 8114 700295 8170 700304
rect 3330 653576 3386 653585
rect 3330 653511 3386 653520
rect 3344 652905 3372 653511
rect 3330 652896 3386 652905
rect 3330 652831 3386 652840
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623801 3464 624815
rect 3422 623792 3478 623801
rect 3422 623727 3478 623736
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610366 3464 610399
rect 3424 610360 3476 610366
rect 3424 610302 3476 610308
rect 3514 596048 3570 596057
rect 3514 595983 3570 595992
rect 3330 509960 3386 509969
rect 3330 509895 3386 509904
rect 3344 509318 3372 509895
rect 3332 509312 3384 509318
rect 3332 509254 3384 509260
rect 3422 495544 3478 495553
rect 3422 495479 3424 495488
rect 3476 495479 3478 495488
rect 3424 495450 3476 495456
rect 2962 481128 3018 481137
rect 2962 481063 3018 481072
rect 2976 480282 3004 481063
rect 2964 480276 3016 480282
rect 2964 480218 3016 480224
rect 3424 478916 3476 478922
rect 3424 478858 3476 478864
rect 3240 425060 3292 425066
rect 3240 425002 3292 425008
rect 3252 423745 3280 425002
rect 3238 423736 3294 423745
rect 3238 423671 3294 423680
rect 3148 396024 3200 396030
rect 3148 395966 3200 395972
rect 3160 395049 3188 395966
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 3056 295316 3108 295322
rect 3056 295258 3108 295264
rect 3068 294409 3096 295258
rect 3054 294400 3110 294409
rect 3054 294335 3110 294344
rect 2688 242956 2740 242962
rect 2688 242898 2740 242904
rect 1308 240168 1360 240174
rect 1308 240110 1360 240116
rect 1320 3534 1348 240110
rect 2700 3534 2728 242898
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 2964 201000 3016 201006
rect 2964 200942 3016 200948
rect 2976 193905 3004 200942
rect 2962 193896 3018 193905
rect 2962 193831 3018 193840
rect 3330 50960 3386 50969
rect 3330 50895 3386 50904
rect 3344 50153 3372 50895
rect 3330 50144 3386 50153
rect 3330 50079 3386 50088
rect 3436 21457 3464 478858
rect 3528 478242 3556 595983
rect 3606 567352 3662 567361
rect 3606 567287 3662 567296
rect 3620 479534 3648 567287
rect 3698 553072 3754 553081
rect 3698 553007 3754 553016
rect 3608 479528 3660 479534
rect 3608 479470 3660 479476
rect 3516 478236 3568 478242
rect 3516 478178 3568 478184
rect 3712 478174 3740 553007
rect 3790 538656 3846 538665
rect 3790 538591 3846 538600
rect 3804 478310 3832 538591
rect 41340 479369 41368 700334
rect 105464 699718 105492 703520
rect 137848 700330 137876 703520
rect 154132 700398 154160 703520
rect 170324 700942 170352 703520
rect 170312 700936 170364 700942
rect 170312 700878 170364 700884
rect 171048 700936 171100 700942
rect 171048 700878 171100 700884
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 71318 479904 71374 479913
rect 71318 479839 71374 479848
rect 71332 479641 71360 479839
rect 61842 479632 61898 479641
rect 61842 479567 61898 479576
rect 71318 479632 71374 479641
rect 106200 479602 106228 699654
rect 171060 479670 171088 700878
rect 202800 700466 202828 703520
rect 218992 700534 219020 703520
rect 218980 700528 219032 700534
rect 218980 700470 219032 700476
rect 202788 700460 202840 700466
rect 202788 700402 202840 700408
rect 235184 699718 235212 703520
rect 267660 700602 267688 703520
rect 283852 700670 283880 703520
rect 283840 700664 283892 700670
rect 283840 700606 283892 700612
rect 267648 700596 267700 700602
rect 267648 700538 267700 700544
rect 300136 699718 300164 703520
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300584 699712 300636 699718
rect 300584 699654 300636 699660
rect 235920 479738 235948 699654
rect 298006 606656 298062 606665
rect 298006 606591 298062 606600
rect 297914 605432 297970 605441
rect 297914 605367 297970 605376
rect 297822 603800 297878 603809
rect 297822 603735 297878 603744
rect 297730 602576 297786 602585
rect 297730 602511 297786 602520
rect 297638 600944 297694 600953
rect 297638 600879 297694 600888
rect 297546 599856 297602 599865
rect 297546 599791 297602 599800
rect 297454 598088 297510 598097
rect 297454 598023 297510 598032
rect 297362 540288 297418 540297
rect 297362 540223 297418 540232
rect 297270 538520 297326 538529
rect 297270 538455 297326 538464
rect 297284 520946 297312 538455
rect 297272 520940 297324 520946
rect 297272 520882 297324 520888
rect 292488 518424 292540 518430
rect 292488 518366 292540 518372
rect 285588 517880 285640 517886
rect 285588 517822 285640 517828
rect 280896 517744 280948 517750
rect 280896 517686 280948 517692
rect 235908 479732 235960 479738
rect 235908 479674 235960 479680
rect 171048 479664 171100 479670
rect 108946 479632 109002 479641
rect 71318 479567 71374 479576
rect 106188 479596 106240 479602
rect 50986 479496 51042 479505
rect 50986 479431 50988 479440
rect 51040 479431 51042 479440
rect 57796 479460 57848 479466
rect 50988 479402 51040 479408
rect 57796 479402 57848 479408
rect 57808 479369 57836 479402
rect 41326 479360 41382 479369
rect 41326 479295 41382 479304
rect 57794 479360 57850 479369
rect 57794 479295 57850 479304
rect 57978 479360 58034 479369
rect 61856 479330 61884 479567
rect 109130 479632 109186 479641
rect 109002 479590 109130 479618
rect 108946 479567 109002 479576
rect 171048 479606 171100 479612
rect 109130 479567 109186 479576
rect 278792 479590 278912 479618
rect 106188 479538 106240 479544
rect 278792 479505 278820 479590
rect 99378 479496 99434 479505
rect 135166 479496 135222 479505
rect 99434 479454 99512 479482
rect 99378 479431 99434 479440
rect 57978 479295 57980 479304
rect 58032 479295 58034 479304
rect 61844 479324 61896 479330
rect 57980 479266 58032 479272
rect 61844 479266 61896 479272
rect 99484 479233 99512 479454
rect 128268 479460 128320 479466
rect 135166 479431 135168 479440
rect 128268 479402 128320 479408
rect 135220 479431 135222 479440
rect 154486 479496 154542 479505
rect 154486 479431 154542 479440
rect 173806 479496 173862 479505
rect 173806 479431 173862 479440
rect 193126 479496 193182 479505
rect 193126 479431 193182 479440
rect 212446 479496 212502 479505
rect 212446 479431 212502 479440
rect 231766 479496 231822 479505
rect 231766 479431 231822 479440
rect 251086 479496 251142 479505
rect 251086 479431 251142 479440
rect 278778 479496 278834 479505
rect 278884 479466 278912 479590
rect 278778 479431 278834 479440
rect 278872 479460 278924 479466
rect 135168 479402 135220 479408
rect 128280 479369 128308 479402
rect 154500 479398 154528 479431
rect 173820 479398 173848 479431
rect 193140 479398 193168 479431
rect 212460 479398 212488 479431
rect 231780 479398 231808 479431
rect 251100 479398 251128 479431
rect 278872 479402 278924 479408
rect 147588 479392 147640 479398
rect 128266 479360 128322 479369
rect 128266 479295 128322 479304
rect 147586 479360 147588 479369
rect 154488 479392 154540 479398
rect 147640 479360 147642 479369
rect 166908 479392 166960 479398
rect 154488 479334 154540 479340
rect 166906 479360 166908 479369
rect 173808 479392 173860 479398
rect 166960 479360 166962 479369
rect 147586 479295 147642 479304
rect 186228 479392 186280 479398
rect 173808 479334 173860 479340
rect 186226 479360 186228 479369
rect 193128 479392 193180 479398
rect 186280 479360 186282 479369
rect 166906 479295 166962 479304
rect 205548 479392 205600 479398
rect 193128 479334 193180 479340
rect 205546 479360 205548 479369
rect 212448 479392 212500 479398
rect 205600 479360 205602 479369
rect 186226 479295 186282 479304
rect 224868 479392 224920 479398
rect 212448 479334 212500 479340
rect 224866 479360 224868 479369
rect 231768 479392 231820 479398
rect 224920 479360 224922 479369
rect 205546 479295 205602 479304
rect 244188 479392 244240 479398
rect 231768 479334 231820 479340
rect 244186 479360 244188 479369
rect 251088 479392 251140 479398
rect 244240 479360 244242 479369
rect 224866 479295 224922 479304
rect 251088 479334 251140 479340
rect 244186 479295 244242 479304
rect 99470 479224 99526 479233
rect 99470 479159 99526 479168
rect 279700 479188 279752 479194
rect 279700 479130 279752 479136
rect 279608 479120 279660 479126
rect 279608 479062 279660 479068
rect 135168 478984 135220 478990
rect 277400 478984 277452 478990
rect 135168 478926 135220 478932
rect 277398 478952 277400 478961
rect 277452 478952 277454 478961
rect 3792 478304 3844 478310
rect 3792 478246 3844 478252
rect 3700 478168 3752 478174
rect 3700 478110 3752 478116
rect 133788 476128 133840 476134
rect 133788 476070 133840 476076
rect 132408 473408 132460 473414
rect 132408 473350 132460 473356
rect 131028 472048 131080 472054
rect 131028 471990 131080 471996
rect 129648 469260 129700 469266
rect 129648 469202 129700 469208
rect 128268 467900 128320 467906
rect 128268 467842 128320 467848
rect 126888 465112 126940 465118
rect 126888 465054 126940 465060
rect 125508 463752 125560 463758
rect 125508 463694 125560 463700
rect 125416 460964 125468 460970
rect 125416 460906 125468 460912
rect 124128 459604 124180 459610
rect 124128 459546 124180 459552
rect 122748 456816 122800 456822
rect 122748 456758 122800 456764
rect 121368 455456 121420 455462
rect 121368 455398 121420 455404
rect 119988 452668 120040 452674
rect 119988 452610 120040 452616
rect 3516 452600 3568 452606
rect 3516 452542 3568 452548
rect 3528 452441 3556 452542
rect 3514 452432 3570 452441
rect 3514 452367 3570 452376
rect 118608 451308 118660 451314
rect 118608 451250 118660 451256
rect 117228 448588 117280 448594
rect 117228 448530 117280 448536
rect 117136 445800 117188 445806
rect 117136 445742 117188 445748
rect 115848 444440 115900 444446
rect 115848 444382 115900 444388
rect 114468 441652 114520 441658
rect 114468 441594 114520 441600
rect 113088 440292 113140 440298
rect 113088 440234 113140 440240
rect 3516 438864 3568 438870
rect 3516 438806 3568 438812
rect 3528 438025 3556 438806
rect 3514 438016 3570 438025
rect 3514 437951 3570 437960
rect 111708 437504 111760 437510
rect 111708 437446 111760 437452
rect 110328 436144 110380 436150
rect 110328 436086 110380 436092
rect 108948 433356 109000 433362
rect 108948 433298 109000 433304
rect 107568 431996 107620 432002
rect 107568 431938 107620 431944
rect 107476 429208 107528 429214
rect 107476 429150 107528 429156
rect 106188 427848 106240 427854
rect 106188 427790 106240 427796
rect 104808 425128 104860 425134
rect 104808 425070 104860 425076
rect 103428 423700 103480 423706
rect 103428 423642 103480 423648
rect 102048 420980 102100 420986
rect 102048 420922 102100 420928
rect 100668 418192 100720 418198
rect 100668 418134 100720 418140
rect 99288 416832 99340 416838
rect 99288 416774 99340 416780
rect 99196 414044 99248 414050
rect 99196 413986 99248 413992
rect 97908 412684 97960 412690
rect 97908 412626 97960 412632
rect 96528 409896 96580 409902
rect 96528 409838 96580 409844
rect 95148 408536 95200 408542
rect 95148 408478 95200 408484
rect 93768 405748 93820 405754
rect 93768 405690 93820 405696
rect 92388 404388 92440 404394
rect 92388 404330 92440 404336
rect 91008 401668 91060 401674
rect 91008 401610 91060 401616
rect 90916 400240 90968 400246
rect 90916 400182 90968 400188
rect 89628 397520 89680 397526
rect 89628 397462 89680 397468
rect 88248 396092 88300 396098
rect 88248 396034 88300 396040
rect 86868 393372 86920 393378
rect 86868 393314 86920 393320
rect 85488 390584 85540 390590
rect 85488 390526 85540 390532
rect 84108 389224 84160 389230
rect 84108 389166 84160 389172
rect 82728 386436 82780 386442
rect 82728 386378 82780 386384
rect 82636 385076 82688 385082
rect 82636 385018 82688 385024
rect 81348 382288 81400 382294
rect 81348 382230 81400 382236
rect 79968 380928 80020 380934
rect 79968 380870 80020 380876
rect 3516 380860 3568 380866
rect 3516 380802 3568 380808
rect 3528 380633 3556 380802
rect 3514 380624 3570 380633
rect 3514 380559 3570 380568
rect 78588 378208 78640 378214
rect 78588 378150 78640 378156
rect 77208 376780 77260 376786
rect 77208 376722 77260 376728
rect 75828 374060 75880 374066
rect 75828 374002 75880 374008
rect 74448 372632 74500 372638
rect 74448 372574 74500 372580
rect 73068 369912 73120 369918
rect 73068 369854 73120 369860
rect 72976 368552 73028 368558
rect 72976 368494 73028 368500
rect 3516 367056 3568 367062
rect 3516 366998 3568 367004
rect 3528 366217 3556 366998
rect 3514 366208 3570 366217
rect 3514 366143 3570 366152
rect 71688 365764 71740 365770
rect 71688 365706 71740 365712
rect 70308 362976 70360 362982
rect 70308 362918 70360 362924
rect 68928 361616 68980 361622
rect 68928 361558 68980 361564
rect 67548 358828 67600 358834
rect 67548 358770 67600 358776
rect 66168 357468 66220 357474
rect 66168 357410 66220 357416
rect 64788 354748 64840 354754
rect 64788 354690 64840 354696
rect 64696 353320 64748 353326
rect 64696 353262 64748 353268
rect 63408 350600 63460 350606
rect 63408 350542 63460 350548
rect 62028 349172 62080 349178
rect 62028 349114 62080 349120
rect 60648 346452 60700 346458
rect 60648 346394 60700 346400
rect 59268 345092 59320 345098
rect 59268 345034 59320 345040
rect 57888 342304 57940 342310
rect 57888 342246 57940 342252
rect 56508 340944 56560 340950
rect 56508 340886 56560 340892
rect 56416 338156 56468 338162
rect 56416 338098 56468 338104
rect 3516 338088 3568 338094
rect 3516 338030 3568 338036
rect 3528 337521 3556 338030
rect 3514 337512 3570 337521
rect 3514 337447 3570 337456
rect 55128 335368 55180 335374
rect 55128 335310 55180 335316
rect 53748 334008 53800 334014
rect 53748 333950 53800 333956
rect 52368 331288 52420 331294
rect 52368 331230 52420 331236
rect 50988 329860 51040 329866
rect 50988 329802 51040 329808
rect 49608 327140 49660 327146
rect 49608 327082 49660 327088
rect 48228 325712 48280 325718
rect 48228 325654 48280 325660
rect 3516 324284 3568 324290
rect 3516 324226 3568 324232
rect 3528 323105 3556 324226
rect 3514 323096 3570 323105
rect 3514 323031 3570 323040
rect 48136 322992 48188 322998
rect 48136 322934 48188 322940
rect 46848 321632 46900 321638
rect 46848 321574 46900 321580
rect 45468 318844 45520 318850
rect 45468 318786 45520 318792
rect 44088 317484 44140 317490
rect 44088 317426 44140 317432
rect 42708 314696 42760 314702
rect 42708 314638 42760 314644
rect 41328 313336 41380 313342
rect 41328 313278 41380 313284
rect 39948 310548 40000 310554
rect 39948 310490 40000 310496
rect 38568 307828 38620 307834
rect 38568 307770 38620 307776
rect 38476 306400 38528 306406
rect 38476 306342 38528 306348
rect 37188 303680 37240 303686
rect 37188 303622 37240 303628
rect 35808 302252 35860 302258
rect 35808 302194 35860 302200
rect 34428 299532 34480 299538
rect 34428 299474 34480 299480
rect 33048 298172 33100 298178
rect 33048 298114 33100 298120
rect 31668 295384 31720 295390
rect 31668 295326 31720 295332
rect 30288 294024 30340 294030
rect 30288 293966 30340 293972
rect 30196 291236 30248 291242
rect 30196 291178 30248 291184
rect 28908 289876 28960 289882
rect 28908 289818 28960 289824
rect 27528 287088 27580 287094
rect 27528 287030 27580 287036
rect 26148 285728 26200 285734
rect 26148 285670 26200 285676
rect 24768 282940 24820 282946
rect 24768 282882 24820 282888
rect 23388 280220 23440 280226
rect 23388 280162 23440 280168
rect 3516 280152 3568 280158
rect 3514 280120 3516 280129
rect 3568 280120 3570 280129
rect 3514 280055 3570 280064
rect 22008 278792 22060 278798
rect 22008 278734 22060 278740
rect 21916 276072 21968 276078
rect 21916 276014 21968 276020
rect 20628 274712 20680 274718
rect 20628 274654 20680 274660
rect 19248 271924 19300 271930
rect 19248 271866 19300 271872
rect 17868 270564 17920 270570
rect 17868 270506 17920 270512
rect 16488 267776 16540 267782
rect 16488 267718 16540 267724
rect 15108 266416 15160 266422
rect 15108 266358 15160 266364
rect 3514 265704 3570 265713
rect 3514 265639 3570 265648
rect 3528 240922 3556 265639
rect 13728 263628 13780 263634
rect 13728 263570 13780 263576
rect 13636 262268 13688 262274
rect 13636 262210 13688 262216
rect 12348 259480 12400 259486
rect 12348 259422 12400 259428
rect 10968 256760 11020 256766
rect 10968 256702 11020 256708
rect 9588 255332 9640 255338
rect 9588 255274 9640 255280
rect 8208 252612 8260 252618
rect 8208 252554 8260 252560
rect 3606 251288 3662 251297
rect 3606 251223 3662 251232
rect 6828 251252 6880 251258
rect 3516 240916 3568 240922
rect 3516 240858 3568 240864
rect 3620 240854 3648 251223
rect 6828 251194 6880 251200
rect 5448 248464 5500 248470
rect 5448 248406 5500 248412
rect 3608 240848 3660 240854
rect 3608 240790 3660 240796
rect 3516 237380 3568 237386
rect 3516 237322 3568 237328
rect 3528 237017 3556 237322
rect 3514 237008 3570 237017
rect 3514 236943 3570 236952
rect 3516 208344 3568 208350
rect 3516 208286 3568 208292
rect 3528 208185 3556 208286
rect 3514 208176 3570 208185
rect 3514 208111 3570 208120
rect 3792 200932 3844 200938
rect 3792 200874 3844 200880
rect 3608 200864 3660 200870
rect 3608 200806 3660 200812
rect 3698 200832 3754 200841
rect 3514 200696 3570 200705
rect 3514 200631 3570 200640
rect 3528 122097 3556 200631
rect 3620 150793 3648 200806
rect 3698 200767 3754 200776
rect 3606 150784 3662 150793
rect 3606 150719 3662 150728
rect 3712 136377 3740 200767
rect 3804 165073 3832 200874
rect 3884 200796 3936 200802
rect 3884 200738 3936 200744
rect 3896 179489 3924 200738
rect 3882 179480 3938 179489
rect 3882 179415 3938 179424
rect 3790 165064 3846 165073
rect 3790 164999 3846 165008
rect 3698 136368 3754 136377
rect 3698 136303 3754 136312
rect 3514 122088 3570 122097
rect 3514 122023 3570 122032
rect 3514 108896 3570 108905
rect 3514 108831 3570 108840
rect 3528 107681 3556 108831
rect 3514 107672 3570 107681
rect 3514 107607 3570 107616
rect 3514 80064 3570 80073
rect 3514 79999 3570 80008
rect 3528 78985 3556 79999
rect 3514 78976 3570 78985
rect 3514 78911 3570 78920
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 584 480 612 3470
rect 1688 480 1716 3470
rect 2884 480 2912 3470
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 5460 610 5488 248406
rect 6840 626 6868 251194
rect 8220 3602 8248 252554
rect 9600 3602 9628 255274
rect 10980 3602 11008 256702
rect 12360 3602 12388 259422
rect 13648 3602 13676 262210
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5448 604 5500 610
rect 5448 546 5500 552
rect 6472 598 6868 626
rect 5276 480 5304 546
rect 6472 480 6500 598
rect 7668 480 7696 3538
rect 8864 480 8892 3538
rect 10060 480 10088 3538
rect 11256 480 11284 3538
rect 12452 480 12480 3538
rect 13740 3482 13768 263570
rect 15120 3482 15148 266358
rect 16500 3602 16528 267718
rect 17880 3602 17908 270506
rect 19260 3602 19288 271866
rect 20640 3602 20668 274654
rect 21928 3602 21956 276014
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 13648 3454 13768 3482
rect 14844 3454 15148 3482
rect 13648 480 13676 3454
rect 14844 480 14872 3454
rect 16040 480 16068 3538
rect 17236 480 17264 3538
rect 18340 480 18368 3538
rect 19536 480 19564 3538
rect 20732 480 20760 3538
rect 22020 3482 22048 278734
rect 23400 3482 23428 280162
rect 24780 3602 24808 282882
rect 26160 3602 26188 285670
rect 27540 3602 27568 287030
rect 28920 3602 28948 289818
rect 30208 3602 30236 291178
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26700 3596 26752 3602
rect 26700 3538 26752 3544
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27896 3596 27948 3602
rect 27896 3538 27948 3544
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 21928 3454 22048 3482
rect 23124 3454 23428 3482
rect 21928 480 21956 3454
rect 23124 480 23152 3454
rect 24320 480 24348 3538
rect 25516 480 25544 3538
rect 26712 480 26740 3538
rect 27908 480 27936 3538
rect 29104 480 29132 3538
rect 30300 480 30328 293966
rect 31680 3482 31708 295326
rect 33060 3482 33088 298114
rect 34440 3602 34468 299474
rect 35820 3602 35848 302194
rect 37200 3602 37228 303622
rect 38488 3602 38516 306342
rect 33876 3596 33928 3602
rect 33876 3538 33928 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34980 3596 35032 3602
rect 34980 3538 35032 3544
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 36176 3596 36228 3602
rect 36176 3538 36228 3544
rect 37188 3596 37240 3602
rect 37188 3538 37240 3544
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 38476 3596 38528 3602
rect 38476 3538 38528 3544
rect 31496 3454 31708 3482
rect 32692 3454 33088 3482
rect 31496 480 31524 3454
rect 32692 480 32720 3454
rect 33888 480 33916 3538
rect 34992 480 35020 3538
rect 36188 480 36216 3538
rect 37384 480 37412 3538
rect 38580 480 38608 307770
rect 39960 3482 39988 310490
rect 41340 3482 41368 313278
rect 42720 3602 42748 314638
rect 44100 3602 44128 317426
rect 45480 3602 45508 318786
rect 46860 3602 46888 321574
rect 48148 3602 48176 322934
rect 42156 3596 42208 3602
rect 42156 3538 42208 3544
rect 42708 3596 42760 3602
rect 42708 3538 42760 3544
rect 43352 3596 43404 3602
rect 43352 3538 43404 3544
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 44548 3596 44600 3602
rect 44548 3538 44600 3544
rect 45468 3596 45520 3602
rect 45468 3538 45520 3544
rect 45744 3596 45796 3602
rect 45744 3538 45796 3544
rect 46848 3596 46900 3602
rect 46848 3538 46900 3544
rect 46940 3596 46992 3602
rect 46940 3538 46992 3544
rect 48136 3596 48188 3602
rect 48136 3538 48188 3544
rect 39776 3454 39988 3482
rect 40972 3454 41368 3482
rect 39776 480 39804 3454
rect 40972 480 41000 3454
rect 42168 480 42196 3538
rect 43364 480 43392 3538
rect 44560 480 44588 3538
rect 45756 480 45784 3538
rect 46952 480 46980 3538
rect 48240 3482 48268 325654
rect 49620 3482 49648 327082
rect 51000 3602 51028 329802
rect 52380 3602 52408 331230
rect 53760 3602 53788 333950
rect 55140 3602 55168 335310
rect 56428 3602 56456 338098
rect 50528 3596 50580 3602
rect 50528 3538 50580 3544
rect 50988 3596 51040 3602
rect 50988 3538 51040 3544
rect 51632 3596 51684 3602
rect 51632 3538 51684 3544
rect 52368 3596 52420 3602
rect 52368 3538 52420 3544
rect 52828 3596 52880 3602
rect 52828 3538 52880 3544
rect 53748 3596 53800 3602
rect 53748 3538 53800 3544
rect 54024 3596 54076 3602
rect 54024 3538 54076 3544
rect 55128 3596 55180 3602
rect 55128 3538 55180 3544
rect 55220 3596 55272 3602
rect 55220 3538 55272 3544
rect 56416 3596 56468 3602
rect 56416 3538 56468 3544
rect 48148 3454 48268 3482
rect 49344 3454 49648 3482
rect 48148 480 48176 3454
rect 49344 480 49372 3454
rect 50540 480 50568 3538
rect 51644 480 51672 3538
rect 52840 480 52868 3538
rect 54036 480 54064 3538
rect 55232 480 55260 3538
rect 56520 3482 56548 340886
rect 57900 3482 57928 342246
rect 59280 3602 59308 345034
rect 60660 3602 60688 346394
rect 62040 3602 62068 349114
rect 58808 3596 58860 3602
rect 58808 3538 58860 3544
rect 59268 3596 59320 3602
rect 59268 3538 59320 3544
rect 60004 3596 60056 3602
rect 60004 3538 60056 3544
rect 60648 3596 60700 3602
rect 60648 3538 60700 3544
rect 61200 3596 61252 3602
rect 61200 3538 61252 3544
rect 62028 3596 62080 3602
rect 62028 3538 62080 3544
rect 56428 3454 56548 3482
rect 57624 3454 57928 3482
rect 56428 480 56456 3454
rect 57624 480 57652 3454
rect 58820 480 58848 3538
rect 60016 480 60044 3538
rect 61212 480 61240 3538
rect 63420 3194 63448 350542
rect 64708 3602 64736 353262
rect 63592 3596 63644 3602
rect 63592 3538 63644 3544
rect 64696 3596 64748 3602
rect 64696 3538 64748 3544
rect 62396 3188 62448 3194
rect 62396 3130 62448 3136
rect 63408 3188 63460 3194
rect 63408 3130 63460 3136
rect 62408 480 62436 3130
rect 63604 480 63632 3538
rect 64800 480 64828 354690
rect 66180 3482 66208 357410
rect 67560 3482 67588 358770
rect 68940 3602 68968 361558
rect 70320 3602 70348 362918
rect 71700 3602 71728 365706
rect 72988 3602 73016 368494
rect 68284 3596 68336 3602
rect 68284 3538 68336 3544
rect 68928 3596 68980 3602
rect 68928 3538 68980 3544
rect 69480 3596 69532 3602
rect 69480 3538 69532 3544
rect 70308 3596 70360 3602
rect 70308 3538 70360 3544
rect 70676 3596 70728 3602
rect 70676 3538 70728 3544
rect 71688 3596 71740 3602
rect 71688 3538 71740 3544
rect 71872 3596 71924 3602
rect 71872 3538 71924 3544
rect 72976 3596 73028 3602
rect 72976 3538 73028 3544
rect 65996 3454 66208 3482
rect 67192 3454 67588 3482
rect 65996 480 66024 3454
rect 67192 480 67220 3454
rect 68296 480 68324 3538
rect 69492 480 69520 3538
rect 70688 480 70716 3538
rect 71884 480 71912 3538
rect 73080 480 73108 369854
rect 74460 3482 74488 372574
rect 75840 3482 75868 374002
rect 77220 3602 77248 376722
rect 78600 3602 78628 378150
rect 79980 3602 80008 380870
rect 81360 3602 81388 382230
rect 82648 3602 82676 385018
rect 76656 3596 76708 3602
rect 76656 3538 76708 3544
rect 77208 3596 77260 3602
rect 77208 3538 77260 3544
rect 77852 3596 77904 3602
rect 77852 3538 77904 3544
rect 78588 3596 78640 3602
rect 78588 3538 78640 3544
rect 79048 3596 79100 3602
rect 79048 3538 79100 3544
rect 79968 3596 80020 3602
rect 79968 3538 80020 3544
rect 80244 3596 80296 3602
rect 80244 3538 80296 3544
rect 81348 3596 81400 3602
rect 81348 3538 81400 3544
rect 81440 3596 81492 3602
rect 81440 3538 81492 3544
rect 82636 3596 82688 3602
rect 82636 3538 82688 3544
rect 74276 3454 74488 3482
rect 75472 3454 75868 3482
rect 74276 480 74304 3454
rect 75472 480 75500 3454
rect 76668 480 76696 3538
rect 77864 480 77892 3538
rect 79060 480 79088 3538
rect 80256 480 80284 3538
rect 81452 480 81480 3538
rect 82740 3482 82768 386378
rect 84120 3482 84148 389166
rect 85500 3602 85528 390526
rect 86880 3602 86908 393314
rect 88260 3602 88288 396034
rect 89640 3602 89668 397462
rect 90928 3602 90956 400182
rect 84936 3596 84988 3602
rect 84936 3538 84988 3544
rect 85488 3596 85540 3602
rect 85488 3538 85540 3544
rect 86132 3596 86184 3602
rect 86132 3538 86184 3544
rect 86868 3596 86920 3602
rect 86868 3538 86920 3544
rect 87328 3596 87380 3602
rect 87328 3538 87380 3544
rect 88248 3596 88300 3602
rect 88248 3538 88300 3544
rect 88524 3596 88576 3602
rect 88524 3538 88576 3544
rect 89628 3596 89680 3602
rect 89628 3538 89680 3544
rect 89720 3596 89772 3602
rect 89720 3538 89772 3544
rect 90916 3596 90968 3602
rect 90916 3538 90968 3544
rect 82648 3454 82768 3482
rect 83844 3454 84148 3482
rect 82648 480 82676 3454
rect 83844 480 83872 3454
rect 84948 480 84976 3538
rect 86144 480 86172 3538
rect 87340 480 87368 3538
rect 88536 480 88564 3538
rect 89732 480 89760 3538
rect 91020 3482 91048 401610
rect 92400 3482 92428 404330
rect 93780 3602 93808 405690
rect 95160 3602 95188 408478
rect 96540 3602 96568 409838
rect 97920 3602 97948 412626
rect 99208 3602 99236 413986
rect 93308 3596 93360 3602
rect 93308 3538 93360 3544
rect 93768 3596 93820 3602
rect 93768 3538 93820 3544
rect 94504 3596 94556 3602
rect 94504 3538 94556 3544
rect 95148 3596 95200 3602
rect 95148 3538 95200 3544
rect 95700 3596 95752 3602
rect 95700 3538 95752 3544
rect 96528 3596 96580 3602
rect 96528 3538 96580 3544
rect 96896 3596 96948 3602
rect 96896 3538 96948 3544
rect 97908 3596 97960 3602
rect 97908 3538 97960 3544
rect 98092 3596 98144 3602
rect 98092 3538 98144 3544
rect 99196 3596 99248 3602
rect 99196 3538 99248 3544
rect 90928 3454 91048 3482
rect 92124 3454 92428 3482
rect 90928 480 90956 3454
rect 92124 480 92152 3454
rect 93320 480 93348 3538
rect 94516 480 94544 3538
rect 95712 480 95740 3538
rect 96908 480 96936 3538
rect 98104 480 98132 3538
rect 99300 480 99328 416774
rect 100680 3482 100708 418134
rect 100496 3454 100708 3482
rect 100496 480 100524 3454
rect 102060 3330 102088 420922
rect 103440 3602 103468 423642
rect 104820 3602 104848 425070
rect 106200 3602 106228 427790
rect 107488 3602 107516 429150
rect 102784 3596 102836 3602
rect 102784 3538 102836 3544
rect 103428 3596 103480 3602
rect 103428 3538 103480 3544
rect 103980 3596 104032 3602
rect 103980 3538 104032 3544
rect 104808 3596 104860 3602
rect 104808 3538 104860 3544
rect 105176 3596 105228 3602
rect 105176 3538 105228 3544
rect 106188 3596 106240 3602
rect 106188 3538 106240 3544
rect 106372 3596 106424 3602
rect 106372 3538 106424 3544
rect 107476 3596 107528 3602
rect 107476 3538 107528 3544
rect 101588 3324 101640 3330
rect 101588 3266 101640 3272
rect 102048 3324 102100 3330
rect 102048 3266 102100 3272
rect 101600 480 101628 3266
rect 102796 480 102824 3538
rect 103992 480 104020 3538
rect 105188 480 105216 3538
rect 106384 480 106412 3538
rect 107580 480 107608 431938
rect 108960 3482 108988 433298
rect 110340 3482 110368 436086
rect 111720 3602 111748 437446
rect 113100 3602 113128 440234
rect 114480 3602 114508 441594
rect 115860 3602 115888 444382
rect 117148 3602 117176 445742
rect 111156 3596 111208 3602
rect 111156 3538 111208 3544
rect 111708 3596 111760 3602
rect 111708 3538 111760 3544
rect 112352 3596 112404 3602
rect 112352 3538 112404 3544
rect 113088 3596 113140 3602
rect 113088 3538 113140 3544
rect 113548 3596 113600 3602
rect 113548 3538 113600 3544
rect 114468 3596 114520 3602
rect 114468 3538 114520 3544
rect 114744 3596 114796 3602
rect 114744 3538 114796 3544
rect 115848 3596 115900 3602
rect 115848 3538 115900 3544
rect 115940 3596 115992 3602
rect 115940 3538 115992 3544
rect 117136 3596 117188 3602
rect 117136 3538 117188 3544
rect 108776 3454 108988 3482
rect 109972 3454 110368 3482
rect 108776 480 108804 3454
rect 109972 480 110000 3454
rect 111168 480 111196 3538
rect 112364 480 112392 3538
rect 113560 480 113588 3538
rect 114756 480 114784 3538
rect 115952 480 115980 3538
rect 117240 3482 117268 448530
rect 118620 3482 118648 451250
rect 120000 3602 120028 452610
rect 121380 3602 121408 455398
rect 122760 3602 122788 456758
rect 124140 3602 124168 459546
rect 125428 3602 125456 460906
rect 119436 3596 119488 3602
rect 119436 3538 119488 3544
rect 119988 3596 120040 3602
rect 119988 3538 120040 3544
rect 120632 3596 120684 3602
rect 120632 3538 120684 3544
rect 121368 3596 121420 3602
rect 121368 3538 121420 3544
rect 121828 3596 121880 3602
rect 121828 3538 121880 3544
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 123024 3596 123076 3602
rect 123024 3538 123076 3544
rect 124128 3596 124180 3602
rect 124128 3538 124180 3544
rect 124220 3596 124272 3602
rect 124220 3538 124272 3544
rect 125416 3596 125468 3602
rect 125416 3538 125468 3544
rect 117148 3454 117268 3482
rect 118252 3454 118648 3482
rect 117148 480 117176 3454
rect 118252 480 118280 3454
rect 119448 480 119476 3538
rect 120644 480 120672 3538
rect 121840 480 121868 3538
rect 123036 480 123064 3538
rect 124232 480 124260 3538
rect 125520 3482 125548 463694
rect 126900 3482 126928 465054
rect 128280 3602 128308 467842
rect 129660 3602 129688 469202
rect 131040 3602 131068 471990
rect 132420 3602 132448 473350
rect 133800 3602 133828 476070
rect 127808 3596 127860 3602
rect 127808 3538 127860 3544
rect 128268 3596 128320 3602
rect 128268 3538 128320 3544
rect 129004 3596 129056 3602
rect 129004 3538 129056 3544
rect 129648 3596 129700 3602
rect 129648 3538 129700 3544
rect 130200 3596 130252 3602
rect 130200 3538 130252 3544
rect 131028 3596 131080 3602
rect 131028 3538 131080 3544
rect 131396 3596 131448 3602
rect 131396 3538 131448 3544
rect 132408 3596 132460 3602
rect 132408 3538 132460 3544
rect 132592 3596 132644 3602
rect 132592 3538 132644 3544
rect 133788 3596 133840 3602
rect 133788 3538 133840 3544
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3538
rect 129016 480 129044 3538
rect 130212 480 130240 3538
rect 131408 480 131436 3538
rect 132604 480 132632 3538
rect 135180 626 135208 478926
rect 277398 478887 277454 478896
rect 279148 478576 279200 478582
rect 279148 478518 279200 478524
rect 277398 476776 277454 476785
rect 277398 476711 277454 476720
rect 277412 476134 277440 476711
rect 277400 476128 277452 476134
rect 277400 476070 277452 476076
rect 278686 474736 278742 474745
rect 278686 474671 278742 474680
rect 278700 473414 278728 474671
rect 278688 473408 278740 473414
rect 278688 473350 278740 473356
rect 278686 472560 278742 472569
rect 278686 472495 278742 472504
rect 278700 472054 278728 472495
rect 278688 472048 278740 472054
rect 278688 471990 278740 471996
rect 277858 470384 277914 470393
rect 277858 470319 277914 470328
rect 277872 469266 277900 470319
rect 277860 469260 277912 469266
rect 277860 469202 277912 469208
rect 278686 468344 278742 468353
rect 278686 468279 278742 468288
rect 278700 467906 278728 468279
rect 278688 467900 278740 467906
rect 278688 467842 278740 467848
rect 278686 466168 278742 466177
rect 278686 466103 278742 466112
rect 278700 465118 278728 466103
rect 278688 465112 278740 465118
rect 278688 465054 278740 465060
rect 278686 464128 278742 464137
rect 278686 464063 278742 464072
rect 278700 463758 278728 464063
rect 278688 463752 278740 463758
rect 278688 463694 278740 463700
rect 278686 461952 278742 461961
rect 278686 461887 278742 461896
rect 278700 460970 278728 461887
rect 278688 460964 278740 460970
rect 278688 460906 278740 460912
rect 278686 459776 278742 459785
rect 278686 459711 278742 459720
rect 278700 459610 278728 459711
rect 278688 459604 278740 459610
rect 278688 459546 278740 459552
rect 278686 457736 278742 457745
rect 278686 457671 278742 457680
rect 278700 456822 278728 457671
rect 278688 456816 278740 456822
rect 278688 456758 278740 456764
rect 278686 455560 278742 455569
rect 278686 455495 278742 455504
rect 278700 455462 278728 455495
rect 278688 455456 278740 455462
rect 278688 455398 278740 455404
rect 278686 453384 278742 453393
rect 278686 453319 278742 453328
rect 278700 452674 278728 453319
rect 278688 452668 278740 452674
rect 278688 452610 278740 452616
rect 279160 452606 279188 478518
rect 279516 478372 279568 478378
rect 279516 478314 279568 478320
rect 279240 478100 279292 478106
rect 279240 478042 279292 478048
rect 279148 452600 279200 452606
rect 279148 452542 279200 452548
rect 278686 451344 278742 451353
rect 278686 451279 278688 451288
rect 278740 451279 278742 451288
rect 278688 451250 278740 451256
rect 278686 449168 278742 449177
rect 278686 449103 278742 449112
rect 278700 448594 278728 449103
rect 278688 448588 278740 448594
rect 278688 448530 278740 448536
rect 278686 447128 278742 447137
rect 278686 447063 278742 447072
rect 278700 445806 278728 447063
rect 278688 445800 278740 445806
rect 278688 445742 278740 445748
rect 278686 444952 278742 444961
rect 278686 444887 278742 444896
rect 278700 444446 278728 444887
rect 278688 444440 278740 444446
rect 278688 444382 278740 444388
rect 277858 442776 277914 442785
rect 277858 442711 277914 442720
rect 277872 441658 277900 442711
rect 277860 441652 277912 441658
rect 277860 441594 277912 441600
rect 278686 440736 278742 440745
rect 278686 440671 278742 440680
rect 278700 440298 278728 440671
rect 278688 440292 278740 440298
rect 278688 440234 278740 440240
rect 279252 438870 279280 478042
rect 279424 478032 279476 478038
rect 279424 477974 279476 477980
rect 279332 477964 279384 477970
rect 279332 477906 279384 477912
rect 279240 438864 279292 438870
rect 279240 438806 279292 438812
rect 278686 438560 278742 438569
rect 278686 438495 278742 438504
rect 278700 437510 278728 438495
rect 278688 437504 278740 437510
rect 278688 437446 278740 437452
rect 278042 436384 278098 436393
rect 278042 436319 278098 436328
rect 278056 436150 278084 436319
rect 278044 436144 278096 436150
rect 278044 436086 278096 436092
rect 278686 434344 278742 434353
rect 278686 434279 278742 434288
rect 278700 433362 278728 434279
rect 278688 433356 278740 433362
rect 278688 433298 278740 433304
rect 278686 432168 278742 432177
rect 278686 432103 278742 432112
rect 278700 432002 278728 432103
rect 278688 431996 278740 432002
rect 278688 431938 278740 431944
rect 277674 430128 277730 430137
rect 277674 430063 277730 430072
rect 277688 429214 277716 430063
rect 277676 429208 277728 429214
rect 277676 429150 277728 429156
rect 278686 427952 278742 427961
rect 278686 427887 278742 427896
rect 278700 427854 278728 427887
rect 278688 427848 278740 427854
rect 278688 427790 278740 427796
rect 278686 425776 278742 425785
rect 278686 425711 278742 425720
rect 278700 425134 278728 425711
rect 278688 425128 278740 425134
rect 278688 425070 278740 425076
rect 279344 425066 279372 477906
rect 279332 425060 279384 425066
rect 279332 425002 279384 425008
rect 278686 423736 278742 423745
rect 278686 423671 278688 423680
rect 278740 423671 278742 423680
rect 278688 423642 278740 423648
rect 278686 421560 278742 421569
rect 278686 421495 278742 421504
rect 278700 420986 278728 421495
rect 278688 420980 278740 420986
rect 278688 420922 278740 420928
rect 278686 419520 278742 419529
rect 278686 419455 278742 419464
rect 278700 418198 278728 419455
rect 278688 418192 278740 418198
rect 278688 418134 278740 418140
rect 278686 417344 278742 417353
rect 278686 417279 278742 417288
rect 278700 416838 278728 417279
rect 278688 416832 278740 416838
rect 278688 416774 278740 416780
rect 277858 415168 277914 415177
rect 277858 415103 277914 415112
rect 277872 414050 277900 415103
rect 277860 414044 277912 414050
rect 277860 413986 277912 413992
rect 278686 413128 278742 413137
rect 278686 413063 278742 413072
rect 278700 412690 278728 413063
rect 278688 412684 278740 412690
rect 278688 412626 278740 412632
rect 278686 410952 278742 410961
rect 278686 410887 278742 410896
rect 278700 409902 278728 410887
rect 278688 409896 278740 409902
rect 278688 409838 278740 409844
rect 278686 408776 278742 408785
rect 278686 408711 278742 408720
rect 278700 408542 278728 408711
rect 278688 408536 278740 408542
rect 278688 408478 278740 408484
rect 278686 406736 278742 406745
rect 278686 406671 278742 406680
rect 278700 405754 278728 406671
rect 278688 405748 278740 405754
rect 278688 405690 278740 405696
rect 278686 404560 278742 404569
rect 278686 404495 278742 404504
rect 278700 404394 278728 404495
rect 278688 404388 278740 404394
rect 278688 404330 278740 404336
rect 278410 402520 278466 402529
rect 278410 402455 278466 402464
rect 278424 401674 278452 402455
rect 278412 401668 278464 401674
rect 278412 401610 278464 401616
rect 278686 400344 278742 400353
rect 278686 400279 278742 400288
rect 278700 400246 278728 400279
rect 278688 400240 278740 400246
rect 278688 400182 278740 400188
rect 278686 398168 278742 398177
rect 278686 398103 278742 398112
rect 278700 397526 278728 398103
rect 278688 397520 278740 397526
rect 278688 397462 278740 397468
rect 278686 396128 278742 396137
rect 278686 396063 278688 396072
rect 278740 396063 278742 396072
rect 278688 396034 278740 396040
rect 278686 393952 278742 393961
rect 278686 393887 278742 393896
rect 278700 393378 278728 393887
rect 278688 393372 278740 393378
rect 278688 393314 278740 393320
rect 278318 391776 278374 391785
rect 278318 391711 278374 391720
rect 278332 390590 278360 391711
rect 278320 390584 278372 390590
rect 278320 390526 278372 390532
rect 278686 389736 278742 389745
rect 278686 389671 278742 389680
rect 278700 389230 278728 389671
rect 278688 389224 278740 389230
rect 278688 389166 278740 389172
rect 277858 387560 277914 387569
rect 277858 387495 277914 387504
rect 277872 386442 277900 387495
rect 277860 386436 277912 386442
rect 277860 386378 277912 386384
rect 277674 385520 277730 385529
rect 277674 385455 277730 385464
rect 277688 385082 277716 385455
rect 277676 385076 277728 385082
rect 277676 385018 277728 385024
rect 278686 383344 278742 383353
rect 278686 383279 278742 383288
rect 278700 382294 278728 383279
rect 278688 382288 278740 382294
rect 278688 382230 278740 382236
rect 278042 381168 278098 381177
rect 278042 381103 278098 381112
rect 278056 380934 278084 381103
rect 278044 380928 278096 380934
rect 278044 380870 278096 380876
rect 278686 379128 278742 379137
rect 278686 379063 278742 379072
rect 278700 378214 278728 379063
rect 278688 378208 278740 378214
rect 278688 378150 278740 378156
rect 278686 376952 278742 376961
rect 278686 376887 278742 376896
rect 278700 376786 278728 376887
rect 278688 376780 278740 376786
rect 278688 376722 278740 376728
rect 278410 374912 278466 374921
rect 278410 374847 278466 374856
rect 278424 374066 278452 374847
rect 278412 374060 278464 374066
rect 278412 374002 278464 374008
rect 278042 372736 278098 372745
rect 278042 372671 278098 372680
rect 278056 372638 278084 372671
rect 278044 372632 278096 372638
rect 278044 372574 278096 372580
rect 278318 370560 278374 370569
rect 278318 370495 278374 370504
rect 278332 369918 278360 370495
rect 278320 369912 278372 369918
rect 278320 369854 278372 369860
rect 278688 368552 278740 368558
rect 278686 368520 278688 368529
rect 278740 368520 278742 368529
rect 278686 368455 278742 368464
rect 278686 366344 278742 366353
rect 278686 366279 278742 366288
rect 278700 365770 278728 366279
rect 278688 365764 278740 365770
rect 278688 365706 278740 365712
rect 277858 364168 277914 364177
rect 277858 364103 277914 364112
rect 277872 362982 277900 364103
rect 277860 362976 277912 362982
rect 277860 362918 277912 362924
rect 278686 362128 278742 362137
rect 278686 362063 278742 362072
rect 278700 361622 278728 362063
rect 278688 361616 278740 361622
rect 278688 361558 278740 361564
rect 277858 359952 277914 359961
rect 277858 359887 277914 359896
rect 277872 358834 277900 359887
rect 277860 358828 277912 358834
rect 277860 358770 277912 358776
rect 278686 357912 278742 357921
rect 278686 357847 278742 357856
rect 278700 357474 278728 357847
rect 278688 357468 278740 357474
rect 278688 357410 278740 357416
rect 278686 355736 278742 355745
rect 278686 355671 278742 355680
rect 278700 354754 278728 355671
rect 278688 354748 278740 354754
rect 278688 354690 278740 354696
rect 278042 353560 278098 353569
rect 278042 353495 278098 353504
rect 278056 353326 278084 353495
rect 278044 353320 278096 353326
rect 278044 353262 278096 353268
rect 278686 351520 278742 351529
rect 278686 351455 278742 351464
rect 278700 350606 278728 351455
rect 278688 350600 278740 350606
rect 278688 350542 278740 350548
rect 278686 349344 278742 349353
rect 278686 349279 278742 349288
rect 278700 349178 278728 349279
rect 278688 349172 278740 349178
rect 278688 349114 278740 349120
rect 278686 347168 278742 347177
rect 278686 347103 278742 347112
rect 278700 346458 278728 347103
rect 278688 346452 278740 346458
rect 278688 346394 278740 346400
rect 278686 345128 278742 345137
rect 278686 345063 278688 345072
rect 278740 345063 278742 345072
rect 278688 345034 278740 345040
rect 278318 342952 278374 342961
rect 278318 342887 278374 342896
rect 278332 342310 278360 342887
rect 278320 342304 278372 342310
rect 278320 342246 278372 342252
rect 278688 340944 278740 340950
rect 278686 340912 278688 340921
rect 278740 340912 278742 340921
rect 278686 340847 278742 340856
rect 278686 338736 278742 338745
rect 278686 338671 278742 338680
rect 278700 338162 278728 338671
rect 278688 338156 278740 338162
rect 278688 338098 278740 338104
rect 277858 336560 277914 336569
rect 277858 336495 277914 336504
rect 277872 335374 277900 336495
rect 277860 335368 277912 335374
rect 277860 335310 277912 335316
rect 278686 334520 278742 334529
rect 278686 334455 278742 334464
rect 278700 334014 278728 334455
rect 278688 334008 278740 334014
rect 278688 333950 278740 333956
rect 278686 332344 278742 332353
rect 278686 332279 278742 332288
rect 278700 331294 278728 332279
rect 278688 331288 278740 331294
rect 278688 331230 278740 331236
rect 278686 330304 278742 330313
rect 278686 330239 278742 330248
rect 278700 329866 278728 330239
rect 278688 329860 278740 329866
rect 278688 329802 278740 329808
rect 278686 328128 278742 328137
rect 278686 328063 278742 328072
rect 278700 327146 278728 328063
rect 278688 327140 278740 327146
rect 278688 327082 278740 327088
rect 278042 325952 278098 325961
rect 278042 325887 278098 325896
rect 278056 325718 278084 325887
rect 278044 325712 278096 325718
rect 278044 325654 278096 325660
rect 277674 323912 277730 323921
rect 277674 323847 277730 323856
rect 277688 322998 277716 323847
rect 277676 322992 277728 322998
rect 277676 322934 277728 322940
rect 278042 321736 278098 321745
rect 278042 321671 278098 321680
rect 278056 321638 278084 321671
rect 278044 321632 278096 321638
rect 278044 321574 278096 321580
rect 278686 319560 278742 319569
rect 278686 319495 278742 319504
rect 278700 318850 278728 319495
rect 278688 318844 278740 318850
rect 278688 318786 278740 318792
rect 278686 317520 278742 317529
rect 278686 317455 278688 317464
rect 278740 317455 278742 317464
rect 278688 317426 278740 317432
rect 278686 315344 278742 315353
rect 278686 315279 278742 315288
rect 278700 314702 278728 315279
rect 278688 314696 278740 314702
rect 278688 314638 278740 314644
rect 278688 313336 278740 313342
rect 278686 313304 278688 313313
rect 278740 313304 278742 313313
rect 278686 313239 278742 313248
rect 278686 311128 278742 311137
rect 278686 311063 278742 311072
rect 278700 310554 278728 311063
rect 278688 310548 278740 310554
rect 278688 310490 278740 310496
rect 277858 308952 277914 308961
rect 277858 308887 277914 308896
rect 277872 307834 277900 308887
rect 277860 307828 277912 307834
rect 277860 307770 277912 307776
rect 278686 306912 278742 306921
rect 278686 306847 278742 306856
rect 278700 306406 278728 306847
rect 278688 306400 278740 306406
rect 278688 306342 278740 306348
rect 278686 304736 278742 304745
rect 278686 304671 278742 304680
rect 278700 303686 278728 304671
rect 278688 303680 278740 303686
rect 278688 303622 278740 303628
rect 278686 302560 278742 302569
rect 278686 302495 278742 302504
rect 278700 302258 278728 302495
rect 278688 302252 278740 302258
rect 278688 302194 278740 302200
rect 278686 300520 278742 300529
rect 278686 300455 278742 300464
rect 278700 299538 278728 300455
rect 278688 299532 278740 299538
rect 278688 299474 278740 299480
rect 278686 298344 278742 298353
rect 278686 298279 278742 298288
rect 278700 298178 278728 298279
rect 278688 298172 278740 298178
rect 278688 298114 278740 298120
rect 278686 296304 278742 296313
rect 278686 296239 278742 296248
rect 278700 295390 278728 296239
rect 278688 295384 278740 295390
rect 278688 295326 278740 295332
rect 278686 294128 278742 294137
rect 278686 294063 278742 294072
rect 278700 294030 278728 294063
rect 278688 294024 278740 294030
rect 278688 293966 278740 293972
rect 278686 291952 278742 291961
rect 278686 291887 278742 291896
rect 278700 291242 278728 291887
rect 278688 291236 278740 291242
rect 278688 291178 278740 291184
rect 278686 289912 278742 289921
rect 278686 289847 278688 289856
rect 278740 289847 278742 289856
rect 278688 289818 278740 289824
rect 278686 287736 278742 287745
rect 278686 287671 278742 287680
rect 278700 287094 278728 287671
rect 278688 287088 278740 287094
rect 278688 287030 278740 287036
rect 278688 285728 278740 285734
rect 278686 285696 278688 285705
rect 278740 285696 278742 285705
rect 278686 285631 278742 285640
rect 278686 283520 278742 283529
rect 278686 283455 278742 283464
rect 278700 282946 278728 283455
rect 278688 282940 278740 282946
rect 278688 282882 278740 282888
rect 277858 281344 277914 281353
rect 277858 281279 277914 281288
rect 277872 280226 277900 281279
rect 277860 280220 277912 280226
rect 277860 280162 277912 280168
rect 279436 280158 279464 477974
rect 279528 295322 279556 478314
rect 279620 309126 279648 479062
rect 279712 324290 279740 479130
rect 279976 479052 280028 479058
rect 279976 478994 280028 479000
rect 279884 478984 279936 478990
rect 279884 478926 279936 478932
rect 279792 478440 279844 478446
rect 279792 478382 279844 478388
rect 279804 338094 279832 478382
rect 279896 367062 279924 478926
rect 279988 380866 280016 478994
rect 280068 478508 280120 478514
rect 280068 478450 280120 478456
rect 280080 396030 280108 478450
rect 280068 396024 280120 396030
rect 280068 395966 280120 395972
rect 279976 380860 280028 380866
rect 279976 380802 280028 380808
rect 279884 367056 279936 367062
rect 279884 366998 279936 367004
rect 279792 338088 279844 338094
rect 279792 338030 279844 338036
rect 279700 324284 279752 324290
rect 279700 324226 279752 324232
rect 279608 309120 279660 309126
rect 279608 309062 279660 309068
rect 279516 295316 279568 295322
rect 279516 295258 279568 295264
rect 279424 280152 279476 280158
rect 279424 280094 279476 280100
rect 278686 279304 278742 279313
rect 278686 279239 278742 279248
rect 278700 278798 278728 279239
rect 278688 278792 278740 278798
rect 278688 278734 278740 278740
rect 278686 277128 278742 277137
rect 278686 277063 278742 277072
rect 278700 276078 278728 277063
rect 278688 276072 278740 276078
rect 278688 276014 278740 276020
rect 278042 274952 278098 274961
rect 278042 274887 278098 274896
rect 278056 274718 278084 274887
rect 278044 274712 278096 274718
rect 278044 274654 278096 274660
rect 278686 272912 278742 272921
rect 278686 272847 278742 272856
rect 278700 271930 278728 272847
rect 278688 271924 278740 271930
rect 278688 271866 278740 271872
rect 278686 270736 278742 270745
rect 278686 270671 278742 270680
rect 278700 270570 278728 270671
rect 278688 270564 278740 270570
rect 278688 270506 278740 270512
rect 278686 268696 278742 268705
rect 278686 268631 278742 268640
rect 278700 267782 278728 268631
rect 278688 267776 278740 267782
rect 278688 267718 278740 267724
rect 278042 266520 278098 266529
rect 278042 266455 278098 266464
rect 278056 266422 278084 266455
rect 278044 266416 278096 266422
rect 278044 266358 278096 266364
rect 278686 264344 278742 264353
rect 278686 264279 278742 264288
rect 278700 263634 278728 264279
rect 278688 263628 278740 263634
rect 278688 263570 278740 263576
rect 278686 262304 278742 262313
rect 278686 262239 278688 262248
rect 278740 262239 278742 262248
rect 278688 262210 278740 262216
rect 278318 260128 278374 260137
rect 278318 260063 278374 260072
rect 278332 259486 278360 260063
rect 278320 259480 278372 259486
rect 278320 259422 278372 259428
rect 277858 257952 277914 257961
rect 277858 257887 277914 257896
rect 277872 256766 277900 257887
rect 277860 256760 277912 256766
rect 277860 256702 277912 256708
rect 278686 255912 278742 255921
rect 278686 255847 278742 255856
rect 278700 255338 278728 255847
rect 278688 255332 278740 255338
rect 278688 255274 278740 255280
rect 277858 253736 277914 253745
rect 277858 253671 277914 253680
rect 277872 252618 277900 253671
rect 277860 252612 277912 252618
rect 277860 252554 277912 252560
rect 278686 251696 278742 251705
rect 278686 251631 278742 251640
rect 278700 251258 278728 251631
rect 278688 251252 278740 251258
rect 278688 251194 278740 251200
rect 278686 249520 278742 249529
rect 278686 249455 278742 249464
rect 278700 248470 278728 249455
rect 278688 248464 278740 248470
rect 278688 248406 278740 248412
rect 278042 247344 278098 247353
rect 278042 247279 278098 247288
rect 277398 243128 277454 243137
rect 277398 243063 277454 243072
rect 277412 242962 277440 243063
rect 277400 242956 277452 242962
rect 277400 242898 277452 242904
rect 278056 3466 278084 247279
rect 278134 245304 278190 245313
rect 278134 245239 278190 245248
rect 278148 3534 278176 245239
rect 278686 241088 278742 241097
rect 278686 241023 278742 241032
rect 278700 240174 278728 241023
rect 280158 240816 280214 240825
rect 280158 240751 280214 240760
rect 280172 240718 280200 240751
rect 280908 240718 280936 517686
rect 283472 482860 283524 482866
rect 283472 482802 283524 482808
rect 281356 482724 281408 482730
rect 281356 482666 281408 482672
rect 281368 479890 281396 482666
rect 283484 479890 283512 482802
rect 285600 479890 285628 517822
rect 288348 517676 288400 517682
rect 288348 517618 288400 517624
rect 288360 482594 288388 517618
rect 289728 517608 289780 517614
rect 289728 517550 289780 517556
rect 287888 482588 287940 482594
rect 287888 482530 287940 482536
rect 288348 482588 288400 482594
rect 288348 482530 288400 482536
rect 287900 479890 287928 482530
rect 289740 480026 289768 517550
rect 289740 479998 289814 480026
rect 281060 479862 281396 479890
rect 283176 479862 283512 479890
rect 285384 479862 285628 479890
rect 287592 479862 287928 479890
rect 289786 479876 289814 479998
rect 292500 479754 292528 518366
rect 295248 518356 295300 518362
rect 295248 518298 295300 518304
rect 295260 482594 295288 518298
rect 296628 517948 296680 517954
rect 296628 517890 296680 517896
rect 294512 482588 294564 482594
rect 294512 482530 294564 482536
rect 295248 482588 295300 482594
rect 295248 482530 295300 482536
rect 294524 479890 294552 482530
rect 296640 479890 296668 517890
rect 297376 482322 297404 540223
rect 297468 482934 297496 598023
rect 297456 482928 297508 482934
rect 297456 482870 297508 482876
rect 297560 482798 297588 599791
rect 297548 482792 297600 482798
rect 297548 482734 297600 482740
rect 297652 482662 297680 600879
rect 297640 482656 297692 482662
rect 297640 482598 297692 482604
rect 297744 482526 297772 602511
rect 297836 483002 297864 603735
rect 297824 482996 297876 483002
rect 297824 482938 297876 482944
rect 297732 482520 297784 482526
rect 297732 482462 297784 482468
rect 297928 482458 297956 605367
rect 297916 482452 297968 482458
rect 297916 482394 297968 482400
rect 298020 482390 298048 606591
rect 299388 518016 299440 518022
rect 299388 517958 299440 517964
rect 299400 482594 299428 517958
rect 299572 482996 299624 483002
rect 299572 482938 299624 482944
rect 298928 482588 298980 482594
rect 298928 482530 298980 482536
rect 299388 482588 299440 482594
rect 299388 482530 299440 482536
rect 298008 482384 298060 482390
rect 298008 482326 298060 482332
rect 297364 482316 297416 482322
rect 297364 482258 297416 482264
rect 298940 479890 298968 482530
rect 299584 482526 299612 482938
rect 299572 482520 299624 482526
rect 299572 482462 299624 482468
rect 294216 479862 294552 479890
rect 296424 479862 296668 479890
rect 298632 479862 298968 479890
rect 300596 479806 300624 699654
rect 332520 610638 332548 703520
rect 348804 700738 348832 703520
rect 348792 700732 348844 700738
rect 348792 700674 348844 700680
rect 364996 699718 365024 703520
rect 397472 699990 397500 703520
rect 413664 700806 413692 703520
rect 413652 700800 413704 700806
rect 413652 700742 413704 700748
rect 397460 699984 397512 699990
rect 397460 699926 397512 699932
rect 398748 699984 398800 699990
rect 398748 699926 398800 699932
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 365628 699712 365680 699718
rect 365628 699654 365680 699660
rect 365640 610706 365668 699654
rect 373632 612808 373684 612814
rect 373630 612776 373632 612785
rect 379612 612808 379664 612814
rect 373684 612776 373686 612785
rect 379612 612750 379664 612756
rect 373630 612711 373686 612720
rect 365628 610700 365680 610706
rect 365628 610642 365680 610648
rect 332508 610632 332560 610638
rect 332508 610574 332560 610580
rect 378048 599004 378100 599010
rect 378048 598946 378100 598952
rect 318708 518900 318760 518906
rect 327172 518900 327224 518906
rect 318708 518842 318760 518848
rect 317328 518832 317380 518838
rect 314566 518800 314622 518809
rect 307576 518764 307628 518770
rect 314566 518735 314622 518744
rect 317326 518800 317328 518809
rect 318720 518809 318748 518842
rect 325436 518838 325464 518869
rect 327172 518842 327224 518848
rect 325424 518832 325476 518838
rect 317380 518800 317382 518809
rect 317326 518735 317382 518744
rect 318706 518800 318762 518809
rect 318706 518735 318762 518744
rect 321742 518800 321798 518809
rect 321742 518735 321798 518744
rect 323122 518800 323178 518809
rect 323122 518735 323178 518744
rect 324318 518800 324374 518809
rect 324318 518735 324320 518744
rect 307576 518706 307628 518712
rect 303618 518256 303674 518265
rect 303618 518191 303620 518200
rect 303672 518191 303674 518200
rect 303620 518162 303672 518168
rect 303528 518084 303580 518090
rect 303528 518026 303580 518032
rect 300676 517812 300728 517818
rect 300676 517754 300728 517760
rect 300688 479890 300716 517754
rect 303540 480026 303568 518026
rect 303632 517750 303660 518162
rect 306288 518152 306340 518158
rect 306288 518094 306340 518100
rect 303620 517744 303672 517750
rect 303620 517686 303672 517692
rect 306300 482254 306328 518094
rect 305552 482248 305604 482254
rect 305552 482190 305604 482196
rect 306288 482248 306340 482254
rect 306288 482190 306340 482196
rect 303356 479998 303568 480026
rect 303356 479890 303384 479998
rect 305564 479890 305592 482190
rect 307588 479890 307616 518706
rect 314580 518702 314608 518735
rect 314568 518696 314620 518702
rect 314568 518638 314620 518644
rect 315946 518664 316002 518673
rect 315946 518599 316002 518608
rect 317326 518664 317382 518673
rect 317326 518599 317382 518608
rect 320086 518664 320142 518673
rect 320086 518599 320088 518608
rect 315960 518498 315988 518599
rect 317340 518566 317368 518599
rect 320140 518599 320142 518608
rect 320088 518570 320140 518576
rect 317328 518560 317380 518566
rect 316038 518528 316094 518537
rect 315948 518492 316000 518498
rect 317328 518502 317380 518508
rect 317510 518528 317566 518537
rect 316038 518463 316094 518472
rect 317510 518463 317566 518472
rect 315948 518434 316000 518440
rect 316052 518430 316080 518463
rect 316040 518424 316092 518430
rect 313186 518392 313242 518401
rect 316040 518366 316092 518372
rect 317418 518392 317474 518401
rect 313186 518327 313242 518336
rect 317418 518327 317420 518336
rect 313200 518294 313228 518327
rect 317472 518327 317474 518336
rect 317420 518298 317472 518304
rect 313188 518288 313240 518294
rect 313188 518230 313240 518236
rect 314658 518256 314714 518265
rect 314658 518191 314714 518200
rect 312082 517984 312138 517993
rect 312082 517919 312138 517928
rect 312096 517886 312124 517919
rect 312084 517880 312136 517886
rect 312084 517822 312136 517828
rect 314568 517880 314620 517886
rect 314568 517822 314620 517828
rect 310428 517744 310480 517750
rect 310334 517712 310390 517721
rect 310428 517686 310480 517692
rect 313278 517712 313334 517721
rect 310334 517647 310390 517656
rect 307666 517576 307722 517585
rect 307666 517511 307722 517520
rect 309046 517576 309102 517585
rect 309046 517511 309102 517520
rect 310242 517576 310298 517585
rect 310242 517511 310298 517520
rect 307680 483002 307708 517511
rect 307668 482996 307720 483002
rect 307668 482938 307720 482944
rect 309060 482050 309088 517511
rect 309968 482248 310020 482254
rect 309968 482190 310020 482196
rect 309048 482044 309100 482050
rect 309048 481986 309100 481992
rect 309980 479890 310008 482190
rect 310256 482186 310284 517511
rect 310244 482180 310296 482186
rect 310244 482122 310296 482128
rect 310348 482118 310376 517647
rect 310440 482254 310468 517686
rect 313278 517647 313280 517656
rect 313332 517647 313334 517656
rect 313280 517618 313332 517624
rect 311714 517576 311770 517585
rect 311714 517511 311770 517520
rect 311808 517540 311860 517546
rect 311728 482254 311756 517511
rect 311808 517482 311860 517488
rect 310428 482248 310480 482254
rect 310428 482190 310480 482196
rect 311716 482248 311768 482254
rect 311716 482190 311768 482196
rect 310336 482112 310388 482118
rect 310336 482054 310388 482060
rect 311820 480026 311848 517482
rect 311820 479998 311894 480026
rect 300688 479862 300840 479890
rect 303048 479862 303384 479890
rect 305256 479862 305592 479890
rect 307464 479862 307616 479890
rect 309672 479862 310008 479890
rect 311866 479876 311894 479998
rect 292008 479726 292528 479754
rect 300584 479800 300636 479806
rect 314580 479754 314608 517822
rect 314672 517614 314700 518191
rect 317524 517954 317552 518463
rect 321098 518392 321154 518401
rect 321098 518327 321100 518336
rect 321152 518327 321154 518336
rect 321100 518298 321152 518304
rect 321756 518294 321784 518735
rect 323136 518702 323164 518735
rect 324372 518735 324374 518744
rect 325422 518800 325424 518809
rect 327184 518809 327212 518842
rect 340524 518838 340552 518869
rect 331220 518832 331272 518838
rect 325476 518800 325478 518809
rect 325422 518735 325478 518744
rect 326434 518800 326490 518809
rect 326434 518735 326436 518744
rect 324320 518706 324372 518712
rect 323124 518696 323176 518702
rect 323124 518638 323176 518644
rect 324410 518664 324466 518673
rect 324410 518599 324466 518608
rect 324424 518498 324452 518599
rect 325436 518498 325464 518735
rect 326488 518735 326490 518744
rect 327170 518800 327226 518809
rect 327170 518735 327226 518744
rect 328918 518800 328974 518809
rect 328918 518735 328974 518744
rect 330114 518800 330170 518809
rect 340512 518832 340564 518838
rect 331220 518774 331272 518780
rect 332322 518800 332378 518809
rect 330114 518735 330170 518744
rect 326436 518706 326488 518712
rect 326448 518566 326476 518706
rect 327184 518566 327212 518735
rect 328932 518634 328960 518735
rect 328920 518628 328972 518634
rect 328920 518570 328972 518576
rect 326436 518560 326488 518566
rect 327172 518560 327224 518566
rect 326436 518502 326488 518508
rect 327078 518528 327134 518537
rect 324412 518492 324464 518498
rect 324412 518434 324464 518440
rect 325424 518492 325476 518498
rect 327172 518502 327224 518508
rect 327078 518463 327134 518472
rect 325424 518434 325476 518440
rect 321744 518288 321796 518294
rect 321744 518230 321796 518236
rect 322938 518256 322994 518265
rect 322938 518191 322994 518200
rect 322952 518158 322980 518191
rect 322940 518152 322992 518158
rect 318798 518120 318854 518129
rect 318798 518055 318854 518064
rect 321834 518120 321890 518129
rect 322940 518094 322992 518100
rect 321834 518055 321836 518064
rect 318812 518022 318840 518055
rect 321888 518055 321890 518064
rect 321836 518026 321888 518032
rect 327092 518022 327120 518463
rect 330128 518362 330156 518735
rect 331232 518673 331260 518774
rect 332322 518735 332378 518744
rect 335542 518800 335598 518809
rect 335542 518735 335544 518744
rect 332336 518702 332364 518735
rect 335596 518735 335598 518744
rect 336738 518800 336794 518809
rect 336738 518735 336794 518744
rect 337198 518800 337254 518809
rect 337198 518735 337254 518744
rect 339958 518800 340014 518809
rect 339958 518735 340014 518744
rect 340510 518800 340512 518809
rect 369860 518832 369912 518838
rect 340564 518800 340566 518809
rect 340510 518735 340566 518744
rect 341614 518800 341670 518809
rect 341614 518735 341670 518744
rect 342994 518800 343050 518809
rect 342994 518735 343050 518744
rect 344190 518800 344246 518809
rect 344190 518735 344246 518744
rect 345478 518800 345534 518809
rect 345478 518735 345480 518744
rect 335544 518706 335596 518712
rect 332324 518696 332376 518702
rect 331218 518664 331274 518673
rect 332324 518638 332376 518644
rect 331218 518599 331274 518608
rect 330116 518356 330168 518362
rect 330116 518298 330168 518304
rect 331232 518294 331260 518599
rect 336648 518560 336700 518566
rect 333426 518528 333482 518537
rect 333426 518463 333482 518472
rect 334162 518528 334218 518537
rect 336752 518514 336780 518735
rect 337212 518702 337240 518735
rect 337200 518696 337252 518702
rect 337200 518638 337252 518644
rect 338118 518664 338174 518673
rect 338118 518599 338174 518608
rect 338132 518566 338160 518599
rect 336700 518508 336780 518514
rect 336648 518502 336780 518508
rect 338120 518560 338172 518566
rect 338120 518502 338172 518508
rect 334162 518463 334164 518472
rect 333440 518430 333468 518463
rect 334216 518463 334218 518472
rect 335176 518492 335228 518498
rect 334164 518434 334216 518440
rect 336660 518486 336780 518502
rect 335176 518434 335228 518440
rect 333428 518424 333480 518430
rect 333428 518366 333480 518372
rect 335188 518294 335216 518434
rect 339972 518362 340000 518735
rect 339960 518356 340012 518362
rect 339960 518298 340012 518304
rect 331220 518288 331272 518294
rect 331220 518230 331272 518236
rect 335176 518288 335228 518294
rect 335176 518230 335228 518236
rect 340524 518022 340552 518735
rect 341628 518634 341656 518735
rect 341616 518628 341668 518634
rect 341616 518570 341668 518576
rect 342168 518628 342220 518634
rect 342168 518570 342220 518576
rect 318800 518016 318852 518022
rect 318800 517958 318852 517964
rect 327080 518016 327132 518022
rect 340512 518016 340564 518022
rect 327080 517958 327132 517964
rect 331218 517984 331274 517993
rect 317512 517948 317564 517954
rect 331218 517919 331220 517928
rect 317512 517890 317564 517896
rect 331272 517919 331274 517928
rect 332598 517984 332654 517993
rect 340512 517958 340564 517964
rect 332598 517919 332654 517928
rect 331220 517890 331272 517896
rect 332612 517886 332640 517919
rect 332600 517880 332652 517886
rect 320178 517848 320234 517857
rect 332600 517822 332652 517828
rect 333978 517848 334034 517857
rect 320178 517783 320180 517792
rect 320232 517783 320234 517792
rect 321468 517812 321520 517818
rect 320180 517754 320232 517760
rect 333978 517783 334034 517792
rect 321468 517754 321520 517760
rect 314660 517608 314712 517614
rect 314660 517550 314712 517556
rect 317328 517608 317380 517614
rect 317328 517550 317380 517556
rect 317340 481982 317368 517550
rect 321480 481982 321508 517754
rect 333992 517750 334020 517783
rect 322848 517744 322900 517750
rect 328368 517744 328420 517750
rect 322848 517686 322900 517692
rect 324318 517712 324374 517721
rect 316500 481976 316552 481982
rect 316500 481918 316552 481924
rect 317328 481976 317380 481982
rect 317328 481918 317380 481924
rect 320916 481976 320968 481982
rect 320916 481918 320968 481924
rect 321468 481976 321520 481982
rect 321468 481918 321520 481924
rect 316512 479890 316540 481918
rect 318708 481840 318760 481846
rect 318708 481782 318760 481788
rect 318720 479890 318748 481782
rect 320928 479890 320956 481918
rect 322860 480162 322888 517686
rect 333980 517744 334032 517750
rect 328368 517686 328420 517692
rect 329838 517712 329894 517721
rect 324318 517647 324320 517656
rect 324372 517647 324374 517656
rect 326344 517676 326396 517682
rect 324320 517618 324372 517624
rect 326344 517618 326396 517624
rect 325698 517576 325754 517585
rect 325698 517511 325700 517520
rect 325752 517511 325754 517520
rect 325700 517482 325752 517488
rect 325332 481908 325384 481914
rect 325332 481850 325384 481856
rect 316204 479862 316540 479890
rect 318412 479862 318748 479890
rect 320620 479862 320956 479890
rect 322814 480134 322888 480162
rect 322814 479876 322842 480134
rect 325344 479890 325372 481850
rect 326356 481846 326384 517618
rect 327724 517608 327776 517614
rect 327724 517550 327776 517556
rect 327540 481976 327592 481982
rect 327540 481918 327592 481924
rect 326344 481840 326396 481846
rect 326344 481782 326396 481788
rect 327552 479890 327580 481918
rect 327736 481914 327764 517550
rect 328380 481982 328408 517686
rect 332598 517712 332654 517721
rect 329838 517647 329840 517656
rect 329892 517647 329894 517656
rect 330484 517676 330536 517682
rect 329840 517618 329892 517624
rect 333980 517686 334032 517692
rect 335726 517712 335782 517721
rect 332598 517647 332654 517656
rect 335726 517647 335728 517656
rect 330484 517618 330536 517624
rect 328458 517576 328514 517585
rect 328458 517511 328460 517520
rect 328512 517511 328514 517520
rect 328460 517482 328512 517488
rect 330496 481982 330524 517618
rect 332612 517614 332640 517647
rect 335780 517647 335782 517656
rect 338118 517712 338174 517721
rect 338118 517647 338174 517656
rect 339498 517712 339554 517721
rect 339498 517647 339554 517656
rect 335728 517618 335780 517624
rect 338132 517614 338160 517647
rect 332600 517608 332652 517614
rect 332600 517550 332652 517556
rect 333888 517608 333940 517614
rect 338120 517608 338172 517614
rect 333888 517550 333940 517556
rect 336738 517576 336794 517585
rect 333244 517540 333296 517546
rect 333244 517482 333296 517488
rect 333256 481982 333284 517482
rect 328368 481976 328420 481982
rect 328368 481918 328420 481924
rect 329748 481976 329800 481982
rect 329748 481918 329800 481924
rect 330484 481976 330536 481982
rect 330484 481918 330536 481924
rect 331956 481976 332008 481982
rect 331956 481918 332008 481924
rect 333244 481976 333296 481982
rect 333244 481918 333296 481924
rect 327724 481908 327776 481914
rect 327724 481850 327776 481856
rect 329760 479890 329788 481918
rect 331968 479890 331996 481918
rect 333900 480162 333928 517550
rect 338120 517550 338172 517556
rect 339406 517576 339462 517585
rect 336738 517511 336740 517520
rect 336792 517511 336794 517520
rect 337384 517540 337436 517546
rect 336740 517482 336792 517488
rect 339512 517546 339540 517647
rect 342180 517614 342208 518570
rect 343008 518430 343036 518735
rect 342996 518424 343048 518430
rect 342996 518366 343048 518372
rect 343548 518424 343600 518430
rect 343548 518366 343600 518372
rect 343560 517954 343588 518366
rect 344204 518294 344232 518735
rect 345532 518735 345534 518744
rect 346490 518800 346546 518809
rect 346490 518735 346546 518744
rect 347686 518800 347742 518809
rect 347686 518735 347742 518744
rect 348606 518800 348662 518809
rect 369860 518774 369912 518780
rect 348606 518735 348662 518744
rect 345480 518706 345532 518712
rect 346504 518702 346532 518735
rect 346492 518696 346544 518702
rect 346492 518638 346544 518644
rect 347700 518566 347728 518735
rect 348620 518634 348648 518735
rect 347780 518628 347832 518634
rect 347780 518570 347832 518576
rect 348608 518628 348660 518634
rect 348608 518570 348660 518576
rect 350540 518628 350592 518634
rect 350540 518570 350592 518576
rect 357440 518628 357492 518634
rect 357440 518570 357492 518576
rect 362224 518628 362276 518634
rect 362224 518570 362276 518576
rect 347688 518560 347740 518566
rect 347688 518502 347740 518508
rect 347792 518362 347820 518570
rect 350552 518430 350580 518570
rect 357452 518430 357480 518570
rect 362236 518498 362264 518570
rect 369872 518498 369900 518774
rect 362224 518492 362276 518498
rect 362224 518434 362276 518440
rect 369860 518492 369912 518498
rect 369860 518434 369912 518440
rect 350540 518424 350592 518430
rect 350540 518366 350592 518372
rect 357440 518424 357492 518430
rect 357440 518366 357492 518372
rect 373908 518424 373960 518430
rect 373908 518366 373960 518372
rect 347780 518356 347832 518362
rect 347780 518298 347832 518304
rect 362868 518356 362920 518362
rect 362868 518298 362920 518304
rect 344192 518288 344244 518294
rect 344192 518230 344244 518236
rect 344928 518288 344980 518294
rect 344928 518230 344980 518236
rect 361488 518288 361540 518294
rect 361488 518230 361540 518236
rect 343548 517948 343600 517954
rect 343548 517890 343600 517896
rect 342902 517712 342958 517721
rect 342902 517647 342958 517656
rect 344282 517712 344338 517721
rect 344940 517682 344968 518230
rect 358728 518152 358780 518158
rect 358728 518094 358780 518100
rect 355968 518084 356020 518090
rect 355968 518026 356020 518032
rect 346306 517712 346362 517721
rect 344282 517647 344338 517656
rect 344928 517676 344980 517682
rect 342168 517608 342220 517614
rect 340786 517576 340842 517585
rect 339406 517511 339462 517520
rect 339500 517540 339552 517546
rect 337384 517482 337436 517488
rect 337396 481982 337424 517482
rect 339420 481982 339448 517511
rect 342168 517550 342220 517556
rect 340786 517511 340842 517520
rect 339500 517482 339552 517488
rect 336372 481976 336424 481982
rect 336372 481918 336424 481924
rect 337384 481976 337436 481982
rect 337384 481918 337436 481924
rect 338580 481976 338632 481982
rect 338580 481918 338632 481924
rect 339408 481976 339460 481982
rect 339408 481918 339460 481924
rect 325036 479862 325372 479890
rect 327244 479862 327580 479890
rect 329452 479862 329788 479890
rect 331660 479862 331996 479890
rect 333854 480134 333928 480162
rect 333854 479876 333882 480134
rect 336384 479890 336412 481918
rect 338592 479890 338620 481918
rect 340800 479890 340828 517511
rect 342916 479890 342944 517647
rect 336076 479862 336412 479890
rect 338284 479862 338620 479890
rect 340492 479862 340828 479890
rect 342700 479862 342944 479890
rect 300584 479742 300636 479748
rect 314088 479726 314608 479754
rect 344296 479754 344324 517647
rect 346306 517647 346362 517656
rect 348422 517712 348478 517721
rect 348422 517647 348478 517656
rect 348974 517712 349030 517721
rect 348974 517647 349030 517656
rect 344928 517618 344980 517624
rect 346320 481982 346348 517647
rect 348436 481982 348464 517647
rect 346308 481976 346360 481982
rect 346308 481918 346360 481924
rect 346768 481976 346820 481982
rect 346768 481918 346820 481924
rect 348424 481976 348476 481982
rect 348424 481918 348476 481924
rect 346780 479890 346808 481918
rect 348988 481846 349016 517647
rect 349066 517576 349122 517585
rect 349066 517511 349122 517520
rect 349080 482066 349108 517511
rect 349080 482038 349292 482066
rect 349264 481982 349292 482038
rect 349160 481976 349212 481982
rect 349160 481918 349212 481924
rect 349252 481976 349304 481982
rect 349252 481918 349304 481924
rect 351092 481976 351144 481982
rect 351092 481918 351144 481924
rect 348976 481840 349028 481846
rect 348976 481782 349028 481788
rect 349172 479890 349200 481918
rect 351104 479890 351132 481918
rect 353300 481840 353352 481846
rect 353300 481782 353352 481788
rect 353312 479890 353340 481782
rect 355980 479890 356008 518026
rect 358740 481982 358768 518094
rect 358268 481976 358320 481982
rect 358268 481918 358320 481924
rect 358728 481976 358780 481982
rect 358728 481918 358780 481924
rect 358280 479890 358308 481918
rect 361500 481914 361528 518230
rect 360568 481908 360620 481914
rect 360568 481850 360620 481856
rect 361488 481908 361540 481914
rect 361488 481850 361540 481856
rect 360580 479890 360608 481850
rect 362222 480040 362278 480049
rect 362222 479975 362278 479984
rect 346780 479862 347116 479890
rect 349172 479862 349324 479890
rect 351104 479862 351440 479890
rect 353312 479862 353648 479890
rect 355856 479862 356008 479890
rect 358064 479862 358308 479890
rect 360272 479862 360608 479890
rect 362236 479777 362264 479975
rect 362880 479890 362908 518298
rect 371240 482248 371292 482254
rect 371240 482190 371292 482196
rect 368756 482180 368808 482186
rect 368756 482122 368808 482128
rect 366548 482112 366600 482118
rect 366548 482054 366600 482060
rect 364340 482044 364392 482050
rect 364340 481986 364392 481992
rect 362480 479862 362908 479890
rect 364352 479890 364380 481986
rect 366560 479890 366588 482054
rect 368768 479890 368796 482122
rect 371252 480162 371280 482190
rect 371252 480134 371326 480162
rect 369950 480040 370006 480049
rect 369950 479975 370006 479984
rect 364352 479862 364688 479890
rect 366560 479862 366896 479890
rect 367192 479868 367244 479874
rect 368768 479862 369104 479890
rect 369964 479874 369992 479975
rect 371298 479876 371326 480134
rect 373920 479890 373948 518366
rect 376024 482248 376076 482254
rect 376024 482190 376076 482196
rect 376036 479890 376064 482190
rect 378060 479890 378088 598946
rect 379624 549409 379652 612750
rect 379980 610428 380032 610434
rect 379980 610370 380032 610376
rect 379992 609657 380020 610370
rect 379702 609648 379758 609657
rect 379702 609583 379758 609592
rect 379978 609648 380034 609657
rect 379978 609583 380034 609592
rect 379610 549400 379666 549409
rect 379610 549335 379666 549344
rect 379520 538280 379572 538286
rect 379520 538222 379572 538228
rect 379532 536110 379560 538222
rect 379520 536104 379572 536110
rect 379520 536046 379572 536052
rect 379612 519580 379664 519586
rect 379612 519522 379664 519528
rect 379428 518832 379480 518838
rect 379428 518774 379480 518780
rect 379520 518832 379572 518838
rect 379520 518774 379572 518780
rect 379440 518634 379468 518774
rect 379532 518634 379560 518774
rect 379428 518628 379480 518634
rect 379428 518570 379480 518576
rect 379520 518628 379572 518634
rect 379520 518570 379572 518576
rect 379624 514078 379652 519522
rect 379612 514072 379664 514078
rect 379612 514014 379664 514020
rect 379612 499588 379664 499594
rect 379612 499530 379664 499536
rect 379624 494766 379652 499530
rect 379612 494760 379664 494766
rect 379612 494702 379664 494708
rect 379716 482866 379744 609583
rect 389088 605872 389140 605878
rect 389088 605814 389140 605820
rect 387708 604512 387760 604518
rect 387708 604454 387760 604460
rect 384948 603152 385000 603158
rect 384948 603094 385000 603100
rect 383568 601724 383620 601730
rect 383568 601666 383620 601672
rect 380808 600364 380860 600370
rect 380808 600306 380860 600312
rect 379794 540968 379850 540977
rect 379794 540903 379850 540912
rect 379808 538286 379836 540903
rect 379796 538280 379848 538286
rect 379796 538222 379848 538228
rect 379796 536104 379848 536110
rect 379796 536046 379848 536052
rect 379808 519586 379836 536046
rect 379796 519580 379848 519586
rect 379796 519522 379848 519528
rect 379796 514072 379848 514078
rect 379796 514014 379848 514020
rect 379808 499594 379836 514014
rect 379796 499588 379848 499594
rect 379796 499530 379848 499536
rect 379796 494760 379848 494766
rect 379796 494702 379848 494708
rect 379704 482860 379756 482866
rect 379704 482802 379756 482808
rect 379808 482730 379836 494702
rect 379796 482724 379848 482730
rect 379796 482666 379848 482672
rect 380820 480026 380848 600306
rect 383580 482730 383608 601666
rect 382648 482724 382700 482730
rect 382648 482666 382700 482672
rect 383568 482724 383620 482730
rect 383568 482666 383620 482672
rect 380452 479998 380848 480026
rect 380452 479890 380480 479998
rect 382660 479890 382688 482666
rect 384960 480026 384988 603094
rect 387616 482860 387668 482866
rect 387616 482802 387668 482808
rect 387340 482792 387392 482798
rect 387340 482734 387392 482740
rect 386972 482724 387024 482730
rect 386972 482666 387024 482672
rect 384776 479998 384988 480026
rect 384776 479890 384804 479998
rect 386984 479890 387012 482666
rect 387352 480146 387380 482734
rect 387628 482186 387656 482802
rect 387720 482730 387748 604454
rect 388996 518832 389048 518838
rect 388996 518774 389048 518780
rect 389008 518498 389036 518774
rect 388996 518492 389048 518498
rect 388996 518434 389048 518440
rect 387708 482724 387760 482730
rect 387708 482666 387760 482672
rect 387616 482180 387668 482186
rect 387616 482122 387668 482128
rect 387340 480140 387392 480146
rect 387340 480082 387392 480088
rect 389100 479890 389128 605814
rect 393320 518832 393372 518838
rect 393320 518774 393372 518780
rect 393332 518498 393360 518774
rect 393320 518492 393372 518498
rect 393320 518434 393372 518440
rect 390744 482928 390796 482934
rect 390744 482870 390796 482876
rect 369952 479868 370004 479874
rect 367192 479810 367244 479816
rect 373520 479862 373948 479890
rect 375728 479862 376064 479890
rect 377936 479862 378088 479890
rect 380144 479862 380480 479890
rect 382352 479862 382688 479890
rect 384468 479862 384804 479890
rect 386676 479862 387012 479890
rect 388884 479862 389128 479890
rect 390756 479890 390784 482870
rect 397460 482656 397512 482662
rect 397460 482598 397512 482604
rect 392952 482180 393004 482186
rect 392952 482122 393004 482128
rect 392964 479890 392992 482122
rect 395482 480140 395534 480146
rect 395482 480082 395534 480088
rect 390756 479862 391092 479890
rect 392964 479862 393300 479890
rect 395494 479876 395522 480082
rect 397472 479890 397500 482598
rect 397472 479862 397716 479890
rect 398760 479874 398788 699926
rect 429856 699718 429884 703520
rect 462332 700126 462360 703520
rect 478524 700874 478552 703520
rect 478512 700868 478564 700874
rect 478512 700810 478564 700816
rect 462320 700120 462372 700126
rect 462320 700062 462372 700068
rect 463608 700120 463660 700126
rect 463608 700062 463660 700068
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 430488 699712 430540 699718
rect 430488 699654 430540 699660
rect 430500 610774 430528 699654
rect 463620 610842 463648 700062
rect 494808 699718 494836 703520
rect 519084 700868 519136 700874
rect 519084 700810 519136 700816
rect 514850 700360 514906 700369
rect 514850 700295 514906 700304
rect 494796 699712 494848 699718
rect 494796 699654 494848 699660
rect 495348 699712 495400 699718
rect 495348 699654 495400 699660
rect 488540 613420 488592 613426
rect 488540 613362 488592 613368
rect 493968 613420 494020 613426
rect 493968 613362 494020 613368
rect 488552 612814 488580 613362
rect 493980 612814 494008 613362
rect 488540 612808 488592 612814
rect 488538 612776 488540 612785
rect 493968 612808 494020 612814
rect 488592 612776 488594 612785
rect 488538 612711 488594 612720
rect 493966 612776 493968 612785
rect 494020 612776 494022 612785
rect 493966 612711 494022 612720
rect 495360 610910 495388 699654
rect 514864 695745 514892 700295
rect 514850 695736 514906 695745
rect 514850 695671 514906 695680
rect 499580 612808 499632 612814
rect 499580 612750 499632 612756
rect 495348 610904 495400 610910
rect 495348 610846 495400 610852
rect 463608 610836 463660 610842
rect 463608 610778 463660 610784
rect 430488 610768 430540 610774
rect 430488 610710 430540 610716
rect 496452 610428 496504 610434
rect 496452 610370 496504 610376
rect 496464 609929 496492 610370
rect 496450 609920 496506 609929
rect 496450 609855 496506 609864
rect 416778 606112 416834 606121
rect 416778 606047 416834 606056
rect 416792 605878 416820 606047
rect 416780 605872 416832 605878
rect 416780 605814 416832 605820
rect 416778 604888 416834 604897
rect 416778 604823 416834 604832
rect 416792 604518 416820 604823
rect 416780 604512 416832 604518
rect 416780 604454 416832 604460
rect 416778 603256 416834 603265
rect 416778 603191 416834 603200
rect 416792 603158 416820 603191
rect 416780 603152 416832 603158
rect 416780 603094 416832 603100
rect 416778 602032 416834 602041
rect 416778 601967 416834 601976
rect 416792 601730 416820 601967
rect 416780 601724 416832 601730
rect 416780 601666 416832 601672
rect 416778 600536 416834 600545
rect 416778 600471 416834 600480
rect 416792 600370 416820 600471
rect 416780 600364 416832 600370
rect 416780 600306 416832 600312
rect 416778 599312 416834 599321
rect 416778 599247 416834 599256
rect 416792 599010 416820 599247
rect 416780 599004 416832 599010
rect 416780 598946 416832 598952
rect 416778 597680 416834 597689
rect 416778 597615 416834 597624
rect 416792 597582 416820 597615
rect 410524 597576 410576 597582
rect 410524 597518 410576 597524
rect 416780 597576 416832 597582
rect 416780 597518 416832 597524
rect 409144 538280 409196 538286
rect 409144 538222 409196 538228
rect 409156 521626 409184 538222
rect 408500 521620 408552 521626
rect 408500 521562 408552 521568
rect 409144 521620 409196 521626
rect 409144 521562 409196 521568
rect 408512 520946 408540 521562
rect 408500 520940 408552 520946
rect 408500 520882 408552 520888
rect 402888 518832 402940 518838
rect 402888 518774 402940 518780
rect 402900 518634 402928 518774
rect 402888 518628 402940 518634
rect 402888 518570 402940 518576
rect 399576 482588 399628 482594
rect 399576 482530 399628 482536
rect 399588 479890 399616 482530
rect 401784 482520 401836 482526
rect 401784 482462 401836 482468
rect 401796 479890 401824 482462
rect 403992 482452 404044 482458
rect 403992 482394 404044 482400
rect 404004 479890 404032 482394
rect 406200 482384 406252 482390
rect 406200 482326 406252 482332
rect 406212 479890 406240 482326
rect 408512 479890 408540 520882
rect 410536 482254 410564 597518
rect 499592 549545 499620 612750
rect 499578 549536 499634 549545
rect 499578 549471 499634 549480
rect 499578 542056 499634 542065
rect 499578 541991 499634 542000
rect 499592 540977 499620 541991
rect 499578 540968 499634 540977
rect 499578 540903 499634 540912
rect 416778 539744 416834 539753
rect 416778 539679 416834 539688
rect 416792 539646 416820 539679
rect 411168 539640 411220 539646
rect 411168 539582 411220 539588
rect 416780 539640 416832 539646
rect 416780 539582 416832 539588
rect 410524 482248 410576 482254
rect 410524 482190 410576 482196
rect 411180 479890 411208 539582
rect 416778 538384 416834 538393
rect 416778 538319 416834 538328
rect 416792 538286 416820 538319
rect 416780 538280 416832 538286
rect 416780 538222 416832 538228
rect 425610 519752 425666 519761
rect 425610 519687 425666 519696
rect 423678 518256 423734 518265
rect 423678 518191 423680 518200
rect 423732 518191 423734 518200
rect 423680 518162 423732 518168
rect 425624 518090 425652 519687
rect 451280 518832 451332 518838
rect 443182 518800 443238 518809
rect 441620 518764 441672 518770
rect 443182 518735 443184 518744
rect 441620 518706 441672 518712
rect 443236 518735 443238 518744
rect 451278 518800 451280 518809
rect 459560 518832 459612 518838
rect 451332 518800 451334 518809
rect 451278 518735 451334 518744
rect 452566 518800 452622 518809
rect 452566 518735 452568 518744
rect 443184 518706 443236 518712
rect 429290 518664 429346 518673
rect 429290 518599 429346 518608
rect 432512 518628 432564 518634
rect 426438 518528 426494 518537
rect 426438 518463 426494 518472
rect 426452 518430 426480 518463
rect 426440 518424 426492 518430
rect 426440 518366 426492 518372
rect 429304 518294 429332 518599
rect 432512 518570 432564 518576
rect 430578 518392 430634 518401
rect 432524 518362 432552 518570
rect 430578 518327 430580 518336
rect 430632 518327 430634 518336
rect 432512 518356 432564 518362
rect 430580 518298 430632 518304
rect 432512 518298 432564 518304
rect 429292 518288 429344 518294
rect 429198 518256 429254 518265
rect 429292 518230 429344 518236
rect 432604 518288 432656 518294
rect 432604 518230 432656 518236
rect 429198 518191 429254 518200
rect 429212 518158 429240 518191
rect 429200 518152 429252 518158
rect 429200 518094 429252 518100
rect 425612 518084 425664 518090
rect 425612 518026 425664 518032
rect 431960 518016 432012 518022
rect 431960 517958 432012 517964
rect 428832 482996 428884 483002
rect 428832 482938 428884 482944
rect 426164 482928 426216 482934
rect 426164 482870 426216 482876
rect 424416 482588 424468 482594
rect 424416 482530 424468 482536
rect 420000 482520 420052 482526
rect 420000 482462 420052 482468
rect 417792 482384 417844 482390
rect 417792 482326 417844 482332
rect 412824 482316 412876 482322
rect 412824 482258 412876 482264
rect 415216 482316 415268 482322
rect 415216 482258 415268 482264
rect 398748 479868 398800 479874
rect 369952 479810 370004 479816
rect 399588 479862 399924 479890
rect 401796 479862 402132 479890
rect 404004 479862 404340 479890
rect 406212 479862 406548 479890
rect 408512 479862 408756 479890
rect 410964 479862 411208 479890
rect 412836 479890 412864 482258
rect 412836 479862 413172 479890
rect 398748 479810 398800 479816
rect 362222 479768 362278 479777
rect 344296 479726 344908 479754
rect 362222 479703 362278 479712
rect 367098 479768 367154 479777
rect 367098 479703 367154 479712
rect 316774 479632 316830 479641
rect 367112 479618 367140 479703
rect 367204 479618 367232 479810
rect 415228 479754 415256 482258
rect 417804 479890 417832 482326
rect 420012 479890 420040 482462
rect 422208 482452 422260 482458
rect 422208 482394 422260 482400
rect 422220 479890 422248 482394
rect 424428 479890 424456 482530
rect 417588 479862 417832 479890
rect 419704 479862 420040 479890
rect 421912 479862 422248 479890
rect 424120 479862 424456 479890
rect 415228 479726 415380 479754
rect 367112 479590 367232 479618
rect 426176 479618 426204 482870
rect 428844 479890 428872 482938
rect 431040 482248 431092 482254
rect 431040 482190 431092 482196
rect 431052 479890 431080 482190
rect 428536 479862 428872 479890
rect 430744 479862 431080 479890
rect 431972 479754 432000 517958
rect 432616 517857 432644 518230
rect 435362 518120 435418 518129
rect 435362 518055 435418 518064
rect 435914 518120 435970 518129
rect 435914 518055 435916 518064
rect 433904 517886 433932 517917
rect 433892 517880 433944 517886
rect 432602 517848 432658 517857
rect 432602 517783 432658 517792
rect 433890 517848 433892 517857
rect 433944 517848 433946 517857
rect 433890 517783 433946 517792
rect 432616 482322 432644 517783
rect 433246 517712 433302 517721
rect 433246 517647 433302 517656
rect 433260 482866 433288 517647
rect 433904 511970 433932 517783
rect 434626 517712 434682 517721
rect 434626 517647 434682 517656
rect 433800 511964 433852 511970
rect 433800 511906 433852 511912
rect 433892 511964 433944 511970
rect 433892 511906 433944 511912
rect 433812 502382 433840 511906
rect 433800 502376 433852 502382
rect 433800 502318 433852 502324
rect 434076 502376 434128 502382
rect 434076 502318 434128 502324
rect 434088 495394 434116 502318
rect 433904 495366 434116 495394
rect 433904 492658 433932 495366
rect 433616 492652 433668 492658
rect 433616 492594 433668 492600
rect 433892 492652 433944 492658
rect 433892 492594 433944 492600
rect 433628 483041 433656 492594
rect 433614 483032 433670 483041
rect 433614 482967 433670 482976
rect 433798 483032 433854 483041
rect 433798 482967 433854 482976
rect 433248 482860 433300 482866
rect 433248 482802 433300 482808
rect 433812 482390 433840 482967
rect 434640 482798 434668 517647
rect 434720 517608 434772 517614
rect 434720 517550 434772 517556
rect 434628 482792 434680 482798
rect 434628 482734 434680 482740
rect 433800 482384 433852 482390
rect 433800 482326 433852 482332
rect 432604 482316 432656 482322
rect 432604 482258 432656 482264
rect 434732 479890 434760 517550
rect 435376 482526 435404 518055
rect 435968 518055 435970 518064
rect 435916 518026 435968 518032
rect 437294 517984 437350 517993
rect 436100 517948 436152 517954
rect 436100 517890 436152 517896
rect 436744 517948 436796 517954
rect 437294 517919 437296 517928
rect 436744 517890 436796 517896
rect 437348 517919 437350 517928
rect 437296 517890 437348 517896
rect 436006 517712 436062 517721
rect 436006 517647 436062 517656
rect 436020 482730 436048 517647
rect 436008 482724 436060 482730
rect 436008 482666 436060 482672
rect 435364 482520 435416 482526
rect 435364 482462 435416 482468
rect 436112 480298 436140 517890
rect 436650 517712 436706 517721
rect 436650 517647 436706 517656
rect 436664 517614 436692 517647
rect 436652 517608 436704 517614
rect 436652 517550 436704 517556
rect 436756 482594 436784 517890
rect 440882 517848 440938 517857
rect 438124 517812 438176 517818
rect 440882 517783 440938 517792
rect 438124 517754 438176 517760
rect 437386 517712 437442 517721
rect 437386 517647 437442 517656
rect 436928 517608 436980 517614
rect 436928 517550 436980 517556
rect 436744 482588 436796 482594
rect 436744 482530 436796 482536
rect 436940 482458 436968 517550
rect 437400 482662 437428 517647
rect 438136 517585 438164 517754
rect 440896 517750 440924 517783
rect 440884 517744 440936 517750
rect 438674 517712 438730 517721
rect 439502 517712 439558 517721
rect 438674 517647 438730 517656
rect 438860 517676 438912 517682
rect 438122 517576 438178 517585
rect 438122 517511 438178 517520
rect 438136 482934 438164 517511
rect 438124 482928 438176 482934
rect 438124 482870 438176 482876
rect 437388 482656 437440 482662
rect 437388 482598 437440 482604
rect 438688 482594 438716 517647
rect 440884 517686 440936 517692
rect 439502 517647 439504 517656
rect 438860 517618 438912 517624
rect 439556 517647 439558 517656
rect 439504 517618 439556 517624
rect 438766 517576 438822 517585
rect 438766 517511 438822 517520
rect 438676 482588 438728 482594
rect 438676 482530 438728 482536
rect 438780 482526 438808 517511
rect 438768 482520 438820 482526
rect 438768 482462 438820 482468
rect 436928 482452 436980 482458
rect 436928 482394 436980 482400
rect 436112 480270 436968 480298
rect 436940 479890 436968 480270
rect 434732 479862 435160 479890
rect 436940 479862 437368 479890
rect 438872 479754 438900 517618
rect 439516 483002 439544 517618
rect 440146 517576 440202 517585
rect 440146 517511 440202 517520
rect 439504 482996 439556 483002
rect 439504 482938 439556 482944
rect 440160 482458 440188 517511
rect 440148 482452 440200 482458
rect 440148 482394 440200 482400
rect 440896 482254 440924 517686
rect 441526 517576 441582 517585
rect 441526 517511 441582 517520
rect 441540 482390 441568 517511
rect 441528 482384 441580 482390
rect 441528 482326 441580 482332
rect 440884 482248 440936 482254
rect 440884 482190 440936 482196
rect 441632 479890 441660 518706
rect 443000 518696 443052 518702
rect 443000 518638 443052 518644
rect 442078 518392 442134 518401
rect 442078 518327 442134 518336
rect 442092 518294 442120 518327
rect 442080 518288 442132 518294
rect 442080 518230 442132 518236
rect 442906 517576 442962 517585
rect 442906 517511 442962 517520
rect 442920 482322 442948 517511
rect 442908 482316 442960 482322
rect 442908 482258 442960 482264
rect 443012 480026 443040 518638
rect 443196 517886 443224 518706
rect 446588 518628 446640 518634
rect 446588 518570 446640 518576
rect 445760 518560 445812 518566
rect 445390 518528 445446 518537
rect 446600 518537 446628 518570
rect 447428 518566 447456 518597
rect 447416 518560 447468 518566
rect 445760 518502 445812 518508
rect 446586 518528 446642 518537
rect 445390 518463 445446 518472
rect 445404 518430 445432 518463
rect 445392 518424 445444 518430
rect 444286 518392 444342 518401
rect 445392 518366 445444 518372
rect 444286 518327 444342 518336
rect 444300 518294 444328 518327
rect 444288 518288 444340 518294
rect 444288 518230 444340 518236
rect 444300 518090 444328 518230
rect 444288 518084 444340 518090
rect 444288 518026 444340 518032
rect 443184 517880 443236 517886
rect 443184 517822 443236 517828
rect 445404 517614 445432 518366
rect 445666 517712 445722 517721
rect 445666 517647 445722 517656
rect 445392 517608 445444 517614
rect 444286 517576 444342 517585
rect 445392 517550 445444 517556
rect 445574 517576 445630 517585
rect 444286 517511 444342 517520
rect 445574 517511 445630 517520
rect 444300 481710 444328 517511
rect 445588 481914 445616 517511
rect 445576 481908 445628 481914
rect 445576 481850 445628 481856
rect 445680 481778 445708 517647
rect 445668 481772 445720 481778
rect 445668 481714 445720 481720
rect 444288 481704 444340 481710
rect 444288 481646 444340 481652
rect 443012 479998 443500 480026
rect 441632 479862 441784 479890
rect 443472 479754 443500 479998
rect 445772 479890 445800 518502
rect 446586 518463 446642 518472
rect 447414 518528 447416 518537
rect 447468 518528 447470 518537
rect 447414 518463 447470 518472
rect 448796 518492 448848 518498
rect 446600 517954 446628 518463
rect 447140 518356 447192 518362
rect 447140 518298 447192 518304
rect 446588 517948 446640 517954
rect 446588 517890 446640 517896
rect 447046 517576 447102 517585
rect 447046 517511 447102 517520
rect 447060 481846 447088 517511
rect 447048 481840 447100 481846
rect 447048 481782 447100 481788
rect 447152 480026 447180 518298
rect 447428 517818 447456 518463
rect 448796 518434 448848 518440
rect 448808 518401 448836 518434
rect 448794 518392 448850 518401
rect 448794 518327 448850 518336
rect 449898 518392 449954 518401
rect 449898 518327 449900 518336
rect 447416 517812 447468 517818
rect 447416 517754 447468 517760
rect 448808 517682 448836 518327
rect 449952 518327 449954 518336
rect 449900 518298 449952 518304
rect 449912 517750 449940 518298
rect 451292 518226 451320 518735
rect 452620 518735 452622 518744
rect 453670 518800 453726 518809
rect 453670 518735 453726 518744
rect 459558 518800 459560 518809
rect 459612 518800 459614 518809
rect 459558 518735 459614 518744
rect 460938 518800 460994 518809
rect 460938 518735 460940 518744
rect 452568 518706 452620 518712
rect 453684 518702 453712 518735
rect 460992 518735 460994 518744
rect 462318 518800 462374 518809
rect 462318 518735 462374 518744
rect 460940 518706 460992 518712
rect 462332 518702 462360 518735
rect 453672 518696 453724 518702
rect 462320 518696 462372 518702
rect 453672 518638 453724 518644
rect 455326 518664 455382 518673
rect 453684 518294 453712 518638
rect 455326 518599 455382 518608
rect 456062 518664 456118 518673
rect 456062 518599 456064 518608
rect 455340 518430 455368 518599
rect 456116 518599 456118 518608
rect 456890 518664 456946 518673
rect 456890 518599 456946 518608
rect 458270 518664 458326 518673
rect 458270 518599 458326 518608
rect 459558 518664 459614 518673
rect 462320 518638 462372 518644
rect 465078 518664 465134 518673
rect 459558 518599 459614 518608
rect 465078 518599 465080 518608
rect 456064 518570 456116 518576
rect 456904 518566 456932 518599
rect 456892 518560 456944 518566
rect 456892 518502 456944 518508
rect 456904 518430 456932 518502
rect 458284 518498 458312 518599
rect 458272 518492 458324 518498
rect 458272 518434 458324 518440
rect 455328 518424 455380 518430
rect 455328 518366 455380 518372
rect 456892 518424 456944 518430
rect 456892 518366 456944 518372
rect 455340 518294 455368 518366
rect 459572 518362 459600 518599
rect 465132 518599 465134 518608
rect 466550 518664 466606 518673
rect 466550 518599 466606 518608
rect 465080 518570 465132 518576
rect 466458 518528 466514 518537
rect 466564 518498 466592 518599
rect 466458 518463 466514 518472
rect 466552 518492 466604 518498
rect 466472 518430 466500 518463
rect 466552 518434 466604 518440
rect 466460 518424 466512 518430
rect 463698 518392 463754 518401
rect 459560 518356 459612 518362
rect 466460 518366 466512 518372
rect 467838 518392 467894 518401
rect 463698 518327 463754 518336
rect 467838 518327 467840 518336
rect 459560 518298 459612 518304
rect 463712 518294 463740 518327
rect 467892 518327 467894 518336
rect 467840 518298 467892 518304
rect 453672 518288 453724 518294
rect 453672 518230 453724 518236
rect 455328 518288 455380 518294
rect 455328 518230 455380 518236
rect 463700 518288 463752 518294
rect 463700 518230 463752 518236
rect 451280 518220 451332 518226
rect 451280 518162 451332 518168
rect 449900 517744 449952 517750
rect 449900 517686 449952 517692
rect 453946 517712 454002 517721
rect 448796 517676 448848 517682
rect 453946 517647 454002 517656
rect 460846 517712 460902 517721
rect 460846 517647 460902 517656
rect 469126 517712 469182 517721
rect 469126 517647 469182 517656
rect 448796 517618 448848 517624
rect 448426 517576 448482 517585
rect 448426 517511 448482 517520
rect 449806 517576 449862 517585
rect 449806 517511 449862 517520
rect 451186 517576 451242 517585
rect 451186 517511 451242 517520
rect 452566 517576 452622 517585
rect 452566 517511 452622 517520
rect 453854 517576 453910 517585
rect 453854 517511 453910 517520
rect 448440 482050 448468 517511
rect 448428 482044 448480 482050
rect 448428 481986 448480 481992
rect 449820 481982 449848 517511
rect 450268 482860 450320 482866
rect 450268 482802 450320 482808
rect 449808 481976 449860 481982
rect 449808 481918 449860 481924
rect 447152 479998 447824 480026
rect 447796 479890 447824 479998
rect 450280 479890 450308 482802
rect 451200 482118 451228 517511
rect 452580 482186 452608 517511
rect 453868 482934 453896 517511
rect 453856 482928 453908 482934
rect 453856 482870 453908 482876
rect 452660 482792 452712 482798
rect 452660 482734 452712 482740
rect 452568 482180 452620 482186
rect 452568 482122 452620 482128
rect 451188 482112 451240 482118
rect 451188 482054 451240 482060
rect 452672 480162 452700 482734
rect 453960 482254 453988 517647
rect 455326 517576 455382 517585
rect 455326 517511 455382 517520
rect 456706 517576 456762 517585
rect 456706 517511 456762 517520
rect 458086 517576 458142 517585
rect 458086 517511 458142 517520
rect 459466 517576 459522 517585
rect 459466 517511 459522 517520
rect 460754 517576 460810 517585
rect 460754 517511 460810 517520
rect 455340 483002 455368 517511
rect 455328 482996 455380 483002
rect 455328 482938 455380 482944
rect 456720 482798 456748 517511
rect 458100 482866 458128 517511
rect 458088 482860 458140 482866
rect 458088 482802 458140 482808
rect 456708 482792 456760 482798
rect 456708 482734 456760 482740
rect 459480 482730 459508 517511
rect 454592 482724 454644 482730
rect 454592 482666 454644 482672
rect 459468 482724 459520 482730
rect 459468 482666 459520 482672
rect 453948 482248 454000 482254
rect 453948 482190 454000 482196
rect 452672 480134 452746 480162
rect 445772 479862 446200 479890
rect 447796 479862 448408 479890
rect 450280 479862 450616 479890
rect 452718 479876 452746 480134
rect 454604 479890 454632 482666
rect 456892 482656 456944 482662
rect 456892 482598 456944 482604
rect 456904 479890 456932 482598
rect 460768 482594 460796 517511
rect 460860 482662 460888 517647
rect 462226 517576 462282 517585
rect 462226 517511 462282 517520
rect 463606 517576 463662 517585
rect 463606 517511 463662 517520
rect 464986 517576 465042 517585
rect 464986 517511 465042 517520
rect 466366 517576 466422 517585
rect 466366 517511 466422 517520
rect 467746 517576 467802 517585
rect 467746 517511 467802 517520
rect 469034 517576 469090 517585
rect 469034 517511 469090 517520
rect 460848 482656 460900 482662
rect 460848 482598 460900 482604
rect 459008 482588 459060 482594
rect 459008 482530 459060 482536
rect 460756 482588 460808 482594
rect 460756 482530 460808 482536
rect 459020 479890 459048 482530
rect 462240 482526 462268 517511
rect 461216 482520 461268 482526
rect 461216 482462 461268 482468
rect 462228 482520 462280 482526
rect 463620 482497 463648 517511
rect 462228 482462 462280 482468
rect 463606 482488 463662 482497
rect 461228 479890 461256 482462
rect 465000 482458 465028 517511
rect 463606 482423 463662 482432
rect 463700 482452 463752 482458
rect 463700 482394 463752 482400
rect 464988 482452 465040 482458
rect 464988 482394 465040 482400
rect 463712 480162 463740 482394
rect 466380 482390 466408 517511
rect 465632 482384 465684 482390
rect 465632 482326 465684 482332
rect 466368 482384 466420 482390
rect 467760 482361 467788 517511
rect 466368 482326 466420 482332
rect 467746 482352 467802 482361
rect 463712 480134 463786 480162
rect 454604 479862 454940 479890
rect 456904 479862 457148 479890
rect 459020 479862 459356 479890
rect 461228 479862 461564 479890
rect 463758 479876 463786 480134
rect 465644 479890 465672 482326
rect 467746 482287 467802 482296
rect 467840 482316 467892 482322
rect 467840 482258 467892 482264
rect 467852 479890 467880 482258
rect 469048 482225 469076 517511
rect 469140 482322 469168 517647
rect 492036 482996 492088 483002
rect 492036 482938 492088 482944
rect 489920 482928 489972 482934
rect 489920 482870 489972 482876
rect 469128 482316 469180 482322
rect 469128 482258 469180 482264
rect 487620 482248 487672 482254
rect 469034 482216 469090 482225
rect 487620 482190 487672 482196
rect 469034 482151 469090 482160
rect 485780 482180 485832 482186
rect 485780 482122 485832 482128
rect 483296 482112 483348 482118
rect 483296 482054 483348 482060
rect 478880 482044 478932 482050
rect 478880 481986 478932 481992
rect 474740 481908 474792 481914
rect 474740 481850 474792 481856
rect 472256 481772 472308 481778
rect 472256 481714 472308 481720
rect 470048 481704 470100 481710
rect 470048 481646 470100 481652
rect 470060 479890 470088 481646
rect 472268 479890 472296 481714
rect 474752 480162 474780 481850
rect 476672 481840 476724 481846
rect 476672 481782 476724 481788
rect 474752 480134 474826 480162
rect 465644 479862 465980 479890
rect 467852 479862 468188 479890
rect 470060 479862 470396 479890
rect 472268 479862 472604 479890
rect 474798 479876 474826 480134
rect 476684 479890 476712 481782
rect 478892 479890 478920 481986
rect 481088 481976 481140 481982
rect 481088 481918 481140 481924
rect 481100 479890 481128 481918
rect 483308 479890 483336 482054
rect 485792 480162 485820 482122
rect 485792 480134 485866 480162
rect 476684 479862 477020 479890
rect 478892 479862 479228 479890
rect 481100 479862 481436 479890
rect 483308 479862 483644 479890
rect 485838 479876 485866 480134
rect 487632 479890 487660 482190
rect 489932 479890 489960 482870
rect 492048 479890 492076 482938
rect 496452 482860 496504 482866
rect 496452 482802 496504 482808
rect 494244 482792 494296 482798
rect 494244 482734 494296 482740
rect 494256 479890 494284 482734
rect 496464 479890 496492 482802
rect 498660 482724 498712 482730
rect 498660 482666 498712 482672
rect 498672 479890 498700 482666
rect 500960 482656 501012 482662
rect 500960 482598 501012 482604
rect 500972 479890 501000 482598
rect 503076 482588 503128 482594
rect 503076 482530 503128 482536
rect 503088 479890 503116 482530
rect 505284 482520 505336 482526
rect 505284 482462 505336 482468
rect 507490 482488 507546 482497
rect 505296 479890 505324 482462
rect 507490 482423 507546 482432
rect 509700 482452 509752 482458
rect 507504 479890 507532 482423
rect 509700 482394 509752 482400
rect 509712 479890 509740 482394
rect 512000 482384 512052 482390
rect 512000 482326 512052 482332
rect 514114 482352 514170 482361
rect 512012 479890 512040 482326
rect 514114 482287 514170 482296
rect 516324 482316 516376 482322
rect 514128 479890 514156 482287
rect 516324 482258 516376 482264
rect 516336 479890 516364 482258
rect 518530 482216 518586 482225
rect 518530 482151 518586 482160
rect 518544 479890 518572 482151
rect 487632 479862 487968 479890
rect 489932 479862 490176 479890
rect 492048 479862 492384 479890
rect 494256 479862 494592 479890
rect 496464 479862 496800 479890
rect 498672 479862 499008 479890
rect 500972 479862 501216 479890
rect 503088 479862 503424 479890
rect 505296 479862 505632 479890
rect 507504 479862 507840 479890
rect 509712 479862 510048 479890
rect 512012 479862 512256 479890
rect 514128 479862 514464 479890
rect 516336 479862 516672 479890
rect 518544 479862 518880 479890
rect 444286 479768 444342 479777
rect 431972 479726 432952 479754
rect 438872 479726 439576 479754
rect 443472 479726 443992 479754
rect 444286 479703 444342 479712
rect 426176 479590 426328 479618
rect 316774 479567 316830 479576
rect 283562 479496 283618 479505
rect 283562 479431 283564 479440
rect 283616 479431 283618 479440
rect 283564 479402 283616 479408
rect 309138 479360 309194 479369
rect 316788 479330 316816 479567
rect 444300 479505 444328 479703
rect 466366 479632 466422 479641
rect 466366 479567 466422 479576
rect 507122 479632 507178 479641
rect 507122 479567 507178 479576
rect 427818 479496 427874 479505
rect 427740 479454 427818 479482
rect 427740 479369 427768 479454
rect 427818 479431 427874 479440
rect 444286 479496 444342 479505
rect 466380 479466 466408 479567
rect 473266 479496 473322 479505
rect 444286 479431 444342 479440
rect 466368 479460 466420 479466
rect 473266 479431 473268 479440
rect 466368 479402 466420 479408
rect 473320 479431 473322 479440
rect 492586 479496 492642 479505
rect 492586 479431 492642 479440
rect 473268 479402 473320 479408
rect 492600 479398 492628 479431
rect 485688 479392 485740 479398
rect 321374 479360 321430 479369
rect 309138 479295 309140 479304
rect 309192 479295 309194 479304
rect 316776 479324 316828 479330
rect 309140 479266 309192 479272
rect 321558 479360 321614 479369
rect 321430 479318 321558 479346
rect 321374 479295 321430 479304
rect 321558 479295 321614 479304
rect 350446 479360 350502 479369
rect 350630 479360 350686 479369
rect 350502 479318 350630 479346
rect 350446 479295 350502 479304
rect 350630 479295 350686 479304
rect 427726 479360 427782 479369
rect 427726 479295 427782 479304
rect 485686 479360 485688 479369
rect 492588 479392 492640 479398
rect 485740 479360 485742 479369
rect 507136 479369 507164 479567
rect 492588 479334 492640 479340
rect 507122 479360 507178 479369
rect 485686 479295 485742 479304
rect 507122 479295 507178 479304
rect 316776 479266 316828 479272
rect 519096 346474 519124 700810
rect 519176 700800 519228 700806
rect 519176 700742 519228 700748
rect 519188 353002 519216 700742
rect 520280 700732 520332 700738
rect 520280 700674 520332 700680
rect 519268 700596 519320 700602
rect 519268 700538 519320 700544
rect 519280 363474 519308 700538
rect 519452 700528 519504 700534
rect 519452 700470 519504 700476
rect 519360 700460 519412 700466
rect 519360 700402 519412 700408
rect 519372 369753 519400 700402
rect 519464 372065 519492 700470
rect 519544 700324 519596 700330
rect 519544 700266 519596 700272
rect 519556 376281 519584 700266
rect 519634 695328 519690 695337
rect 519634 695263 519690 695272
rect 519648 686089 519676 695263
rect 519634 686080 519690 686089
rect 519634 686015 519690 686024
rect 519910 684312 519966 684321
rect 519910 684247 519966 684256
rect 519924 666641 519952 684247
rect 519910 666632 519966 666641
rect 519910 666567 519966 666576
rect 519636 610836 519688 610842
rect 519636 610778 519688 610784
rect 519542 376272 519598 376281
rect 519542 376207 519598 376216
rect 519450 372056 519506 372065
rect 519450 371991 519506 372000
rect 519358 369744 519414 369753
rect 519358 369679 519414 369688
rect 519358 363488 519414 363497
rect 519280 363446 519358 363474
rect 519358 363423 519414 363432
rect 519358 353016 519414 353025
rect 519188 352974 519358 353002
rect 519358 352951 519414 352960
rect 519266 346488 519322 346497
rect 519096 346446 519266 346474
rect 519266 346423 519322 346432
rect 519648 344593 519676 610778
rect 519728 610632 519780 610638
rect 519728 610574 519780 610580
rect 519740 357377 519768 610574
rect 520004 509312 520056 509318
rect 520004 509254 520056 509260
rect 519912 479188 519964 479194
rect 519912 479130 519964 479136
rect 519818 479088 519874 479097
rect 519818 479023 519874 479032
rect 519832 478922 519860 479023
rect 519820 478916 519872 478922
rect 519820 478858 519872 478864
rect 519924 478802 519952 479130
rect 519832 478774 519952 478802
rect 519832 437617 519860 478774
rect 519912 478712 519964 478718
rect 519912 478654 519964 478660
rect 519818 437608 519874 437617
rect 519818 437543 519874 437552
rect 519820 437504 519872 437510
rect 519820 437446 519872 437452
rect 519726 357368 519782 357377
rect 519726 357303 519782 357312
rect 519634 344584 519690 344593
rect 519634 344519 519690 344528
rect 519832 240854 519860 437446
rect 519924 351121 519952 478654
rect 520016 412185 520044 509254
rect 520188 480276 520240 480282
rect 520188 480218 520240 480224
rect 520096 479868 520148 479874
rect 520096 479810 520148 479816
rect 520108 478786 520136 479810
rect 520096 478780 520148 478786
rect 520096 478722 520148 478728
rect 520200 478666 520228 480218
rect 520108 478638 520228 478666
rect 520108 476241 520136 478638
rect 520188 478576 520240 478582
rect 520188 478518 520240 478524
rect 520094 476232 520150 476241
rect 520094 476167 520150 476176
rect 520094 476096 520150 476105
rect 520094 476031 520150 476040
rect 520108 413681 520136 476031
rect 520200 417897 520228 478518
rect 520186 417888 520242 417897
rect 520186 417823 520242 417832
rect 520186 414896 520242 414905
rect 520186 414831 520242 414840
rect 520094 413672 520150 413681
rect 520094 413607 520150 413616
rect 520002 412176 520058 412185
rect 520002 412111 520058 412120
rect 520002 409184 520058 409193
rect 520002 409119 520058 409128
rect 520016 406065 520044 409119
rect 520200 406201 520228 414831
rect 520186 406192 520242 406201
rect 520186 406127 520242 406136
rect 520002 406056 520058 406065
rect 520002 405991 520058 406000
rect 520002 396400 520058 396409
rect 520002 396335 520058 396344
rect 520016 393145 520044 396335
rect 520094 395584 520150 395593
rect 520094 395519 520150 395528
rect 520002 393136 520058 393145
rect 520002 393071 520058 393080
rect 520108 390697 520136 395519
rect 520094 390688 520150 390697
rect 520094 390623 520150 390632
rect 520292 359009 520320 700674
rect 520372 700664 520424 700670
rect 520372 700606 520424 700612
rect 520384 365265 520412 700606
rect 520464 700392 520516 700398
rect 520464 700334 520516 700340
rect 520476 377913 520504 700334
rect 525064 626612 525116 626618
rect 525064 626554 525116 626560
rect 520556 610904 520608 610910
rect 520556 610846 520608 610852
rect 520462 377904 520518 377913
rect 520462 377839 520518 377848
rect 520370 365256 520426 365265
rect 520370 365191 520426 365200
rect 520278 359000 520334 359009
rect 520278 358935 520334 358944
rect 519910 351112 519966 351121
rect 519910 351047 519966 351056
rect 520568 342145 520596 610846
rect 520648 610768 520700 610774
rect 520648 610710 520700 610716
rect 520660 348401 520688 610710
rect 520740 610700 520792 610706
rect 520740 610642 520792 610648
rect 520752 354793 520780 610642
rect 520832 610360 520884 610366
rect 520832 610302 520884 610308
rect 520844 403209 520872 610302
rect 523684 579692 523736 579698
rect 523684 579634 523736 579640
rect 521292 495508 521344 495514
rect 521292 495450 521344 495456
rect 520924 479800 520976 479806
rect 520924 479742 520976 479748
rect 520830 403200 520886 403209
rect 520830 403135 520886 403144
rect 520936 361049 520964 479742
rect 521016 479732 521068 479738
rect 521016 479674 521068 479680
rect 521028 367305 521056 479674
rect 521108 479664 521160 479670
rect 521108 479606 521160 479612
rect 521120 373697 521148 479606
rect 521200 479596 521252 479602
rect 521200 479538 521252 479544
rect 521212 379953 521240 479538
rect 521304 415857 521332 495450
rect 521384 479528 521436 479534
rect 521384 479470 521436 479476
rect 521290 415848 521346 415857
rect 521290 415783 521346 415792
rect 521396 405249 521424 479470
rect 521568 479120 521620 479126
rect 521568 479062 521620 479068
rect 521476 478508 521528 478514
rect 521476 478450 521528 478456
rect 521488 424153 521516 478450
rect 521580 432585 521608 479062
rect 523132 479052 523184 479058
rect 523132 478994 523184 479000
rect 523040 478984 523092 478990
rect 523040 478926 523092 478932
rect 522672 478440 522724 478446
rect 522672 478382 522724 478388
rect 522488 478304 522540 478310
rect 522488 478246 522540 478252
rect 522304 478236 522356 478242
rect 522304 478178 522356 478184
rect 521658 460048 521714 460057
rect 521658 459983 521714 459992
rect 521566 432576 521622 432585
rect 521566 432511 521622 432520
rect 521474 424144 521530 424153
rect 521474 424079 521530 424088
rect 521382 405240 521438 405249
rect 521382 405175 521438 405184
rect 521198 379944 521254 379953
rect 521198 379879 521254 379888
rect 521106 373688 521162 373697
rect 521106 373623 521162 373632
rect 521014 367296 521070 367305
rect 521014 367231 521070 367240
rect 520922 361040 520978 361049
rect 520922 360975 520978 360984
rect 520738 354784 520794 354793
rect 520738 354719 520794 354728
rect 520646 348392 520702 348401
rect 520646 348327 520702 348336
rect 520554 342136 520610 342145
rect 520554 342071 520610 342080
rect 519820 240848 519872 240854
rect 519820 240790 519872 240796
rect 280160 240712 280212 240718
rect 280160 240654 280212 240660
rect 280896 240712 280948 240718
rect 280896 240654 280948 240660
rect 306380 240712 306432 240718
rect 306380 240654 306432 240660
rect 315948 240712 316000 240718
rect 325608 240712 325660 240718
rect 315948 240654 316000 240660
rect 316038 240680 316094 240689
rect 306392 240514 306420 240654
rect 315960 240514 315988 240654
rect 316038 240615 316040 240624
rect 316092 240615 316094 240624
rect 325606 240680 325608 240689
rect 340880 240712 340932 240718
rect 325660 240680 325662 240689
rect 340800 240660 340880 240666
rect 340800 240654 340932 240660
rect 350448 240712 350500 240718
rect 369676 240712 369728 240718
rect 357438 240680 357494 240689
rect 350500 240660 350672 240666
rect 350448 240654 350672 240660
rect 340800 240650 340920 240654
rect 325606 240615 325662 240624
rect 340788 240644 340920 240650
rect 316040 240586 316092 240592
rect 340840 240638 340920 240644
rect 350460 240650 350672 240654
rect 350460 240644 350684 240650
rect 350460 240638 350632 240644
rect 340788 240586 340840 240592
rect 357438 240615 357440 240624
rect 350632 240586 350684 240592
rect 357492 240615 357494 240624
rect 360382 240680 360438 240689
rect 369676 240654 369728 240660
rect 360382 240615 360384 240624
rect 357440 240586 357492 240592
rect 360436 240615 360438 240624
rect 360384 240586 360436 240592
rect 306380 240508 306432 240514
rect 306380 240450 306432 240456
rect 315948 240508 316000 240514
rect 315948 240450 316000 240456
rect 369688 240446 369716 240654
rect 369676 240440 369728 240446
rect 369676 240382 369728 240388
rect 373264 240440 373316 240446
rect 373264 240382 373316 240388
rect 278688 240168 278740 240174
rect 278688 240110 278740 240116
rect 281060 240094 281396 240122
rect 283176 240094 283512 240122
rect 285384 240094 285628 240122
rect 287592 240094 287928 240122
rect 281368 238134 281396 240094
rect 283484 238202 283512 240094
rect 283472 238196 283524 238202
rect 283472 238138 283524 238144
rect 281356 238128 281408 238134
rect 281356 238070 281408 238076
rect 285600 238066 285628 240094
rect 285588 238060 285640 238066
rect 285588 238002 285640 238008
rect 287900 237454 287928 240094
rect 289786 239850 289814 240108
rect 292008 240094 292528 240122
rect 294216 240094 294552 240122
rect 296424 240094 296668 240122
rect 298632 240094 298968 240122
rect 289740 239822 289814 239850
rect 287888 237448 287940 237454
rect 287888 237390 287940 237396
rect 288348 237448 288400 237454
rect 288348 237390 288400 237396
rect 288360 203969 288388 237390
rect 288346 203960 288402 203969
rect 288346 203895 288402 203904
rect 289740 203833 289768 239822
rect 292500 204105 292528 240094
rect 294524 238474 294552 240094
rect 294512 238468 294564 238474
rect 294512 238410 294564 238416
rect 295248 238468 295300 238474
rect 295248 238410 295300 238416
rect 292486 204096 292542 204105
rect 292486 204031 292542 204040
rect 289726 203824 289782 203833
rect 289726 203759 289782 203768
rect 295260 202910 295288 238410
rect 296640 203046 296668 240094
rect 297824 238196 297876 238202
rect 297824 238138 297876 238144
rect 297364 238128 297416 238134
rect 297364 238070 297416 238076
rect 296628 203040 296680 203046
rect 296628 202982 296680 202988
rect 295248 202904 295300 202910
rect 295248 202846 295300 202852
rect 297376 202842 297404 238070
rect 297364 202836 297416 202842
rect 297364 202778 297416 202784
rect 297836 111761 297864 238138
rect 298940 237454 298968 240094
rect 300826 239850 300854 240108
rect 303048 240094 303384 240122
rect 305256 240094 305592 240122
rect 307464 240094 307708 240122
rect 309672 240094 310008 240122
rect 300780 239822 300854 239850
rect 298928 237448 298980 237454
rect 298928 237390 298980 237396
rect 299388 237448 299440 237454
rect 299388 237390 299440 237396
rect 299400 204202 299428 237390
rect 299388 204196 299440 204202
rect 299388 204138 299440 204144
rect 300780 204066 300808 239822
rect 303356 238202 303384 240094
rect 305564 238270 305592 240094
rect 305552 238264 305604 238270
rect 305552 238206 305604 238212
rect 303344 238196 303396 238202
rect 303344 238138 303396 238144
rect 307680 238134 307708 240094
rect 309980 238338 310008 240094
rect 311866 239850 311894 240108
rect 314088 240094 314608 240122
rect 316204 240094 316540 240122
rect 318412 240094 318748 240122
rect 320620 240094 320956 240122
rect 311820 239822 311894 239850
rect 311820 238406 311848 239822
rect 311808 238400 311860 238406
rect 311808 238342 311860 238348
rect 309968 238332 310020 238338
rect 309968 238274 310020 238280
rect 307668 238128 307720 238134
rect 307668 238070 307720 238076
rect 300768 204060 300820 204066
rect 300768 204002 300820 204008
rect 314580 203998 314608 240094
rect 316512 237454 316540 240094
rect 316500 237448 316552 237454
rect 316500 237390 316552 237396
rect 317328 237448 317380 237454
rect 317328 237390 317380 237396
rect 317340 204270 317368 237390
rect 317328 204264 317380 204270
rect 317328 204206 317380 204212
rect 314568 203992 314620 203998
rect 314568 203934 314620 203940
rect 318720 203862 318748 240094
rect 320928 237454 320956 240094
rect 322814 239850 322842 240108
rect 325036 240094 325648 240122
rect 327244 240094 327580 240122
rect 329452 240094 329788 240122
rect 331660 240094 331996 240122
rect 322814 239822 322888 239850
rect 320916 237448 320968 237454
rect 320916 237390 320968 237396
rect 321468 237448 321520 237454
rect 321468 237390 321520 237396
rect 318708 203856 318760 203862
rect 318708 203798 318760 203804
rect 321480 203794 321508 237390
rect 321468 203788 321520 203794
rect 321468 203730 321520 203736
rect 322860 203726 322888 239822
rect 322848 203720 322900 203726
rect 322848 203662 322900 203668
rect 325620 203658 325648 240094
rect 327552 237454 327580 240094
rect 329564 238536 329616 238542
rect 329564 238478 329616 238484
rect 328368 238468 328420 238474
rect 328368 238410 328420 238416
rect 327540 237448 327592 237454
rect 327540 237390 327592 237396
rect 328276 237448 328328 237454
rect 328276 237390 328328 237396
rect 325608 203652 325660 203658
rect 325608 203594 325660 203600
rect 328288 203590 328316 237390
rect 328276 203584 328328 203590
rect 328276 203526 328328 203532
rect 328276 203380 328328 203386
rect 328276 203322 328328 203328
rect 328288 203153 328316 203322
rect 328380 203289 328408 238410
rect 329576 234598 329604 238478
rect 329760 237454 329788 240094
rect 331128 238604 331180 238610
rect 331128 238546 331180 238552
rect 329748 237448 329800 237454
rect 329748 237390 329800 237396
rect 329564 234592 329616 234598
rect 329564 234534 329616 234540
rect 329748 234592 329800 234598
rect 329748 234534 329800 234540
rect 329760 231826 329788 234534
rect 329668 231798 329788 231826
rect 329668 222222 329696 231798
rect 329472 222216 329524 222222
rect 329472 222158 329524 222164
rect 329656 222216 329708 222222
rect 329656 222158 329708 222164
rect 329484 215370 329512 222158
rect 329392 215342 329512 215370
rect 329392 212537 329420 215342
rect 329378 212528 329434 212537
rect 329378 212463 329434 212472
rect 330944 204128 330996 204134
rect 330944 204070 330996 204076
rect 330956 203697 330984 204070
rect 330942 203688 330998 203697
rect 330942 203623 330998 203632
rect 329748 203448 329800 203454
rect 329746 203416 329748 203425
rect 331140 203425 331168 238546
rect 331968 237726 331996 240094
rect 333854 239850 333882 240108
rect 336076 240094 336688 240122
rect 333854 239822 333928 239850
rect 333704 238740 333756 238746
rect 333704 238682 333756 238688
rect 332508 238672 332560 238678
rect 332508 238614 332560 238620
rect 331956 237720 332008 237726
rect 331956 237662 332008 237668
rect 331220 203652 331272 203658
rect 331220 203594 331272 203600
rect 329800 203416 329802 203425
rect 329746 203351 329802 203360
rect 331126 203416 331182 203425
rect 331126 203351 331182 203360
rect 328366 203280 328422 203289
rect 331232 203250 331260 203594
rect 332416 203312 332468 203318
rect 332520 203289 332548 238614
rect 333716 237454 333744 238682
rect 333900 237590 333928 239822
rect 335176 237856 335228 237862
rect 335176 237798 335228 237804
rect 333888 237584 333940 237590
rect 333888 237526 333940 237532
rect 333704 237448 333756 237454
rect 333704 237390 333756 237396
rect 333888 237448 333940 237454
rect 333888 237390 333940 237396
rect 333796 203924 333848 203930
rect 333796 203866 333848 203872
rect 332416 203254 332468 203260
rect 332506 203280 332562 203289
rect 328366 203215 328422 203224
rect 331220 203244 331272 203250
rect 331220 203186 331272 203192
rect 332428 203153 332456 203254
rect 332506 203215 332562 203224
rect 333808 203153 333836 203866
rect 333900 203289 333928 237390
rect 335084 203856 335136 203862
rect 335084 203798 335136 203804
rect 335096 203522 335124 203798
rect 335084 203516 335136 203522
rect 335084 203458 335136 203464
rect 335188 203425 335216 237798
rect 335268 237652 335320 237658
rect 335268 237594 335320 237600
rect 335174 203416 335230 203425
rect 335174 203351 335230 203360
rect 335280 203289 335308 237594
rect 336556 237448 336608 237454
rect 336556 237390 336608 237396
rect 336660 237402 336688 240094
rect 338132 240094 338284 240122
rect 340156 240094 340492 240122
rect 342364 240094 342700 240122
rect 344572 240094 344908 240122
rect 346780 240094 347116 240122
rect 349172 240094 349324 240122
rect 351104 240094 351440 240122
rect 353312 240094 353648 240122
rect 355856 240094 356008 240122
rect 358064 240094 358768 240122
rect 360272 240094 360608 240122
rect 362480 240094 362908 240122
rect 364688 240094 365024 240122
rect 337384 237516 337436 237522
rect 337384 237458 337436 237464
rect 336568 230518 336596 237390
rect 336660 237374 336780 237402
rect 336372 230512 336424 230518
rect 336372 230454 336424 230460
rect 336556 230512 336608 230518
rect 336556 230454 336608 230460
rect 336384 222290 336412 230454
rect 336372 222284 336424 222290
rect 336372 222226 336424 222232
rect 336648 222284 336700 222290
rect 336648 222226 336700 222232
rect 336660 220833 336688 222226
rect 336646 220824 336702 220833
rect 336646 220759 336702 220768
rect 335820 203788 335872 203794
rect 335820 203730 335872 203736
rect 335832 203386 335860 203730
rect 336004 203720 336056 203726
rect 336004 203662 336056 203668
rect 336016 203454 336044 203662
rect 336004 203448 336056 203454
rect 336752 203425 336780 237374
rect 337396 204134 337424 237458
rect 338132 237454 338160 240094
rect 339592 237720 339644 237726
rect 339592 237662 339644 237668
rect 338212 237584 338264 237590
rect 338212 237526 338264 237532
rect 338120 237448 338172 237454
rect 338120 237390 338172 237396
rect 337292 204128 337344 204134
rect 337292 204070 337344 204076
rect 337384 204128 337436 204134
rect 337384 204070 337436 204076
rect 337304 203794 337332 204070
rect 337292 203788 337344 203794
rect 337292 203730 337344 203736
rect 337936 203720 337988 203726
rect 337936 203662 337988 203668
rect 336004 203390 336056 203396
rect 336738 203416 336794 203425
rect 335820 203380 335872 203386
rect 336738 203351 336794 203360
rect 335820 203322 335872 203328
rect 333886 203280 333942 203289
rect 333886 203215 333942 203224
rect 335266 203280 335322 203289
rect 335266 203215 335322 203224
rect 336556 203244 336608 203250
rect 336556 203186 336608 203192
rect 336568 203153 336596 203186
rect 328274 203144 328330 203153
rect 328274 203079 328330 203088
rect 332414 203144 332470 203153
rect 332414 203079 332470 203088
rect 333794 203144 333850 203153
rect 336554 203144 336610 203153
rect 333794 203079 333850 203088
rect 335268 203108 335320 203114
rect 336554 203079 336610 203088
rect 335268 203050 335320 203056
rect 335280 203017 335308 203050
rect 337948 203017 337976 203662
rect 338224 203289 338252 237526
rect 339224 203380 339276 203386
rect 339224 203322 339276 203328
rect 338210 203280 338266 203289
rect 338210 203215 338266 203224
rect 339236 203017 339264 203322
rect 339604 203289 339632 237662
rect 340156 237658 340184 240094
rect 341524 238196 341576 238202
rect 341524 238138 341576 238144
rect 340144 237652 340196 237658
rect 340144 237594 340196 237600
rect 340972 204128 341024 204134
rect 340972 204070 341024 204076
rect 340052 203788 340104 203794
rect 340052 203730 340104 203736
rect 340064 203561 340092 203730
rect 340696 203720 340748 203726
rect 340984 203697 341012 204070
rect 340970 203688 341026 203697
rect 340748 203668 340828 203674
rect 340696 203662 340828 203668
rect 340604 203652 340656 203658
rect 340708 203646 340828 203662
rect 340604 203594 340656 203600
rect 340050 203552 340106 203561
rect 340050 203487 340106 203496
rect 339590 203280 339646 203289
rect 339590 203215 339646 203224
rect 340616 203182 340644 203594
rect 340800 203182 340828 203646
rect 341536 203658 341564 238138
rect 342364 237862 342392 240094
rect 344572 238746 344600 240094
rect 344560 238740 344612 238746
rect 344560 238682 344612 238688
rect 346780 238678 346808 240094
rect 346768 238672 346820 238678
rect 346768 238614 346820 238620
rect 349172 238610 349200 240094
rect 349160 238604 349212 238610
rect 349160 238546 349212 238552
rect 351104 238542 351132 240094
rect 351092 238536 351144 238542
rect 351092 238478 351144 238484
rect 353312 238474 353340 240094
rect 353300 238468 353352 238474
rect 353300 238410 353352 238416
rect 342904 238400 342956 238406
rect 342904 238342 342956 238348
rect 342352 237856 342404 237862
rect 342352 237798 342404 237804
rect 342812 204264 342864 204270
rect 342812 204206 342864 204212
rect 342824 204134 342852 204206
rect 342812 204128 342864 204134
rect 342812 204070 342864 204076
rect 341708 203924 341760 203930
rect 341708 203866 341760 203872
rect 340970 203623 341026 203632
rect 341524 203652 341576 203658
rect 341524 203594 341576 203600
rect 341720 203425 341748 203866
rect 342260 203720 342312 203726
rect 342258 203688 342260 203697
rect 342812 203720 342864 203726
rect 342312 203688 342314 203697
rect 342812 203662 342864 203668
rect 342258 203623 342314 203632
rect 342260 203584 342312 203590
rect 342258 203552 342260 203561
rect 342720 203584 342772 203590
rect 342312 203552 342314 203561
rect 342720 203526 342772 203532
rect 342258 203487 342314 203496
rect 341706 203416 341762 203425
rect 342732 203386 342760 203526
rect 341706 203351 341762 203360
rect 342720 203380 342772 203386
rect 342720 203322 342772 203328
rect 341340 203312 341392 203318
rect 341340 203254 341392 203260
rect 340604 203176 340656 203182
rect 340604 203118 340656 203124
rect 340788 203176 340840 203182
rect 340788 203118 340840 203124
rect 341352 203017 341380 203254
rect 342824 203114 342852 203662
rect 342916 203318 342944 238342
rect 344284 238332 344336 238338
rect 344284 238274 344336 238280
rect 342996 238264 343048 238270
rect 342996 238206 343048 238212
rect 342904 203312 342956 203318
rect 342904 203254 342956 203260
rect 342812 203108 342864 203114
rect 342812 203050 342864 203056
rect 342904 203108 342956 203114
rect 342904 203050 342956 203056
rect 335266 203008 335322 203017
rect 335266 202943 335322 202952
rect 336646 203008 336702 203017
rect 336646 202943 336648 202952
rect 336700 202943 336702 202952
rect 337934 203008 337990 203017
rect 337934 202943 337990 202952
rect 339222 203008 339278 203017
rect 339222 202943 339278 202952
rect 341338 203008 341394 203017
rect 342916 202978 342944 203050
rect 343008 202978 343036 238206
rect 343640 203720 343692 203726
rect 343640 203662 343692 203668
rect 343652 203561 343680 203662
rect 343638 203552 343694 203561
rect 343638 203487 343694 203496
rect 343640 203448 343692 203454
rect 343640 203390 343692 203396
rect 344192 203448 344244 203454
rect 344192 203390 344244 203396
rect 343652 203153 343680 203390
rect 344204 203182 344232 203390
rect 344296 203182 344324 238274
rect 347044 238128 347096 238134
rect 347044 238070 347096 238076
rect 345664 238060 345716 238066
rect 345664 238002 345716 238008
rect 345020 203856 345072 203862
rect 345020 203798 345072 203804
rect 345572 203856 345624 203862
rect 345572 203798 345624 203804
rect 344192 203176 344244 203182
rect 343638 203144 343694 203153
rect 344192 203118 344244 203124
rect 344284 203176 344336 203182
rect 345032 203153 345060 203798
rect 345584 203425 345612 203798
rect 345676 203794 345704 238002
rect 347056 204270 347084 238070
rect 347780 204332 347832 204338
rect 347780 204274 347832 204280
rect 347044 204264 347096 204270
rect 347792 204241 347820 204274
rect 351920 204264 351972 204270
rect 347044 204206 347096 204212
rect 347778 204232 347834 204241
rect 351920 204206 351972 204212
rect 347778 204167 347834 204176
rect 347780 204128 347832 204134
rect 347780 204070 347832 204076
rect 345664 203788 345716 203794
rect 345664 203730 345716 203736
rect 347792 203697 347820 204070
rect 349160 203992 349212 203998
rect 349160 203934 349212 203940
rect 349172 203697 349200 203934
rect 349436 203924 349488 203930
rect 349436 203866 349488 203872
rect 347778 203688 347834 203697
rect 347778 203623 347834 203632
rect 349158 203688 349214 203697
rect 349158 203623 349214 203632
rect 348424 203584 348476 203590
rect 348424 203526 348476 203532
rect 346400 203516 346452 203522
rect 346400 203458 346452 203464
rect 345570 203416 345626 203425
rect 345570 203351 345626 203360
rect 346412 203289 346440 203458
rect 347044 203448 347096 203454
rect 347044 203390 347096 203396
rect 346398 203280 346454 203289
rect 345940 203244 345992 203250
rect 346398 203215 346454 203224
rect 345940 203186 345992 203192
rect 344284 203118 344336 203124
rect 345018 203144 345074 203153
rect 343638 203079 343694 203088
rect 344928 203108 344980 203114
rect 345018 203079 345074 203088
rect 344928 203050 344980 203056
rect 344940 203017 344968 203050
rect 345952 203017 345980 203186
rect 347056 203017 347084 203390
rect 348436 203017 348464 203526
rect 349160 203312 349212 203318
rect 349158 203280 349160 203289
rect 349212 203280 349214 203289
rect 349158 203215 349214 203224
rect 349448 203017 349476 203866
rect 351644 203856 351696 203862
rect 351644 203798 351696 203804
rect 351184 203312 351236 203318
rect 351184 203254 351236 203260
rect 351196 203182 351224 203254
rect 351092 203176 351144 203182
rect 351090 203144 351092 203153
rect 351184 203176 351236 203182
rect 351144 203144 351146 203153
rect 351184 203118 351236 203124
rect 351090 203079 351146 203088
rect 351196 203017 351224 203118
rect 351656 203017 351684 203798
rect 351932 203697 351960 204206
rect 354036 204128 354088 204134
rect 354036 204070 354088 204076
rect 354048 203930 354076 204070
rect 355322 203960 355378 203969
rect 354036 203924 354088 203930
rect 355322 203895 355378 203904
rect 354036 203866 354088 203872
rect 354588 203856 354640 203862
rect 354588 203798 354640 203804
rect 353024 203720 353076 203726
rect 351918 203688 351974 203697
rect 353024 203662 353076 203668
rect 351918 203623 351974 203632
rect 353036 203017 353064 203662
rect 354600 203114 354628 203798
rect 354680 203652 354732 203658
rect 354680 203594 354732 203600
rect 354692 203561 354720 203594
rect 354678 203552 354734 203561
rect 354678 203487 354734 203496
rect 355336 203425 355364 203895
rect 355600 203652 355652 203658
rect 355600 203594 355652 203600
rect 355322 203416 355378 203425
rect 355322 203351 355378 203360
rect 355612 203250 355640 203594
rect 355980 203561 356008 240094
rect 357348 204332 357400 204338
rect 357348 204274 357400 204280
rect 357360 204241 357388 204274
rect 357346 204232 357402 204241
rect 357346 204167 357402 204176
rect 357440 204196 357492 204202
rect 357440 204138 357492 204144
rect 357992 204196 358044 204202
rect 357992 204138 358044 204144
rect 356060 204060 356112 204066
rect 356060 204002 356112 204008
rect 355966 203552 356022 203561
rect 355966 203487 356022 203496
rect 356072 203289 356100 204002
rect 357452 203969 357480 204138
rect 357438 203960 357494 203969
rect 357438 203895 357494 203904
rect 358004 203590 358032 204138
rect 358636 204128 358688 204134
rect 358636 204070 358688 204076
rect 357992 203584 358044 203590
rect 357992 203526 358044 203532
rect 356428 203448 356480 203454
rect 356428 203390 356480 203396
rect 356058 203280 356114 203289
rect 355600 203244 355652 203250
rect 356058 203215 356114 203224
rect 355600 203186 355652 203192
rect 354588 203108 354640 203114
rect 354588 203050 354640 203056
rect 354600 203017 354628 203050
rect 355612 203017 355640 203186
rect 356440 203017 356468 203390
rect 358004 203153 358032 203526
rect 357990 203144 358046 203153
rect 357990 203079 358046 203088
rect 357440 203040 357492 203046
rect 344926 203008 344982 203017
rect 341338 202943 341394 202952
rect 342904 202972 342956 202978
rect 336648 202914 336700 202920
rect 342904 202914 342956 202920
rect 342996 202972 343048 202978
rect 344926 202943 344982 202952
rect 345938 203008 345994 203017
rect 345938 202943 345994 202952
rect 347042 203008 347098 203017
rect 347042 202943 347098 202952
rect 348422 203008 348478 203017
rect 348422 202943 348478 202952
rect 349434 203008 349490 203017
rect 349434 202943 349490 202952
rect 351182 203008 351238 203017
rect 351182 202943 351238 202952
rect 351642 203008 351698 203017
rect 351642 202943 351698 202952
rect 353022 203008 353078 203017
rect 353022 202943 353078 202952
rect 353298 203008 353354 203017
rect 353298 202943 353300 202952
rect 342996 202914 343048 202920
rect 353352 202943 353354 202952
rect 354586 203008 354642 203017
rect 354586 202943 354642 202952
rect 355598 203008 355654 203017
rect 355598 202943 355654 202952
rect 356426 203008 356482 203017
rect 356426 202943 356482 202952
rect 357438 203008 357440 203017
rect 358648 203017 358676 204070
rect 358740 203697 358768 240094
rect 360580 238066 360608 240094
rect 360568 238060 360620 238066
rect 360568 238002 360620 238008
rect 362880 204241 362908 240094
rect 364996 237454 365024 240094
rect 366882 239850 366910 240108
rect 366836 239822 366910 239850
rect 368768 240094 369104 240122
rect 364984 237448 365036 237454
rect 364984 237390 365036 237396
rect 366364 237448 366416 237454
rect 366364 237390 366416 237396
rect 362866 204232 362922 204241
rect 362866 204167 362922 204176
rect 364984 204128 365036 204134
rect 364984 204070 365036 204076
rect 360016 204060 360068 204066
rect 360016 204002 360068 204008
rect 358726 203688 358782 203697
rect 358726 203623 358782 203632
rect 360028 203182 360056 204002
rect 361304 203992 361356 203998
rect 361304 203934 361356 203940
rect 360198 203552 360254 203561
rect 360198 203487 360254 203496
rect 360016 203176 360068 203182
rect 360212 203153 360240 203487
rect 360016 203118 360068 203124
rect 360198 203144 360254 203153
rect 360028 203017 360056 203118
rect 360198 203079 360254 203088
rect 361316 203017 361344 203934
rect 362868 203924 362920 203930
rect 362868 203866 362920 203872
rect 362880 203726 362908 203866
rect 363420 203856 363472 203862
rect 363420 203798 363472 203804
rect 362868 203720 362920 203726
rect 362868 203662 362920 203668
rect 362880 203017 362908 203662
rect 363432 203017 363460 203798
rect 364340 203788 364392 203794
rect 364340 203730 364392 203736
rect 364352 203425 364380 203730
rect 364996 203590 365024 204070
rect 365076 203652 365128 203658
rect 365076 203594 365128 203600
rect 364984 203584 365036 203590
rect 364984 203526 365036 203532
rect 364338 203416 364394 203425
rect 364338 203351 364394 203360
rect 365088 203017 365116 203594
rect 366376 203318 366404 237390
rect 366836 203425 366864 239822
rect 367008 237516 367060 237522
rect 367008 237458 367060 237464
rect 366916 237448 366968 237454
rect 366916 237390 366968 237396
rect 366822 203416 366878 203425
rect 366822 203351 366878 203360
rect 366364 203312 366416 203318
rect 366928 203289 366956 237390
rect 366364 203254 366416 203260
rect 366914 203280 366970 203289
rect 366914 203215 366970 203224
rect 367020 203153 367048 237458
rect 368768 237454 368796 240094
rect 371298 239850 371326 240108
rect 371252 239822 371326 239850
rect 371148 238264 371200 238270
rect 371148 238206 371200 238212
rect 368756 237448 368808 237454
rect 368756 237390 368808 237396
rect 367098 204232 367154 204241
rect 367098 204167 367154 204176
rect 367112 204134 367140 204167
rect 367100 204128 367152 204134
rect 367100 204070 367152 204076
rect 369860 203652 369912 203658
rect 369860 203594 369912 203600
rect 369872 203522 369900 203594
rect 369860 203516 369912 203522
rect 369860 203458 369912 203464
rect 368480 203312 368532 203318
rect 368478 203280 368480 203289
rect 371160 203289 371188 238206
rect 371252 237522 371280 239822
rect 371240 237516 371292 237522
rect 371240 237458 371292 237464
rect 368532 203280 368534 203289
rect 368478 203215 368534 203224
rect 371146 203280 371202 203289
rect 371146 203215 371202 203224
rect 373276 203153 373304 240382
rect 373520 240094 373948 240122
rect 375728 240094 376064 240122
rect 377936 240094 378088 240122
rect 380144 240094 380848 240122
rect 382352 240094 382688 240122
rect 384468 240094 384988 240122
rect 386676 240094 387012 240122
rect 388884 240094 389128 240122
rect 373920 204950 373948 240094
rect 376036 237454 376064 240094
rect 376024 237448 376076 237454
rect 376024 237390 376076 237396
rect 376668 237448 376720 237454
rect 376668 237390 376720 237396
rect 373908 204944 373960 204950
rect 373908 204886 373960 204892
rect 374644 204264 374696 204270
rect 374644 204206 374696 204212
rect 374656 203590 374684 204206
rect 376576 204128 376628 204134
rect 376576 204070 376628 204076
rect 376588 203833 376616 204070
rect 376574 203824 376630 203833
rect 376574 203759 376630 203768
rect 376390 203688 376446 203697
rect 376300 203652 376352 203658
rect 376574 203688 376630 203697
rect 376446 203646 376574 203674
rect 376390 203623 376446 203632
rect 376574 203623 376630 203632
rect 376300 203594 376352 203600
rect 374644 203584 374696 203590
rect 374644 203526 374696 203532
rect 376312 203522 376340 203594
rect 376300 203516 376352 203522
rect 376300 203458 376352 203464
rect 375654 203280 375710 203289
rect 375654 203215 375710 203224
rect 367006 203144 367062 203153
rect 367006 203079 367062 203088
rect 373262 203144 373318 203153
rect 373262 203079 373318 203088
rect 375668 203017 375696 203215
rect 357492 203008 357494 203017
rect 357438 202943 357494 202952
rect 358634 203008 358690 203017
rect 358634 202943 358690 202952
rect 358818 203008 358874 203017
rect 358818 202943 358874 202952
rect 360014 203008 360070 203017
rect 360014 202943 360070 202952
rect 361302 203008 361358 203017
rect 361302 202943 361358 202952
rect 362866 203008 362922 203017
rect 362866 202943 362922 202952
rect 363418 203008 363474 203017
rect 363418 202943 363474 202952
rect 365074 203008 365130 203017
rect 365074 202943 365130 202952
rect 375654 203008 375710 203017
rect 375654 202943 375710 202952
rect 353300 202914 353352 202920
rect 358832 202910 358860 202943
rect 358820 202904 358872 202910
rect 358820 202846 358872 202852
rect 297916 202836 297968 202842
rect 297916 202778 297968 202784
rect 297928 201550 297956 202778
rect 297916 201544 297968 201550
rect 297916 201486 297968 201492
rect 297928 180305 297956 201486
rect 376680 201074 376708 237390
rect 378060 201142 378088 240094
rect 380440 238536 380492 238542
rect 380440 238478 380492 238484
rect 380348 238468 380400 238474
rect 380348 238410 380400 238416
rect 380256 238400 380308 238406
rect 380256 238342 380308 238348
rect 380164 238128 380216 238134
rect 380164 238070 380216 238076
rect 379520 204264 379572 204270
rect 379520 204206 379572 204212
rect 379532 204134 379560 204206
rect 379520 204128 379572 204134
rect 379520 204070 379572 204076
rect 378048 201136 378100 201142
rect 378048 201078 378100 201084
rect 376668 201068 376720 201074
rect 376668 201010 376720 201016
rect 379796 183524 379848 183530
rect 379796 183466 379848 183472
rect 379808 182753 379836 183466
rect 379794 182744 379850 182753
rect 379794 182679 379850 182688
rect 297914 180296 297970 180305
rect 297914 180231 297970 180240
rect 297914 171864 297970 171873
rect 297914 171799 297970 171808
rect 297822 111752 297878 111761
rect 297822 111687 297878 111696
rect 297928 109002 297956 171799
rect 379980 124160 380032 124166
rect 379980 124102 380032 124108
rect 379992 123185 380020 124102
rect 379978 123176 380034 123185
rect 379978 123111 380034 123120
rect 380072 118652 380124 118658
rect 380072 118594 380124 118600
rect 380084 118153 380112 118594
rect 380070 118144 380126 118153
rect 380070 118079 380126 118088
rect 379980 115932 380032 115938
rect 379980 115874 380032 115880
rect 379992 114753 380020 115874
rect 380176 115841 380204 238070
rect 380268 118697 380296 238342
rect 380360 120329 380388 238410
rect 380452 122097 380480 238478
rect 380532 238196 380584 238202
rect 380532 238138 380584 238144
rect 380544 180985 380572 238138
rect 380820 201210 380848 240094
rect 382660 237454 382688 240094
rect 382648 237448 382700 237454
rect 382648 237390 382700 237396
rect 383568 237448 383620 237454
rect 383568 237390 383620 237396
rect 383580 201278 383608 237390
rect 384960 201346 384988 240094
rect 386984 237454 387012 240094
rect 389100 238338 389128 240094
rect 390756 240094 391092 240122
rect 392964 240094 393300 240122
rect 395172 240094 395508 240122
rect 397472 240094 397716 240122
rect 399588 240094 399924 240122
rect 401796 240094 402132 240122
rect 404004 240094 404340 240122
rect 406212 240094 406548 240122
rect 408512 240094 408756 240122
rect 410964 240094 411208 240122
rect 389088 238332 389140 238338
rect 389088 238274 389140 238280
rect 390756 238270 390784 240094
rect 390744 238264 390796 238270
rect 390744 238206 390796 238212
rect 392964 237454 392992 240094
rect 395172 238542 395200 240094
rect 395160 238536 395212 238542
rect 395160 238478 395212 238484
rect 397472 238474 397500 240094
rect 397460 238468 397512 238474
rect 397460 238410 397512 238416
rect 399588 238406 399616 240094
rect 399576 238400 399628 238406
rect 399576 238342 399628 238348
rect 395344 238264 395396 238270
rect 395344 238206 395396 238212
rect 386972 237448 387024 237454
rect 386972 237390 387024 237396
rect 387708 237448 387760 237454
rect 387708 237390 387760 237396
rect 391204 237448 391256 237454
rect 391204 237390 391256 237396
rect 392952 237448 393004 237454
rect 392952 237390 393004 237396
rect 393964 237448 394016 237454
rect 393964 237390 394016 237396
rect 387720 201414 387748 237390
rect 389824 204332 389876 204338
rect 389824 204274 389876 204280
rect 389836 204134 389864 204274
rect 389824 204128 389876 204134
rect 389824 204070 389876 204076
rect 387708 201408 387760 201414
rect 387708 201350 387760 201356
rect 384948 201340 385000 201346
rect 384948 201282 385000 201288
rect 383568 201272 383620 201278
rect 383568 201214 383620 201220
rect 380808 201204 380860 201210
rect 380808 201146 380860 201152
rect 380530 180976 380586 180985
rect 380530 180911 380586 180920
rect 391216 124166 391244 237390
rect 391204 124160 391256 124166
rect 391204 124102 391256 124108
rect 380438 122088 380494 122097
rect 380438 122023 380494 122032
rect 380346 120320 380402 120329
rect 380346 120255 380402 120264
rect 380254 118688 380310 118697
rect 393976 118658 394004 237390
rect 394424 204332 394476 204338
rect 394424 204274 394476 204280
rect 394436 204134 394464 204274
rect 394528 204202 394648 204218
rect 394516 204196 394660 204202
rect 394568 204190 394608 204196
rect 394516 204138 394568 204144
rect 394608 204138 394660 204144
rect 394424 204128 394476 204134
rect 394424 204070 394476 204076
rect 380254 118623 380310 118632
rect 393964 118652 394016 118658
rect 393964 118594 394016 118600
rect 395356 115938 395384 238206
rect 401796 237454 401824 240094
rect 404004 238134 404032 240094
rect 406212 238270 406240 240094
rect 406200 238264 406252 238270
rect 406200 238206 406252 238212
rect 403992 238128 404044 238134
rect 403992 238070 404044 238076
rect 401784 237448 401836 237454
rect 401784 237390 401836 237396
rect 402900 204190 403020 204218
rect 402900 204134 402928 204190
rect 402992 204134 403020 204190
rect 402888 204128 402940 204134
rect 402888 204070 402940 204076
rect 402980 204128 403032 204134
rect 402980 204070 403032 204076
rect 408512 201618 408540 240094
rect 411180 238134 411208 240094
rect 412836 240094 413172 240122
rect 412836 238202 412864 240094
rect 415366 239850 415394 240108
rect 417588 240094 417924 240122
rect 419704 240094 420040 240122
rect 421912 240094 422248 240122
rect 424120 240094 424456 240122
rect 415320 239822 415394 239850
rect 415320 238474 415348 239822
rect 417896 238542 417924 240094
rect 417884 238536 417936 238542
rect 417884 238478 417936 238484
rect 415308 238468 415360 238474
rect 415308 238410 415360 238416
rect 420012 238406 420040 240094
rect 422220 238610 422248 240094
rect 424428 238678 424456 240094
rect 426314 239850 426342 240108
rect 428536 240094 428872 240122
rect 430744 240094 431080 240122
rect 426314 239822 426388 239850
rect 426360 238746 426388 239822
rect 426348 238740 426400 238746
rect 426348 238682 426400 238688
rect 424416 238672 424468 238678
rect 424416 238614 424468 238620
rect 422208 238604 422260 238610
rect 422208 238546 422260 238552
rect 420000 238400 420052 238406
rect 420000 238342 420052 238348
rect 428844 238270 428872 240094
rect 428832 238264 428884 238270
rect 428832 238206 428884 238212
rect 431052 238202 431080 240094
rect 432708 240094 432952 240122
rect 434732 240094 435160 240122
rect 436112 240094 437368 240122
rect 438872 240094 439576 240122
rect 441632 240094 441784 240122
rect 443012 240094 443992 240122
rect 445772 240094 446200 240122
rect 447152 240094 448408 240122
rect 450616 240094 451228 240122
rect 452732 240094 453068 240122
rect 454940 240094 455276 240122
rect 457148 240094 457484 240122
rect 459356 240094 459508 240122
rect 461564 240094 461900 240122
rect 463772 240094 464108 240122
rect 465980 240094 466316 240122
rect 468188 240094 468524 240122
rect 470396 240094 470548 240122
rect 412824 238196 412876 238202
rect 412824 238138 412876 238144
rect 431040 238196 431092 238202
rect 431040 238138 431092 238144
rect 411168 238128 411220 238134
rect 411168 238070 411220 238076
rect 432708 232218 432736 240094
rect 431960 232212 432012 232218
rect 431960 232154 432012 232160
rect 432696 232212 432748 232218
rect 432696 232154 432748 232160
rect 431972 231849 432000 232154
rect 431774 231840 431830 231849
rect 431774 231775 431830 231784
rect 431958 231840 432014 231849
rect 431958 231775 432014 231784
rect 431788 222222 431816 231775
rect 431776 222216 431828 222222
rect 431776 222158 431828 222164
rect 432052 222216 432104 222222
rect 432052 222158 432104 222164
rect 432064 215422 432092 222158
rect 432052 215416 432104 215422
rect 432052 215358 432104 215364
rect 432144 215348 432196 215354
rect 432144 215290 432196 215296
rect 416044 204264 416096 204270
rect 416044 204206 416096 204212
rect 427820 204264 427872 204270
rect 427872 204212 427952 204218
rect 427820 204206 427952 204212
rect 412548 204196 412600 204202
rect 412640 204196 412692 204202
rect 412600 204156 412640 204184
rect 412548 204138 412600 204144
rect 412640 204138 412692 204144
rect 416056 204134 416084 204206
rect 427832 204190 427952 204206
rect 427924 204134 427952 204190
rect 416044 204128 416096 204134
rect 416044 204070 416096 204076
rect 427912 204128 427964 204134
rect 427912 204070 427964 204076
rect 432156 203794 432184 215290
rect 434732 203862 434760 240094
rect 436112 203930 436140 240094
rect 438872 203998 438900 240094
rect 441632 204066 441660 240094
rect 443012 204134 443040 240094
rect 445772 204202 445800 240094
rect 445760 204196 445812 204202
rect 445760 204138 445812 204144
rect 443000 204128 443052 204134
rect 443000 204070 443052 204076
rect 441620 204060 441672 204066
rect 441620 204002 441672 204008
rect 438860 203992 438912 203998
rect 437478 203960 437534 203969
rect 436100 203924 436152 203930
rect 438860 203934 438912 203940
rect 437478 203895 437534 203904
rect 436100 203866 436152 203872
rect 434720 203856 434772 203862
rect 434720 203798 434772 203804
rect 432144 203788 432196 203794
rect 432144 203730 432196 203736
rect 408592 203720 408644 203726
rect 408684 203720 408736 203726
rect 408644 203668 408684 203674
rect 437492 203697 437520 203895
rect 442262 203824 442318 203833
rect 442262 203759 442318 203768
rect 408592 203662 408736 203668
rect 437478 203688 437534 203697
rect 408604 203646 408724 203662
rect 437478 203623 437534 203632
rect 442276 203289 442304 203759
rect 447152 203454 447180 240094
rect 450544 238740 450596 238746
rect 450544 238682 450596 238688
rect 449164 238264 449216 238270
rect 449164 238206 449216 238212
rect 449808 238264 449860 238270
rect 449808 238206 449860 238212
rect 447784 238196 447836 238202
rect 447784 238138 447836 238144
rect 448428 238196 448480 238202
rect 448428 238138 448480 238144
rect 447796 204066 447824 238138
rect 448440 204241 448468 238138
rect 448426 204232 448482 204241
rect 448426 204167 448482 204176
rect 449176 204134 449204 238206
rect 449820 204241 449848 238206
rect 449806 204232 449862 204241
rect 450556 204202 450584 238682
rect 451200 205018 451228 240094
rect 452016 238672 452068 238678
rect 452016 238614 452068 238620
rect 451924 238332 451976 238338
rect 451924 238274 451976 238280
rect 451188 205012 451240 205018
rect 451188 204954 451240 204960
rect 449806 204167 449862 204176
rect 450544 204196 450596 204202
rect 450544 204138 450596 204144
rect 450912 204196 450964 204202
rect 450912 204138 450964 204144
rect 449164 204128 449216 204134
rect 449162 204096 449164 204105
rect 450924 204105 450952 204138
rect 449216 204096 449218 204105
rect 447784 204060 447836 204066
rect 447784 204002 447836 204008
rect 448428 204060 448480 204066
rect 449162 204031 449218 204040
rect 450910 204096 450966 204105
rect 450910 204031 450966 204040
rect 448428 204002 448480 204008
rect 447140 203448 447192 203454
rect 447140 203390 447192 203396
rect 442262 203280 442318 203289
rect 442262 203215 442318 203224
rect 408500 201612 408552 201618
rect 408500 201554 408552 201560
rect 409144 201612 409196 201618
rect 409144 201554 409196 201560
rect 409156 183530 409184 201554
rect 417424 201544 417476 201550
rect 417424 201486 417476 201492
rect 409144 183524 409196 183530
rect 409144 183466 409196 183472
rect 417436 180577 417464 201486
rect 448440 201385 448468 204002
rect 451094 203960 451150 203969
rect 451150 203918 451228 203946
rect 451094 203895 451150 203904
rect 451094 203824 451150 203833
rect 451094 203759 451150 203768
rect 451108 203289 451136 203759
rect 451200 203697 451228 203918
rect 451186 203688 451242 203697
rect 451186 203623 451242 203632
rect 451094 203280 451150 203289
rect 451094 203215 451150 203224
rect 451004 203108 451056 203114
rect 451004 203050 451056 203056
rect 451016 203017 451044 203050
rect 451002 203008 451058 203017
rect 451002 202943 451058 202952
rect 451936 201482 451964 238274
rect 452028 204270 452056 238614
rect 452568 238332 452620 238338
rect 452568 238274 452620 238280
rect 452016 204264 452068 204270
rect 452580 204241 452608 238274
rect 453040 237454 453068 240094
rect 453304 238604 453356 238610
rect 453304 238546 453356 238552
rect 453028 237448 453080 237454
rect 453028 237390 453080 237396
rect 453316 204241 453344 238546
rect 454684 238400 454736 238406
rect 454684 238342 454736 238348
rect 455144 238400 455196 238406
rect 455144 238342 455196 238348
rect 453948 237448 454000 237454
rect 453948 237390 454000 237396
rect 452016 204206 452068 204212
rect 452566 204232 452622 204241
rect 452028 204105 452056 204206
rect 452566 204167 452622 204176
rect 453302 204232 453358 204241
rect 453302 204167 453358 204176
rect 452014 204096 452070 204105
rect 452014 204031 452070 204040
rect 453316 203182 453344 204167
rect 453960 203930 453988 237390
rect 454696 204105 454724 238342
rect 455156 204241 455184 238342
rect 455142 204232 455198 204241
rect 455142 204167 455198 204176
rect 454682 204096 454738 204105
rect 454682 204031 454738 204040
rect 453948 203924 454000 203930
rect 453948 203866 454000 203872
rect 453304 203176 453356 203182
rect 453304 203118 453356 203124
rect 453948 203040 454000 203046
rect 453946 203008 453948 203017
rect 454000 203008 454002 203017
rect 453946 202943 454002 202952
rect 454696 202910 454724 204031
rect 455248 203862 455276 240094
rect 456248 238536 456300 238542
rect 456248 238478 456300 238484
rect 456064 238468 456116 238474
rect 456064 238410 456116 238416
rect 456076 204105 456104 238410
rect 456062 204096 456118 204105
rect 456062 204031 456118 204040
rect 455236 203856 455288 203862
rect 455236 203798 455288 203804
rect 456076 203590 456104 204031
rect 456064 203584 456116 203590
rect 456064 203526 456116 203532
rect 456260 203425 456288 238478
rect 456708 238468 456760 238474
rect 456708 238410 456760 238416
rect 456720 204241 456748 238410
rect 457456 237454 457484 240094
rect 459480 238746 459508 240094
rect 459468 238740 459520 238746
rect 459468 238682 459520 238688
rect 459468 238536 459520 238542
rect 459468 238478 459520 238484
rect 457444 237448 457496 237454
rect 457444 237390 457496 237396
rect 458088 237448 458140 237454
rect 458088 237390 458140 237396
rect 456706 204232 456762 204241
rect 456706 204167 456762 204176
rect 457904 204060 457956 204066
rect 457904 204002 457956 204008
rect 457996 204060 458048 204066
rect 457996 204002 458048 204008
rect 456708 203652 456760 203658
rect 456708 203594 456760 203600
rect 456720 203425 456748 203594
rect 456246 203416 456302 203425
rect 456246 203351 456302 203360
rect 456706 203416 456762 203425
rect 456706 203351 456762 203360
rect 457916 203318 457944 204002
rect 458008 203969 458036 204002
rect 457994 203960 458050 203969
rect 457994 203895 458050 203904
rect 458100 203794 458128 237390
rect 459100 204128 459152 204134
rect 459100 204070 459152 204076
rect 458088 203788 458140 203794
rect 458088 203730 458140 203736
rect 457904 203312 457956 203318
rect 457904 203254 457956 203260
rect 457916 203017 457944 203254
rect 459112 203250 459140 204070
rect 459480 203289 459508 238478
rect 461872 237998 461900 240094
rect 463608 238672 463660 238678
rect 463608 238614 463660 238620
rect 462228 238604 462280 238610
rect 462228 238546 462280 238552
rect 461860 237992 461912 237998
rect 461860 237934 461912 237940
rect 461492 204264 461544 204270
rect 461492 204206 461544 204212
rect 460664 204196 460716 204202
rect 460664 204138 460716 204144
rect 460676 203386 460704 204138
rect 460848 203992 460900 203998
rect 460846 203960 460848 203969
rect 460900 203960 460902 203969
rect 460846 203895 460902 203904
rect 461504 203522 461532 204206
rect 461582 203960 461638 203969
rect 461582 203895 461638 203904
rect 461492 203516 461544 203522
rect 461492 203458 461544 203464
rect 460664 203380 460716 203386
rect 460664 203322 460716 203328
rect 459466 203280 459522 203289
rect 459100 203244 459152 203250
rect 459466 203215 459522 203224
rect 459100 203186 459152 203192
rect 459112 203017 459140 203186
rect 460676 203017 460704 203322
rect 461504 203017 461532 203458
rect 461596 203425 461624 203895
rect 461582 203416 461638 203425
rect 461582 203351 461638 203360
rect 462240 203289 462268 238546
rect 463516 203720 463568 203726
rect 463516 203662 463568 203668
rect 463056 203448 463108 203454
rect 463056 203390 463108 203396
rect 462226 203280 462282 203289
rect 462226 203215 462282 203224
rect 462412 203176 462464 203182
rect 462412 203118 462464 203124
rect 462424 203017 462452 203118
rect 463068 203017 463096 203390
rect 463528 203289 463556 203662
rect 463620 203425 463648 238614
rect 464080 237930 464108 240094
rect 464068 237924 464120 237930
rect 464068 237866 464120 237872
rect 466288 237794 466316 240094
rect 466276 237788 466328 237794
rect 466276 237730 466328 237736
rect 468496 237658 468524 240094
rect 470520 237862 470548 240094
rect 472590 239850 472618 240108
rect 474798 239850 474826 240108
rect 472590 239822 472664 239850
rect 470508 237856 470560 237862
rect 470508 237798 470560 237804
rect 468484 237652 468536 237658
rect 468484 237594 468536 237600
rect 471888 237448 471940 237454
rect 471888 237390 471940 237396
rect 470508 205284 470560 205290
rect 470508 205226 470560 205232
rect 470416 205148 470468 205154
rect 470416 205090 470468 205096
rect 469128 205080 469180 205086
rect 469128 205022 469180 205028
rect 464988 204264 465040 204270
rect 469140 204241 469168 205022
rect 464988 204206 465040 204212
rect 469126 204232 469182 204241
rect 465000 204105 465028 204206
rect 466276 204196 466328 204202
rect 469126 204167 469182 204176
rect 466276 204138 466328 204144
rect 466288 204105 466316 204138
rect 467288 204128 467340 204134
rect 464986 204096 465042 204105
rect 464986 204031 465042 204040
rect 466274 204096 466330 204105
rect 470428 204105 470456 205090
rect 470520 204241 470548 205226
rect 470506 204232 470562 204241
rect 470506 204167 470562 204176
rect 467288 204070 467340 204076
rect 470414 204096 470470 204105
rect 466274 204031 466330 204040
rect 466366 203960 466422 203969
rect 466366 203895 466422 203904
rect 464712 203652 464764 203658
rect 464712 203594 464764 203600
rect 464724 203425 464752 203594
rect 465908 203584 465960 203590
rect 466380 203561 466408 203895
rect 467300 203590 467328 204070
rect 470414 204031 470470 204040
rect 471242 203960 471298 203969
rect 471242 203895 471298 203904
rect 471060 203856 471112 203862
rect 471112 203804 471192 203810
rect 471060 203798 471192 203804
rect 470784 203788 470836 203794
rect 471072 203782 471192 203798
rect 470784 203730 470836 203736
rect 470508 203720 470560 203726
rect 470560 203668 470732 203674
rect 470508 203662 470732 203668
rect 470520 203646 470732 203662
rect 470796 203658 470824 203730
rect 470704 203590 470732 203646
rect 470784 203652 470836 203658
rect 470784 203594 470836 203600
rect 467288 203584 467340 203590
rect 465908 203526 465960 203532
rect 466366 203552 466422 203561
rect 463606 203416 463662 203425
rect 463606 203351 463662 203360
rect 464710 203416 464766 203425
rect 464710 203351 464766 203360
rect 463514 203280 463570 203289
rect 463514 203215 463570 203224
rect 465920 203017 465948 203526
rect 467288 203526 467340 203532
rect 470416 203584 470468 203590
rect 470692 203584 470744 203590
rect 470468 203532 470640 203538
rect 470416 203526 470640 203532
rect 470692 203526 470744 203532
rect 470428 203510 470640 203526
rect 466366 203487 466422 203496
rect 467562 203416 467618 203425
rect 467562 203351 467564 203360
rect 467616 203351 467618 203360
rect 469494 203416 469550 203425
rect 469494 203351 469550 203360
rect 467564 203322 467616 203328
rect 467196 203312 467248 203318
rect 467748 203312 467800 203318
rect 467196 203254 467248 203260
rect 467746 203280 467748 203289
rect 467800 203280 467802 203289
rect 467208 203017 467236 203254
rect 467746 203215 467802 203224
rect 468484 203244 468536 203250
rect 468484 203186 468536 203192
rect 468496 203017 468524 203186
rect 455326 203008 455382 203017
rect 455326 202943 455328 202952
rect 455380 202943 455382 202952
rect 457902 203008 457958 203017
rect 457902 202943 457958 202952
rect 459098 203008 459154 203017
rect 459098 202943 459154 202952
rect 460662 203008 460718 203017
rect 460662 202943 460718 202952
rect 461490 203008 461546 203017
rect 461490 202943 461546 202952
rect 462410 203008 462466 203017
rect 462410 202943 462466 202952
rect 463054 203008 463110 203017
rect 463054 202943 463110 202952
rect 465906 203008 465962 203017
rect 465906 202943 465962 202952
rect 467194 203008 467250 203017
rect 467194 202943 467250 202952
rect 468482 203008 468538 203017
rect 468482 202943 468538 202952
rect 455328 202914 455380 202920
rect 463068 202910 463096 202943
rect 469508 202910 469536 203351
rect 470612 203289 470640 203510
rect 470598 203280 470654 203289
rect 470598 203215 470654 203224
rect 471164 203182 471192 203782
rect 471256 203561 471284 203895
rect 471336 203788 471388 203794
rect 471336 203730 471388 203736
rect 471242 203552 471298 203561
rect 471242 203487 471298 203496
rect 471348 203289 471376 203730
rect 471796 203448 471848 203454
rect 471796 203390 471848 203396
rect 471334 203280 471390 203289
rect 471334 203215 471390 203224
rect 471060 203176 471112 203182
rect 471060 203118 471112 203124
rect 471152 203176 471204 203182
rect 471152 203118 471204 203124
rect 471072 203017 471100 203118
rect 471808 203017 471836 203390
rect 471900 203289 471928 237390
rect 472636 203289 472664 239822
rect 474752 239822 474826 239850
rect 476132 240094 477020 240122
rect 478892 240094 479228 240122
rect 480272 240094 481436 240122
rect 483308 240094 483644 240122
rect 474004 238740 474056 238746
rect 474004 238682 474056 238688
rect 473360 237856 473412 237862
rect 473360 237798 473412 237804
rect 472900 203516 472952 203522
rect 472900 203458 472952 203464
rect 472912 203289 472940 203458
rect 473372 203289 473400 237798
rect 474016 203726 474044 238682
rect 474096 237992 474148 237998
rect 474096 237934 474148 237940
rect 474108 203862 474136 237934
rect 474280 237856 474332 237862
rect 474280 237798 474332 237804
rect 474188 237720 474240 237726
rect 474188 237662 474240 237668
rect 474096 203856 474148 203862
rect 474096 203798 474148 203804
rect 473912 203720 473964 203726
rect 473912 203662 473964 203668
rect 474004 203720 474056 203726
rect 474004 203662 474056 203668
rect 473924 203561 473952 203662
rect 473910 203552 473966 203561
rect 473910 203487 473966 203496
rect 474200 203318 474228 237662
rect 474292 204202 474320 237798
rect 474752 237454 474780 239822
rect 475568 238740 475620 238746
rect 475568 238682 475620 238688
rect 475476 237992 475528 237998
rect 475476 237934 475528 237940
rect 475384 237924 475436 237930
rect 475384 237866 475436 237872
rect 474832 237652 474884 237658
rect 474832 237594 474884 237600
rect 474740 237448 474792 237454
rect 474740 237390 474792 237396
rect 474280 204196 474332 204202
rect 474280 204138 474332 204144
rect 474372 203788 474424 203794
rect 474372 203730 474424 203736
rect 474464 203788 474516 203794
rect 474464 203730 474516 203736
rect 474384 203386 474412 203730
rect 474476 203561 474504 203730
rect 474462 203552 474518 203561
rect 474462 203487 474518 203496
rect 474372 203380 474424 203386
rect 474372 203322 474424 203328
rect 474188 203312 474240 203318
rect 471886 203280 471942 203289
rect 471886 203215 471942 203224
rect 472622 203280 472678 203289
rect 472622 203215 472678 203224
rect 472898 203280 472954 203289
rect 472898 203215 472954 203224
rect 473358 203280 473414 203289
rect 474844 203289 474872 237594
rect 475396 204202 475424 237866
rect 475488 204270 475516 237934
rect 475476 204264 475528 204270
rect 475476 204206 475528 204212
rect 475384 204196 475436 204202
rect 475384 204138 475436 204144
rect 475580 203590 475608 238682
rect 475660 237788 475712 237794
rect 475660 237730 475712 237736
rect 475672 204105 475700 237730
rect 476132 205290 476160 240094
rect 476764 238060 476816 238066
rect 476764 238002 476816 238008
rect 476120 205284 476172 205290
rect 476120 205226 476172 205232
rect 476776 204270 476804 238002
rect 478892 205154 478920 240094
rect 478880 205148 478932 205154
rect 478880 205090 478932 205096
rect 480272 205086 480300 240094
rect 483308 237726 483336 240094
rect 485838 239850 485866 240108
rect 485792 239822 485866 239850
rect 487632 240094 487968 240122
rect 489932 240094 490176 240122
rect 492048 240094 492384 240122
rect 494256 240094 494592 240122
rect 495452 240094 496800 240122
rect 498672 240094 499008 240122
rect 500972 240094 501216 240122
rect 503088 240094 503424 240122
rect 505112 240094 505632 240122
rect 507504 240094 507840 240122
rect 509252 240094 510048 240122
rect 512104 240094 512256 240122
rect 513392 240094 514464 240122
rect 516336 240094 516672 240122
rect 518544 240094 518880 240122
rect 485792 237862 485820 239822
rect 487632 237998 487660 240094
rect 489932 238746 489960 240094
rect 489920 238740 489972 238746
rect 489920 238682 489972 238688
rect 492048 238678 492076 240094
rect 492036 238672 492088 238678
rect 492036 238614 492088 238620
rect 494256 238610 494284 240094
rect 494244 238604 494296 238610
rect 494244 238546 494296 238552
rect 487620 237992 487672 237998
rect 487620 237934 487672 237940
rect 485780 237856 485832 237862
rect 485780 237798 485832 237804
rect 483296 237720 483348 237726
rect 483296 237662 483348 237668
rect 480260 205080 480312 205086
rect 480260 205022 480312 205028
rect 484400 205012 484452 205018
rect 484400 204954 484452 204960
rect 476764 204264 476816 204270
rect 484412 204241 484440 204954
rect 490196 204944 490248 204950
rect 490196 204886 490248 204892
rect 485780 204264 485832 204270
rect 476764 204206 476816 204212
rect 484398 204232 484454 204241
rect 477500 204196 477552 204202
rect 485780 204206 485832 204212
rect 484398 204167 484454 204176
rect 477500 204138 477552 204144
rect 475752 204128 475804 204134
rect 475658 204096 475714 204105
rect 475752 204070 475804 204076
rect 475844 204128 475896 204134
rect 477512 204105 477540 204138
rect 483020 204128 483072 204134
rect 475844 204070 475896 204076
rect 477498 204096 477554 204105
rect 475658 204031 475714 204040
rect 475764 203590 475792 204070
rect 475856 203794 475884 204070
rect 477498 204031 477554 204040
rect 483018 204096 483020 204105
rect 485792 204105 485820 204206
rect 483072 204096 483074 204105
rect 483018 204031 483074 204040
rect 485778 204096 485834 204105
rect 485778 204031 485834 204040
rect 490208 203969 490236 204886
rect 495452 203998 495480 240094
rect 498672 238542 498700 240094
rect 498660 238536 498712 238542
rect 498660 238478 498712 238484
rect 496360 238128 496412 238134
rect 496360 238070 496412 238076
rect 495440 203992 495492 203998
rect 480166 203960 480222 203969
rect 490194 203960 490250 203969
rect 480166 203895 480222 203904
rect 483020 203924 483072 203930
rect 477500 203856 477552 203862
rect 477500 203798 477552 203804
rect 475844 203788 475896 203794
rect 475844 203730 475896 203736
rect 475568 203584 475620 203590
rect 475568 203526 475620 203532
rect 475752 203584 475804 203590
rect 475752 203526 475804 203532
rect 474188 203254 474240 203260
rect 474830 203280 474886 203289
rect 473358 203215 473414 203224
rect 474830 203215 474886 203224
rect 475764 203017 475792 203526
rect 477512 203425 477540 203798
rect 478880 203720 478932 203726
rect 478880 203662 478932 203668
rect 478892 203425 478920 203662
rect 480180 203561 480208 203895
rect 495440 203934 495492 203940
rect 490194 203895 490250 203904
rect 483020 203866 483072 203872
rect 480628 203652 480680 203658
rect 480628 203594 480680 203600
rect 480640 203561 480668 203594
rect 480166 203552 480222 203561
rect 480166 203487 480222 203496
rect 480626 203552 480682 203561
rect 480626 203487 480682 203496
rect 481640 203448 481692 203454
rect 477498 203416 477554 203425
rect 477498 203351 477554 203360
rect 478878 203416 478934 203425
rect 481640 203390 481692 203396
rect 478878 203351 478934 203360
rect 478972 203380 479024 203386
rect 478972 203322 479024 203328
rect 480536 203380 480588 203386
rect 480536 203322 480588 203328
rect 476120 203312 476172 203318
rect 478984 203289 479012 203322
rect 476120 203254 476172 203260
rect 477498 203280 477554 203289
rect 476132 203017 476160 203254
rect 477498 203215 477500 203224
rect 477552 203215 477554 203224
rect 478970 203280 479026 203289
rect 478970 203215 479026 203224
rect 477500 203186 477552 203192
rect 480548 203017 480576 203322
rect 481652 203289 481680 203390
rect 481638 203280 481694 203289
rect 481638 203215 481694 203224
rect 481640 203176 481692 203182
rect 481640 203118 481692 203124
rect 481652 203017 481680 203118
rect 483032 203017 483060 203866
rect 484400 203584 484452 203590
rect 484398 203552 484400 203561
rect 484452 203552 484454 203561
rect 484398 203487 484454 203496
rect 471058 203008 471114 203017
rect 471058 202943 471114 202952
rect 471794 203008 471850 203017
rect 471794 202943 471850 202952
rect 475750 203008 475806 203017
rect 475750 202943 475806 202952
rect 476118 203008 476174 203017
rect 476118 202943 476174 202952
rect 477498 203008 477554 203017
rect 477498 202943 477554 202952
rect 480534 203008 480590 203017
rect 480534 202943 480590 202952
rect 481638 203008 481694 203017
rect 481638 202943 481694 202952
rect 483018 203008 483074 203017
rect 483018 202943 483074 202952
rect 477512 202910 477540 202943
rect 454684 202904 454736 202910
rect 454684 202846 454736 202852
rect 463056 202904 463108 202910
rect 463056 202846 463108 202852
rect 469496 202904 469548 202910
rect 469496 202846 469548 202852
rect 477500 202904 477552 202910
rect 477500 202846 477552 202852
rect 451924 201476 451976 201482
rect 451924 201418 451976 201424
rect 448426 201376 448482 201385
rect 448426 201311 448482 201320
rect 496372 181370 496400 238070
rect 500972 204066 501000 240094
rect 503088 238474 503116 240094
rect 503076 238468 503128 238474
rect 503076 238410 503128 238416
rect 500960 204060 501012 204066
rect 500960 204002 501012 204008
rect 505112 202978 505140 240094
rect 507504 238406 507532 240094
rect 507492 238400 507544 238406
rect 507492 238342 507544 238348
rect 509252 203046 509280 240094
rect 512104 238338 512132 240094
rect 512092 238332 512144 238338
rect 512092 238274 512144 238280
rect 513392 203114 513420 240094
rect 516336 238270 516364 240094
rect 516324 238264 516376 238270
rect 516324 238206 516376 238212
rect 518544 238202 518572 240094
rect 518532 238196 518584 238202
rect 518532 238138 518584 238144
rect 513380 203108 513432 203114
rect 513380 203050 513432 203056
rect 509240 203040 509292 203046
rect 509240 202982 509292 202988
rect 505100 202972 505152 202978
rect 505100 202914 505152 202920
rect 500316 201612 500368 201618
rect 500316 201554 500368 201560
rect 499672 201476 499724 201482
rect 499672 201418 499724 201424
rect 496450 181384 496506 181393
rect 496372 181342 496450 181370
rect 496450 181319 496506 181328
rect 417422 180568 417478 180577
rect 417422 180503 417478 180512
rect 418066 171728 418122 171737
rect 418066 171663 418122 171672
rect 395344 115932 395396 115938
rect 395344 115874 395396 115880
rect 380162 115832 380218 115841
rect 380162 115767 380218 115776
rect 379978 114744 380034 114753
rect 379978 114679 380034 114688
rect 300766 111344 300822 111353
rect 300766 111279 300822 111288
rect 416778 111344 416834 111353
rect 416778 111279 416834 111288
rect 300780 110974 300808 111279
rect 416792 110974 416820 111279
rect 300768 110968 300820 110974
rect 300768 110910 300820 110916
rect 416780 110968 416832 110974
rect 416780 110910 416832 110916
rect 303618 109032 303674 109041
rect 297916 108996 297968 109002
rect 307758 109032 307814 109041
rect 303618 108967 303620 108976
rect 297916 108938 297968 108944
rect 303672 108967 303674 108976
rect 305644 108996 305696 109002
rect 303620 108938 303672 108944
rect 418080 109002 418108 171663
rect 499684 115297 499712 201418
rect 500224 201408 500276 201414
rect 500224 201350 500276 201356
rect 499856 201340 499908 201346
rect 499856 201282 499908 201288
rect 499764 201272 499816 201278
rect 499764 201214 499816 201220
rect 499776 118697 499804 201214
rect 499762 118688 499818 118697
rect 499762 118623 499818 118632
rect 499868 118153 499896 201282
rect 499948 201204 500000 201210
rect 499948 201146 500000 201152
rect 499960 120873 499988 201146
rect 500040 201136 500092 201142
rect 500040 201078 500092 201084
rect 500052 122097 500080 201078
rect 500132 201068 500184 201074
rect 500132 201010 500184 201016
rect 500144 123729 500172 201010
rect 500130 123720 500186 123729
rect 500130 123655 500186 123664
rect 500038 122088 500094 122097
rect 500038 122023 500094 122032
rect 499946 120864 500002 120873
rect 499946 120799 500002 120808
rect 499854 118144 499910 118153
rect 499854 118079 499910 118088
rect 500236 115841 500264 201350
rect 500328 183161 500356 201554
rect 521672 200870 521700 459983
rect 521750 455832 521806 455841
rect 521750 455767 521806 455776
rect 521764 200938 521792 455767
rect 521842 453656 521898 453665
rect 521842 453591 521898 453600
rect 521856 201006 521884 453591
rect 521934 451616 521990 451625
rect 521934 451551 521990 451560
rect 521844 201000 521896 201006
rect 521844 200942 521896 200948
rect 521752 200932 521804 200938
rect 521752 200874 521804 200880
rect 521660 200864 521712 200870
rect 521660 200806 521712 200812
rect 521948 200802 521976 451551
rect 522026 449440 522082 449449
rect 522026 449375 522082 449384
rect 522040 208350 522068 449375
rect 522118 447400 522174 447409
rect 522118 447335 522174 447344
rect 522132 237386 522160 447335
rect 522210 443184 522266 443193
rect 522210 443119 522266 443128
rect 522224 437646 522252 443119
rect 522212 437640 522264 437646
rect 522212 437582 522264 437588
rect 522212 437504 522264 437510
rect 522212 437446 522264 437452
rect 522120 237380 522172 237386
rect 522120 237322 522172 237328
rect 522118 237144 522174 237153
rect 522118 237079 522174 237088
rect 522028 208344 522080 208350
rect 522028 208286 522080 208292
rect 521936 200796 521988 200802
rect 521936 200738 521988 200744
rect 500314 183152 500370 183161
rect 500314 183087 500370 183096
rect 500222 115832 500278 115841
rect 500222 115767 500278 115776
rect 499670 115288 499726 115297
rect 499670 115223 499726 115232
rect 424230 109032 424286 109041
rect 307758 108967 307760 108976
rect 305644 108938 305696 108944
rect 307812 108967 307814 108976
rect 418068 108996 418120 109002
rect 307760 108938 307812 108944
rect 424230 108967 424232 108976
rect 418068 108938 418120 108944
rect 424284 108967 424286 108976
rect 427818 109032 427874 109041
rect 427818 108967 427820 108976
rect 424232 108938 424284 108944
rect 427872 108967 427874 108976
rect 427820 108938 427872 108944
rect 278136 3528 278188 3534
rect 278136 3470 278188 3476
rect 278044 3460 278096 3466
rect 278044 3402 278096 3408
rect 305656 2854 305684 108938
rect 522132 8294 522160 237079
rect 522224 223582 522252 437446
rect 522316 401033 522344 478178
rect 522396 478032 522448 478038
rect 522396 477974 522448 477980
rect 522408 441017 522436 477974
rect 522394 441008 522450 441017
rect 522394 440943 522450 440952
rect 522394 438968 522450 438977
rect 522394 438903 522450 438912
rect 522302 401024 522358 401033
rect 522302 400959 522358 400968
rect 522304 324148 522356 324154
rect 522304 324090 522356 324096
rect 522316 323105 522344 324090
rect 522302 323096 522358 323105
rect 522302 323031 522358 323040
rect 522304 316940 522356 316946
rect 522304 316882 522356 316888
rect 522316 316849 522344 316882
rect 522302 316840 522358 316849
rect 522302 316775 522358 316784
rect 522304 310480 522356 310486
rect 522302 310448 522304 310457
rect 522356 310448 522358 310457
rect 522302 310383 522358 310392
rect 522304 304836 522356 304842
rect 522304 304778 522356 304784
rect 522316 304201 522344 304778
rect 522302 304192 522358 304201
rect 522302 304127 522358 304136
rect 522304 294636 522356 294642
rect 522304 294578 522356 294584
rect 522316 278905 522344 294578
rect 522302 278896 522358 278905
rect 522302 278831 522358 278840
rect 522302 272640 522358 272649
rect 522302 272575 522358 272584
rect 522316 252550 522344 272575
rect 522304 252544 522356 252550
rect 522304 252486 522356 252492
rect 522302 249384 522358 249393
rect 522302 249319 522358 249328
rect 522316 248470 522344 249319
rect 522304 248464 522356 248470
rect 522304 248406 522356 248412
rect 522302 247344 522358 247353
rect 522302 247279 522358 247288
rect 522316 247110 522344 247279
rect 522304 247104 522356 247110
rect 522304 247046 522356 247052
rect 522302 245168 522358 245177
rect 522302 245103 522358 245112
rect 522212 223576 522264 223582
rect 522212 223518 522264 223524
rect 522316 30326 522344 245103
rect 522408 243234 522436 438903
rect 522500 407425 522528 478246
rect 522580 478168 522632 478174
rect 522580 478110 522632 478116
rect 522592 409465 522620 478110
rect 522684 430545 522712 478382
rect 522856 478372 522908 478378
rect 522856 478314 522908 478320
rect 522764 478100 522816 478106
rect 522764 478042 522816 478048
rect 522670 430536 522726 430545
rect 522670 430471 522726 430480
rect 522776 422113 522804 478042
rect 522868 436801 522896 478314
rect 522946 445224 523002 445233
rect 522946 445159 523002 445168
rect 522960 437510 522988 445159
rect 522948 437504 523000 437510
rect 522948 437446 523000 437452
rect 522854 436792 522910 436801
rect 522854 436727 522910 436736
rect 522946 426320 523002 426329
rect 523052 426306 523080 478926
rect 523144 428369 523172 478994
rect 523130 428360 523186 428369
rect 523130 428295 523186 428304
rect 523002 426278 523080 426306
rect 522946 426255 523002 426264
rect 522762 422104 522818 422113
rect 522762 422039 522818 422048
rect 522672 420096 522724 420102
rect 522670 420064 522672 420073
rect 522724 420064 522726 420073
rect 522670 419999 522726 420008
rect 522578 409456 522634 409465
rect 522578 409391 522634 409400
rect 522486 407416 522542 407425
rect 522486 407351 522542 407360
rect 522948 340876 523000 340882
rect 522948 340818 523000 340824
rect 522960 339969 522988 340818
rect 522946 339960 523002 339969
rect 522946 339895 523002 339904
rect 522948 337952 523000 337958
rect 522946 337920 522948 337929
rect 523000 337920 523002 337929
rect 522946 337855 523002 337864
rect 522580 336728 522632 336734
rect 522580 336670 522632 336676
rect 522592 335753 522620 336670
rect 522578 335744 522634 335753
rect 522578 335679 522634 335688
rect 522948 333940 523000 333946
rect 522948 333882 523000 333888
rect 522960 333713 522988 333882
rect 522946 333704 523002 333713
rect 522946 333639 523002 333648
rect 522580 332580 522632 332586
rect 522580 332522 522632 332528
rect 522592 331537 522620 332522
rect 522578 331528 522634 331537
rect 522578 331463 522634 331472
rect 522946 329488 523002 329497
rect 522946 329423 523002 329432
rect 522960 328574 522988 329423
rect 522948 328568 523000 328574
rect 522948 328510 523000 328516
rect 522948 328432 523000 328438
rect 522948 328374 523000 328380
rect 522960 327321 522988 328374
rect 522946 327312 523002 327321
rect 522946 327247 523002 327256
rect 522948 325644 523000 325650
rect 522948 325586 523000 325592
rect 522960 325281 522988 325586
rect 522946 325272 523002 325281
rect 522946 325207 523002 325216
rect 522672 321564 522724 321570
rect 522672 321506 522724 321512
rect 522684 321065 522712 321506
rect 522670 321056 522726 321065
rect 522670 320991 522726 321000
rect 522948 320136 523000 320142
rect 522948 320078 523000 320084
rect 522960 318889 522988 320078
rect 522946 318880 523002 318889
rect 522946 318815 523002 318824
rect 523696 316946 523724 579634
rect 523776 532772 523828 532778
rect 523776 532714 523828 532720
rect 523684 316940 523736 316946
rect 523684 316882 523736 316888
rect 522946 314664 523002 314673
rect 522946 314599 522948 314608
rect 523000 314599 523002 314608
rect 522948 314570 523000 314576
rect 522948 313268 523000 313274
rect 522948 313210 523000 313216
rect 522960 312633 522988 313210
rect 522946 312624 523002 312633
rect 522946 312559 523002 312568
rect 523788 310486 523816 532714
rect 523868 485852 523920 485858
rect 523868 485794 523920 485800
rect 523776 310480 523828 310486
rect 523776 310422 523828 310428
rect 522948 309120 523000 309126
rect 522948 309062 523000 309068
rect 522960 308417 522988 309062
rect 522946 308408 523002 308417
rect 522946 308343 523002 308352
rect 522948 306332 523000 306338
rect 522948 306274 523000 306280
rect 522960 306241 522988 306274
rect 522946 306232 523002 306241
rect 522946 306167 523002 306176
rect 523880 304842 523908 485794
rect 524420 477964 524472 477970
rect 524420 477906 524472 477912
rect 524432 420102 524460 477906
rect 524420 420096 524472 420102
rect 524420 420038 524472 420044
rect 523960 392012 524012 392018
rect 523960 391954 524012 391960
rect 523868 304836 523920 304842
rect 523868 304778 523920 304784
rect 522948 302184 523000 302190
rect 522948 302126 523000 302132
rect 522960 302025 522988 302126
rect 522946 302016 523002 302025
rect 522946 301951 523002 301960
rect 522948 300824 523000 300830
rect 522948 300766 523000 300772
rect 522960 299985 522988 300766
rect 522946 299976 523002 299985
rect 522946 299911 523002 299920
rect 522948 298104 523000 298110
rect 522948 298046 523000 298052
rect 522960 297945 522988 298046
rect 522946 297936 523002 297945
rect 522946 297871 523002 297880
rect 522948 296676 523000 296682
rect 522948 296618 523000 296624
rect 522960 295769 522988 296618
rect 522946 295760 523002 295769
rect 522946 295695 523002 295704
rect 522488 294704 522540 294710
rect 522488 294646 522540 294652
rect 522500 283121 522528 294646
rect 522948 293956 523000 293962
rect 522948 293898 523000 293904
rect 522960 293729 522988 293898
rect 522946 293720 523002 293729
rect 522946 293655 523002 293664
rect 523972 292058 524000 391954
rect 525076 324154 525104 626554
rect 527192 337958 527220 703520
rect 543476 703474 543504 703520
rect 543476 703446 543596 703474
rect 531964 700324 532016 700330
rect 531964 700266 532016 700272
rect 529204 673532 529256 673538
rect 529204 673474 529256 673480
rect 527180 337952 527232 337958
rect 527180 337894 527232 337900
rect 529216 328574 529244 673474
rect 531976 336734 532004 700266
rect 543568 698290 543596 703446
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 542728 698284 542780 698290
rect 542728 698226 542780 698232
rect 543556 698284 543608 698290
rect 543556 698226 543608 698232
rect 542740 694142 542768 698226
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 545764 696992 545816 696998
rect 545764 696934 545816 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 542544 694136 542596 694142
rect 542544 694078 542596 694084
rect 542728 694136 542780 694142
rect 542728 694078 542780 694084
rect 542556 684554 542584 694078
rect 542452 684548 542504 684554
rect 542452 684490 542504 684496
rect 542544 684548 542596 684554
rect 542544 684490 542596 684496
rect 542464 684457 542492 684490
rect 542450 684448 542506 684457
rect 542450 684383 542506 684392
rect 542542 678872 542598 678881
rect 542542 678807 542598 678816
rect 542556 666602 542584 678807
rect 542544 666596 542596 666602
rect 542544 666538 542596 666544
rect 542820 666596 542872 666602
rect 542820 666538 542872 666544
rect 542832 661774 542860 666538
rect 542544 661768 542596 661774
rect 542544 661710 542596 661716
rect 542820 661768 542872 661774
rect 542820 661710 542872 661716
rect 542556 656946 542584 661710
rect 542544 656940 542596 656946
rect 542544 656882 542596 656888
rect 542636 656940 542688 656946
rect 542636 656882 542688 656888
rect 540244 650072 540296 650078
rect 540244 650014 540296 650020
rect 538864 603152 538916 603158
rect 538864 603094 538916 603100
rect 537484 556232 537536 556238
rect 537484 556174 537536 556180
rect 536104 509312 536156 509318
rect 536104 509254 536156 509260
rect 534724 438932 534776 438938
rect 534724 438874 534776 438880
rect 531964 336728 532016 336734
rect 531964 336670 532016 336676
rect 529204 328568 529256 328574
rect 529204 328510 529256 328516
rect 525064 324148 525116 324154
rect 525064 324090 525116 324096
rect 534736 298110 534764 438874
rect 536116 306338 536144 509254
rect 537496 313274 537524 556174
rect 538876 320142 538904 603094
rect 540256 325650 540284 650014
rect 542648 647290 542676 656882
rect 542544 647284 542596 647290
rect 542544 647226 542596 647232
rect 542636 647284 542688 647290
rect 542636 647226 542688 647232
rect 542556 640422 542584 647226
rect 542544 640416 542596 640422
rect 542544 640358 542596 640364
rect 542636 640416 542688 640422
rect 542636 640358 542688 640364
rect 542648 630698 542676 640358
rect 542452 630692 542504 630698
rect 542452 630634 542504 630640
rect 542636 630692 542688 630698
rect 542636 630634 542688 630640
rect 542464 630578 542492 630634
rect 542464 630550 542584 630578
rect 542556 621058 542584 630550
rect 542556 621030 542676 621058
rect 542648 611386 542676 621030
rect 542452 611380 542504 611386
rect 542452 611322 542504 611328
rect 542636 611380 542688 611386
rect 542636 611322 542688 611328
rect 542464 611266 542492 611322
rect 542464 611238 542584 611266
rect 542556 608598 542584 611238
rect 542452 608592 542504 608598
rect 542452 608534 542504 608540
rect 542544 608592 542596 608598
rect 542544 608534 542596 608540
rect 542464 601730 542492 608534
rect 542452 601724 542504 601730
rect 542452 601666 542504 601672
rect 542728 601724 542780 601730
rect 542728 601666 542780 601672
rect 542740 598942 542768 601666
rect 542544 598936 542596 598942
rect 542544 598878 542596 598884
rect 542728 598936 542780 598942
rect 542728 598878 542780 598884
rect 542556 589354 542584 598878
rect 542544 589348 542596 589354
rect 542544 589290 542596 589296
rect 542820 589348 542872 589354
rect 542820 589290 542872 589296
rect 542832 582486 542860 589290
rect 542820 582480 542872 582486
rect 542820 582422 542872 582428
rect 542728 582344 542780 582350
rect 542728 582286 542780 582292
rect 542740 572642 542768 582286
rect 542556 572614 542768 572642
rect 542556 569922 542584 572614
rect 542464 569894 542584 569922
rect 542464 563174 542492 569894
rect 542452 563168 542504 563174
rect 542452 563110 542504 563116
rect 542452 563032 542504 563038
rect 542452 562974 542504 562980
rect 542464 560266 542492 562974
rect 542372 560238 542492 560266
rect 542372 553450 542400 560238
rect 542360 553444 542412 553450
rect 542360 553386 542412 553392
rect 542452 553376 542504 553382
rect 542452 553318 542504 553324
rect 542464 550662 542492 553318
rect 542360 550656 542412 550662
rect 542360 550598 542412 550604
rect 542452 550656 542504 550662
rect 542452 550598 542504 550604
rect 542372 543794 542400 550598
rect 542360 543788 542412 543794
rect 542360 543730 542412 543736
rect 542452 543652 542504 543658
rect 542452 543594 542504 543600
rect 542464 534070 542492 543594
rect 542452 534064 542504 534070
rect 542452 534006 542504 534012
rect 542636 534064 542688 534070
rect 542636 534006 542688 534012
rect 542648 524482 542676 534006
rect 542636 524476 542688 524482
rect 542636 524418 542688 524424
rect 542728 524408 542780 524414
rect 542728 524350 542780 524356
rect 542740 521665 542768 524350
rect 542542 521656 542598 521665
rect 542542 521591 542598 521600
rect 542726 521656 542782 521665
rect 542726 521591 542782 521600
rect 542556 512038 542584 521591
rect 542544 512032 542596 512038
rect 542544 511974 542596 511980
rect 542820 512032 542872 512038
rect 542820 511974 542872 511980
rect 542832 502382 542860 511974
rect 542636 502376 542688 502382
rect 542636 502318 542688 502324
rect 542820 502376 542872 502382
rect 542820 502318 542872 502324
rect 542648 492833 542676 502318
rect 542634 492824 542690 492833
rect 542634 492759 542690 492768
rect 542542 492688 542598 492697
rect 542542 492623 542544 492632
rect 542596 492623 542598 492632
rect 542636 492652 542688 492658
rect 542544 492594 542596 492600
rect 542636 492594 542688 492600
rect 542648 485790 542676 492594
rect 542544 485784 542596 485790
rect 542544 485726 542596 485732
rect 542636 485784 542688 485790
rect 542636 485726 542688 485732
rect 542556 483018 542584 485726
rect 542556 482990 542676 483018
rect 542648 476134 542676 482990
rect 542452 476128 542504 476134
rect 542636 476128 542688 476134
rect 542504 476076 542584 476082
rect 542452 476070 542584 476076
rect 542636 476070 542688 476076
rect 542464 476054 542584 476070
rect 542556 473346 542584 476054
rect 542544 473340 542596 473346
rect 542544 473282 542596 473288
rect 542636 473340 542688 473346
rect 542636 473282 542688 473288
rect 542648 466478 542676 473282
rect 542636 466472 542688 466478
rect 542636 466414 542688 466420
rect 542544 466404 542596 466410
rect 542544 466346 542596 466352
rect 542556 463706 542584 466346
rect 542556 463678 542676 463706
rect 542648 454073 542676 463678
rect 542358 454064 542414 454073
rect 542358 453999 542414 454008
rect 542634 454064 542690 454073
rect 542634 453999 542690 454008
rect 542372 447166 542400 453999
rect 542360 447160 542412 447166
rect 542360 447102 542412 447108
rect 542452 447092 542504 447098
rect 542452 447034 542504 447040
rect 542464 444378 542492 447034
rect 542176 444372 542228 444378
rect 542176 444314 542228 444320
rect 542452 444372 542504 444378
rect 542452 444314 542504 444320
rect 542188 434761 542216 444314
rect 542174 434752 542230 434761
rect 542174 434687 542230 434696
rect 542358 434752 542414 434761
rect 542358 434687 542414 434696
rect 542372 427854 542400 434687
rect 542360 427848 542412 427854
rect 542360 427790 542412 427796
rect 542452 427780 542504 427786
rect 542452 427722 542504 427728
rect 542464 425066 542492 427722
rect 542176 425060 542228 425066
rect 542176 425002 542228 425008
rect 542452 425060 542504 425066
rect 542452 425002 542504 425008
rect 542188 415449 542216 425002
rect 542174 415440 542230 415449
rect 542174 415375 542230 415384
rect 542358 415440 542414 415449
rect 542358 415375 542414 415384
rect 542372 408542 542400 415375
rect 542360 408536 542412 408542
rect 542360 408478 542412 408484
rect 542452 408400 542504 408406
rect 542452 408342 542504 408348
rect 542464 404326 542492 408342
rect 542084 404320 542136 404326
rect 542084 404262 542136 404268
rect 542452 404320 542504 404326
rect 542452 404262 542504 404268
rect 542096 394777 542124 404262
rect 542082 394768 542138 394777
rect 542082 394703 542138 394712
rect 542266 394768 542322 394777
rect 542322 394726 542400 394754
rect 542266 394703 542322 394712
rect 542372 393310 542400 394726
rect 542176 393304 542228 393310
rect 542176 393246 542228 393252
rect 542360 393304 542412 393310
rect 542360 393246 542412 393252
rect 542188 383722 542216 393246
rect 542176 383716 542228 383722
rect 542176 383658 542228 383664
rect 542452 383716 542504 383722
rect 542452 383658 542504 383664
rect 542464 379506 542492 383658
rect 542452 379500 542504 379506
rect 542452 379442 542504 379448
rect 542636 379500 542688 379506
rect 542636 379442 542688 379448
rect 542648 371906 542676 379442
rect 542648 371878 542768 371906
rect 542740 367062 542768 371878
rect 542452 367056 542504 367062
rect 542452 366998 542504 367004
rect 542728 367056 542780 367062
rect 542728 366998 542780 367004
rect 542464 357474 542492 366998
rect 542452 357468 542504 357474
rect 542452 357410 542504 357416
rect 542544 357468 542596 357474
rect 542544 357410 542596 357416
rect 542556 350606 542584 357410
rect 542544 350600 542596 350606
rect 542544 350542 542596 350548
rect 542728 350532 542780 350538
rect 542728 350474 542780 350480
rect 542740 340882 542768 350474
rect 542728 340876 542780 340882
rect 542728 340818 542780 340824
rect 545776 332586 545804 696934
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 560944 685908 560996 685914
rect 560944 685850 560996 685856
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 558184 638988 558236 638994
rect 558184 638930 558236 638936
rect 556804 592068 556856 592074
rect 556804 592010 556856 592016
rect 555424 545148 555476 545154
rect 555424 545090 555476 545096
rect 554044 498228 554096 498234
rect 554044 498170 554096 498176
rect 549904 462392 549956 462398
rect 549904 462334 549956 462340
rect 547144 415472 547196 415478
rect 547144 415414 547196 415420
rect 545764 332580 545816 332586
rect 545764 332522 545816 332528
rect 540244 325644 540296 325650
rect 540244 325586 540296 325592
rect 538864 320136 538916 320142
rect 538864 320078 538916 320084
rect 537484 313268 537536 313274
rect 537484 313210 537536 313216
rect 536104 306332 536156 306338
rect 536104 306274 536156 306280
rect 534724 298104 534776 298110
rect 534724 298046 534776 298052
rect 547156 293962 547184 415414
rect 549916 300830 549944 462334
rect 554056 309126 554084 498170
rect 555436 314634 555464 545090
rect 556816 321570 556844 592010
rect 558196 328438 558224 638930
rect 560956 333946 560984 685850
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 563704 451308 563756 451314
rect 563704 451250 563756 451256
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 560944 333940 560996 333946
rect 560944 333882 560996 333888
rect 558184 328432 558236 328438
rect 558184 328374 558236 328380
rect 556804 321564 556856 321570
rect 556804 321506 556856 321512
rect 555424 314628 555476 314634
rect 555424 314570 555476 314576
rect 554044 309120 554096 309126
rect 554044 309062 554096 309068
rect 563716 302190 563744 451250
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 580184 415478 580212 416463
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 580262 404832 580318 404841
rect 580262 404767 580318 404776
rect 579894 393000 579950 393009
rect 579894 392935 579950 392944
rect 579908 392018 579936 392935
rect 579896 392012 579948 392018
rect 579896 391954 579948 391960
rect 563704 302184 563756 302190
rect 563704 302126 563756 302132
rect 549904 300824 549956 300830
rect 549904 300766 549956 300772
rect 579986 299160 580042 299169
rect 579986 299095 580042 299104
rect 580000 294642 580028 299095
rect 580276 296682 580304 404767
rect 580354 369608 580410 369617
rect 580354 369543 580410 369552
rect 580264 296676 580316 296682
rect 580264 296618 580316 296624
rect 579988 294636 580040 294642
rect 579988 294578 580040 294584
rect 547144 293956 547196 293962
rect 547144 293898 547196 293904
rect 522580 292052 522632 292058
rect 522580 291994 522632 292000
rect 523960 292052 524012 292058
rect 523960 291994 524012 292000
rect 522592 291553 522620 291994
rect 522578 291544 522634 291553
rect 522578 291479 522634 291488
rect 522948 289808 523000 289814
rect 522948 289750 523000 289756
rect 522960 289513 522988 289750
rect 522946 289504 523002 289513
rect 522946 289439 523002 289448
rect 580368 288386 580396 369543
rect 580446 357912 580502 357921
rect 580446 357847 580502 357856
rect 580460 289814 580488 357847
rect 580538 346080 580594 346089
rect 580538 346015 580594 346024
rect 580448 289808 580500 289814
rect 580448 289750 580500 289756
rect 522580 288380 522632 288386
rect 522580 288322 522632 288328
rect 580356 288380 580408 288386
rect 580356 288322 580408 288328
rect 522592 287337 522620 288322
rect 522578 287328 522634 287337
rect 522578 287263 522634 287272
rect 580552 285666 580580 346015
rect 580630 322688 580686 322697
rect 580630 322623 580686 322632
rect 522580 285660 522632 285666
rect 522580 285602 522632 285608
rect 580540 285660 580592 285666
rect 580540 285602 580592 285608
rect 522592 285297 522620 285602
rect 522578 285288 522634 285297
rect 522578 285223 522634 285232
rect 522486 283112 522542 283121
rect 522486 283047 522542 283056
rect 580644 281518 580672 322623
rect 580722 310856 580778 310865
rect 580722 310791 580778 310800
rect 580736 294710 580764 310791
rect 580724 294704 580776 294710
rect 580724 294646 580776 294652
rect 522948 281512 523000 281518
rect 522948 281454 523000 281460
rect 580632 281512 580684 281518
rect 580632 281454 580684 281460
rect 522960 281081 522988 281454
rect 522946 281072 523002 281081
rect 522946 281007 523002 281016
rect 522486 276856 522542 276865
rect 522486 276791 522542 276800
rect 522500 265674 522528 276791
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580184 275330 580212 275703
rect 522948 275324 523000 275330
rect 522948 275266 523000 275272
rect 580172 275324 580224 275330
rect 580172 275266 580224 275272
rect 522960 274689 522988 275266
rect 522946 274680 523002 274689
rect 522946 274615 523002 274624
rect 522854 270464 522910 270473
rect 522854 270399 522910 270408
rect 522578 266248 522634 266257
rect 522578 266183 522634 266192
rect 522488 265668 522540 265674
rect 522488 265610 522540 265616
rect 522592 264994 522620 266183
rect 522580 264988 522632 264994
rect 522580 264930 522632 264936
rect 522762 264208 522818 264217
rect 522762 264143 522818 264152
rect 522578 262032 522634 262041
rect 522578 261967 522634 261976
rect 522592 260914 522620 261967
rect 522580 260908 522632 260914
rect 522580 260850 522632 260856
rect 522578 259992 522634 260001
rect 522578 259927 522634 259936
rect 522592 259486 522620 259927
rect 522580 259480 522632 259486
rect 522580 259422 522632 259428
rect 522578 257816 522634 257825
rect 522578 257751 522634 257760
rect 522486 251560 522542 251569
rect 522486 251495 522542 251504
rect 522396 243228 522448 243234
rect 522396 243170 522448 243176
rect 522394 243128 522450 243137
rect 522394 243063 522450 243072
rect 522408 242962 522436 243063
rect 522396 242956 522448 242962
rect 522396 242898 522448 242904
rect 522396 242820 522448 242826
rect 522396 242762 522448 242768
rect 522408 240922 522436 242762
rect 522396 240916 522448 240922
rect 522396 240858 522448 240864
rect 522394 240544 522450 240553
rect 522394 240479 522450 240488
rect 522408 240174 522436 240479
rect 522396 240168 522448 240174
rect 522396 240110 522448 240116
rect 522500 77246 522528 251495
rect 522592 124166 522620 257751
rect 522670 255776 522726 255785
rect 522670 255711 522726 255720
rect 522684 135250 522712 255711
rect 522776 171086 522804 264143
rect 522868 218006 522896 270399
rect 522946 268424 523002 268433
rect 522946 268359 523002 268368
rect 522960 229090 522988 268359
rect 580172 265668 580224 265674
rect 580172 265610 580224 265616
rect 523960 264988 524012 264994
rect 523960 264930 524012 264936
rect 523868 260908 523920 260914
rect 523868 260850 523920 260856
rect 523776 259480 523828 259486
rect 523776 259422 523828 259428
rect 523682 253600 523738 253609
rect 523682 253535 523738 253544
rect 522948 229084 523000 229090
rect 522948 229026 523000 229032
rect 522856 218000 522908 218006
rect 522856 217942 522908 217948
rect 522764 171080 522816 171086
rect 522764 171022 522816 171028
rect 522672 135244 522724 135250
rect 522672 135186 522724 135192
rect 522580 124160 522632 124166
rect 522580 124102 522632 124108
rect 523696 111790 523724 253535
rect 523788 158710 523816 259422
rect 523880 182170 523908 260850
rect 523972 205630 524000 264930
rect 580184 263945 580212 265610
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 531964 248464 532016 248470
rect 531964 248406 532016 248412
rect 527824 247104 527876 247110
rect 527824 247046 527876 247052
rect 525064 240168 525116 240174
rect 525064 240110 525116 240116
rect 523960 205624 524012 205630
rect 523960 205566 524012 205572
rect 523868 182164 523920 182170
rect 523868 182106 523920 182112
rect 523776 158704 523828 158710
rect 523776 158646 523828 158652
rect 523684 111784 523736 111790
rect 523684 111726 523736 111732
rect 522488 77240 522540 77246
rect 522488 77182 522540 77188
rect 522304 30320 522356 30326
rect 522304 30262 522356 30268
rect 525076 17950 525104 240110
rect 527836 64870 527864 247046
rect 529204 242956 529256 242962
rect 529204 242898 529256 242904
rect 527824 64864 527876 64870
rect 527824 64806 527876 64812
rect 529216 41410 529244 242898
rect 531976 88330 532004 248406
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 531964 88324 532016 88330
rect 531964 88266 532016 88272
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 529204 41404 529256 41410
rect 529204 41346 529256 41352
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 525064 17944 525116 17950
rect 525064 17886 525116 17892
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 522120 8288 522172 8294
rect 522120 8230 522172 8236
rect 142068 2848 142120 2854
rect 142068 2790 142120 2796
rect 145656 2848 145708 2854
rect 145656 2790 145708 2796
rect 149244 2848 149296 2854
rect 149244 2790 149296 2796
rect 152740 2848 152792 2854
rect 152740 2790 152792 2796
rect 156328 2848 156380 2854
rect 156328 2790 156380 2796
rect 159916 2848 159968 2854
rect 159916 2790 159968 2796
rect 163504 2848 163556 2854
rect 163504 2790 163556 2796
rect 167092 2848 167144 2854
rect 167092 2790 167144 2796
rect 170588 2848 170640 2854
rect 170588 2790 170640 2796
rect 174176 2848 174228 2854
rect 174176 2790 174228 2796
rect 177764 2848 177816 2854
rect 177764 2790 177816 2796
rect 181352 2848 181404 2854
rect 181352 2790 181404 2796
rect 184848 2848 184900 2854
rect 184848 2790 184900 2796
rect 188436 2848 188488 2854
rect 188436 2790 188488 2796
rect 192024 2848 192076 2854
rect 192024 2790 192076 2796
rect 195612 2848 195664 2854
rect 195612 2790 195664 2796
rect 199200 2848 199252 2854
rect 199200 2790 199252 2796
rect 202696 2848 202748 2854
rect 202696 2790 202748 2796
rect 206284 2848 206336 2854
rect 206284 2790 206336 2796
rect 209872 2848 209924 2854
rect 209872 2790 209924 2796
rect 213460 2848 213512 2854
rect 213460 2790 213512 2796
rect 217048 2848 217100 2854
rect 217048 2790 217100 2796
rect 220544 2848 220596 2854
rect 220544 2790 220596 2796
rect 224132 2848 224184 2854
rect 224132 2790 224184 2796
rect 227720 2848 227772 2854
rect 227720 2790 227772 2796
rect 231308 2848 231360 2854
rect 231308 2790 231360 2796
rect 234804 2848 234856 2854
rect 234804 2790 234856 2796
rect 238392 2848 238444 2854
rect 238392 2790 238444 2796
rect 241980 2848 242032 2854
rect 241980 2790 242032 2796
rect 245568 2848 245620 2854
rect 245568 2790 245620 2796
rect 249156 2848 249208 2854
rect 249156 2790 249208 2796
rect 252652 2848 252704 2854
rect 252652 2790 252704 2796
rect 256240 2848 256292 2854
rect 256240 2790 256292 2796
rect 259828 2848 259880 2854
rect 259828 2790 259880 2796
rect 263416 2848 263468 2854
rect 263416 2790 263468 2796
rect 267004 2848 267056 2854
rect 267004 2790 267056 2796
rect 270500 2848 270552 2854
rect 270500 2790 270552 2796
rect 274088 2848 274140 2854
rect 274088 2790 274140 2796
rect 277676 2848 277728 2854
rect 277676 2790 277728 2796
rect 281264 2848 281316 2854
rect 281264 2790 281316 2796
rect 284760 2848 284812 2854
rect 284760 2790 284812 2796
rect 288348 2848 288400 2854
rect 288348 2790 288400 2796
rect 291936 2848 291988 2854
rect 291936 2790 291988 2796
rect 295524 2848 295576 2854
rect 295524 2790 295576 2796
rect 299112 2848 299164 2854
rect 299112 2790 299164 2796
rect 302608 2848 302660 2854
rect 302608 2790 302660 2796
rect 305644 2848 305696 2854
rect 305644 2790 305696 2796
rect 306196 2848 306248 2854
rect 306196 2790 306248 2796
rect 309784 2848 309836 2854
rect 309784 2790 309836 2796
rect 313372 2848 313424 2854
rect 313372 2790 313424 2796
rect 316960 2848 317012 2854
rect 316960 2790 317012 2796
rect 320456 2848 320508 2854
rect 320456 2790 320508 2796
rect 324044 2848 324096 2854
rect 324044 2790 324096 2796
rect 327632 2848 327684 2854
rect 327632 2790 327684 2796
rect 331220 2848 331272 2854
rect 331220 2790 331272 2796
rect 334716 2848 334768 2854
rect 334716 2790 334768 2796
rect 338304 2848 338356 2854
rect 338304 2790 338356 2796
rect 341892 2848 341944 2854
rect 341892 2790 341944 2796
rect 345480 2848 345532 2854
rect 345480 2790 345532 2796
rect 349068 2848 349120 2854
rect 349068 2790 349120 2796
rect 352564 2848 352616 2854
rect 352564 2790 352616 2796
rect 356152 2848 356204 2854
rect 356152 2790 356204 2796
rect 359740 2848 359792 2854
rect 359740 2790 359792 2796
rect 363328 2848 363380 2854
rect 363328 2790 363380 2796
rect 366916 2848 366968 2854
rect 366916 2790 366968 2796
rect 370412 2848 370464 2854
rect 370412 2790 370464 2796
rect 374000 2848 374052 2854
rect 374000 2790 374052 2796
rect 377588 2848 377640 2854
rect 377588 2790 377640 2796
rect 381176 2848 381228 2854
rect 381176 2790 381228 2796
rect 384672 2848 384724 2854
rect 384672 2790 384724 2796
rect 388260 2848 388312 2854
rect 388260 2790 388312 2796
rect 391848 2848 391900 2854
rect 391848 2790 391900 2796
rect 395436 2848 395488 2854
rect 395436 2790 395488 2796
rect 399024 2848 399076 2854
rect 399024 2790 399076 2796
rect 402520 2848 402572 2854
rect 402520 2790 402572 2796
rect 406108 2848 406160 2854
rect 406108 2790 406160 2796
rect 409696 2848 409748 2854
rect 409696 2790 409748 2796
rect 413284 2848 413336 2854
rect 413284 2790 413336 2796
rect 416872 2848 416924 2854
rect 416872 2790 416924 2796
rect 420368 2848 420420 2854
rect 420368 2790 420420 2796
rect 423956 2848 424008 2854
rect 423956 2790 424008 2796
rect 427544 2848 427596 2854
rect 427544 2790 427596 2796
rect 431132 2848 431184 2854
rect 431132 2790 431184 2796
rect 434628 2848 434680 2854
rect 434628 2790 434680 2796
rect 438216 2848 438268 2854
rect 438216 2790 438268 2796
rect 441804 2848 441856 2854
rect 441804 2790 441856 2796
rect 445392 2848 445444 2854
rect 445392 2790 445444 2796
rect 448980 2848 449032 2854
rect 448980 2790 449032 2796
rect 452476 2848 452528 2854
rect 452476 2790 452528 2796
rect 456064 2848 456116 2854
rect 456064 2790 456116 2796
rect 459652 2848 459704 2854
rect 459652 2790 459704 2796
rect 463240 2848 463292 2854
rect 463240 2790 463292 2796
rect 466828 2848 466880 2854
rect 466828 2790 466880 2796
rect 470324 2848 470376 2854
rect 470324 2790 470376 2796
rect 473912 2848 473964 2854
rect 473912 2790 473964 2796
rect 477500 2848 477552 2854
rect 477500 2790 477552 2796
rect 481088 2848 481140 2854
rect 481088 2790 481140 2796
rect 484584 2848 484636 2854
rect 484584 2790 484636 2796
rect 488172 2848 488224 2854
rect 488172 2790 488224 2796
rect 491760 2848 491812 2854
rect 491760 2790 491812 2796
rect 495348 2848 495400 2854
rect 495348 2790 495400 2796
rect 498936 2848 498988 2854
rect 498936 2790 498988 2796
rect 502432 2848 502484 2854
rect 502432 2790 502484 2796
rect 506020 2848 506072 2854
rect 506020 2790 506072 2796
rect 509608 2848 509660 2854
rect 509608 2790 509660 2796
rect 513196 2848 513248 2854
rect 513196 2790 513248 2796
rect 516784 2848 516836 2854
rect 516784 2790 516836 2796
rect 520280 2848 520332 2854
rect 520280 2790 520332 2796
rect 523868 2848 523920 2854
rect 523868 2790 523920 2796
rect 527456 2848 527508 2854
rect 527456 2790 527508 2796
rect 531044 2848 531096 2854
rect 531044 2790 531096 2796
rect 534540 2848 534592 2854
rect 534540 2790 534592 2796
rect 538128 2848 538180 2854
rect 538128 2790 538180 2796
rect 541716 2848 541768 2854
rect 541716 2790 541768 2796
rect 545304 2848 545356 2854
rect 545304 2790 545356 2796
rect 548892 2848 548944 2854
rect 548892 2790 548944 2796
rect 552388 2848 552440 2854
rect 552388 2790 552440 2796
rect 555976 2848 556028 2854
rect 555976 2790 556028 2796
rect 559564 2848 559616 2854
rect 559564 2790 559616 2796
rect 563152 2848 563204 2854
rect 563152 2790 563204 2796
rect 566740 2848 566792 2854
rect 566740 2790 566792 2796
rect 570236 2848 570288 2854
rect 570236 2790 570288 2796
rect 573824 2848 573876 2854
rect 573824 2790 573876 2796
rect 577412 2848 577464 2854
rect 577412 2790 577464 2796
rect 581000 2848 581052 2854
rect 581000 2790 581052 2796
rect 134904 598 135208 626
rect 142080 610 142108 2790
rect 138480 604 138532 610
rect 134904 480 134932 598
rect 138480 546 138532 552
rect 142068 604 142120 610
rect 142068 546 142120 552
rect 138492 480 138520 546
rect 142080 480 142108 546
rect 145668 480 145696 2790
rect 149256 480 149284 2790
rect 152752 480 152780 2790
rect 156340 480 156368 2790
rect 159928 480 159956 2790
rect 163516 480 163544 2790
rect 167104 480 167132 2790
rect 170600 480 170628 2790
rect 174188 480 174216 2790
rect 177776 480 177804 2790
rect 181364 480 181392 2790
rect 184860 480 184888 2790
rect 188448 480 188476 2790
rect 192036 480 192064 2790
rect 195624 480 195652 2790
rect 199212 480 199240 2790
rect 202708 480 202736 2790
rect 206296 480 206324 2790
rect 209884 480 209912 2790
rect 213472 480 213500 2790
rect 217060 480 217088 2790
rect 220556 480 220584 2790
rect 224144 480 224172 2790
rect 227732 480 227760 2790
rect 231320 480 231348 2790
rect 234816 480 234844 2790
rect 238404 480 238432 2790
rect 241992 480 242020 2790
rect 245580 480 245608 2790
rect 249168 480 249196 2790
rect 252664 480 252692 2790
rect 256252 480 256280 2790
rect 259840 480 259868 2790
rect 263428 480 263456 2790
rect 267016 480 267044 2790
rect 270512 480 270540 2790
rect 274100 480 274128 2790
rect 277688 480 277716 2790
rect 281276 480 281304 2790
rect 284772 480 284800 2790
rect 288360 480 288388 2790
rect 291948 480 291976 2790
rect 295536 480 295564 2790
rect 299124 480 299152 2790
rect 302620 480 302648 2790
rect 306208 480 306236 2790
rect 309796 480 309824 2790
rect 313384 480 313412 2790
rect 316972 480 317000 2790
rect 320468 480 320496 2790
rect 324056 480 324084 2790
rect 327644 480 327672 2790
rect 331232 480 331260 2790
rect 334728 480 334756 2790
rect 338316 480 338344 2790
rect 341904 480 341932 2790
rect 345492 480 345520 2790
rect 349080 480 349108 2790
rect 352576 480 352604 2790
rect 356164 480 356192 2790
rect 359752 480 359780 2790
rect 363340 480 363368 2790
rect 366928 480 366956 2790
rect 370424 480 370452 2790
rect 374012 480 374040 2790
rect 377600 480 377628 2790
rect 381188 480 381216 2790
rect 384684 480 384712 2790
rect 388272 480 388300 2790
rect 391860 480 391888 2790
rect 395448 480 395476 2790
rect 399036 480 399064 2790
rect 402532 480 402560 2790
rect 406120 480 406148 2790
rect 409708 480 409736 2790
rect 413296 480 413324 2790
rect 416884 480 416912 2790
rect 420380 480 420408 2790
rect 423968 480 423996 2790
rect 427556 480 427584 2790
rect 431144 480 431172 2790
rect 434640 480 434668 2790
rect 438228 480 438256 2790
rect 441816 480 441844 2790
rect 445404 480 445432 2790
rect 448992 480 449020 2790
rect 452488 480 452516 2790
rect 456076 480 456104 2790
rect 459664 480 459692 2790
rect 463252 480 463280 2790
rect 466840 480 466868 2790
rect 470336 480 470364 2790
rect 473924 480 473952 2790
rect 477512 480 477540 2790
rect 481100 480 481128 2790
rect 484596 480 484624 2790
rect 488184 480 488212 2790
rect 491772 480 491800 2790
rect 495360 480 495388 2790
rect 498948 480 498976 2790
rect 502444 480 502472 2790
rect 506032 480 506060 2790
rect 509620 480 509648 2790
rect 513208 480 513236 2790
rect 516796 480 516824 2790
rect 520292 480 520320 2790
rect 523880 480 523908 2790
rect 527468 480 527496 2790
rect 531056 480 531084 2790
rect 534552 480 534580 2790
rect 538140 480 538168 2790
rect 541728 480 541756 2790
rect 545316 480 545344 2790
rect 548904 480 548932 2790
rect 552400 480 552428 2790
rect 555988 480 556016 2790
rect 559576 480 559604 2790
rect 563164 480 563192 2790
rect 566752 480 566780 2790
rect 570248 480 570276 2790
rect 573836 480 573864 2790
rect 577424 480 577452 2790
rect 581012 480 581040 2790
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 24306 700440 24362 700496
rect 89166 700712 89222 700768
rect 72974 700576 73030 700632
rect 8114 700304 8170 700360
rect 3330 653520 3386 653576
rect 3330 652840 3386 652896
rect 3422 624824 3478 624880
rect 3422 623736 3478 623792
rect 3422 610408 3478 610464
rect 3514 595992 3570 596048
rect 3330 509904 3386 509960
rect 3422 495508 3478 495544
rect 3422 495488 3424 495508
rect 3424 495488 3476 495508
rect 3476 495488 3478 495508
rect 2962 481072 3018 481128
rect 3238 423680 3294 423736
rect 3146 394984 3202 395040
rect 3330 308760 3386 308816
rect 3054 294344 3110 294400
rect 3146 222536 3202 222592
rect 2962 193840 3018 193896
rect 3330 50904 3386 50960
rect 3330 50088 3386 50144
rect 3606 567296 3662 567352
rect 3698 553016 3754 553072
rect 3790 538600 3846 538656
rect 71318 479848 71374 479904
rect 61842 479576 61898 479632
rect 71318 479576 71374 479632
rect 298006 606600 298062 606656
rect 297914 605376 297970 605432
rect 297822 603744 297878 603800
rect 297730 602520 297786 602576
rect 297638 600888 297694 600944
rect 297546 599800 297602 599856
rect 297454 598032 297510 598088
rect 297362 540232 297418 540288
rect 297270 538464 297326 538520
rect 50986 479460 51042 479496
rect 50986 479440 50988 479460
rect 50988 479440 51040 479460
rect 51040 479440 51042 479460
rect 41326 479304 41382 479360
rect 57794 479304 57850 479360
rect 57978 479324 58034 479360
rect 108946 479576 109002 479632
rect 109130 479576 109186 479632
rect 99378 479440 99434 479496
rect 57978 479304 57980 479324
rect 57980 479304 58032 479324
rect 58032 479304 58034 479324
rect 135166 479460 135222 479496
rect 135166 479440 135168 479460
rect 135168 479440 135220 479460
rect 135220 479440 135222 479460
rect 154486 479440 154542 479496
rect 173806 479440 173862 479496
rect 193126 479440 193182 479496
rect 212446 479440 212502 479496
rect 231766 479440 231822 479496
rect 251086 479440 251142 479496
rect 278778 479440 278834 479496
rect 128266 479304 128322 479360
rect 147586 479340 147588 479360
rect 147588 479340 147640 479360
rect 147640 479340 147642 479360
rect 147586 479304 147642 479340
rect 166906 479340 166908 479360
rect 166908 479340 166960 479360
rect 166960 479340 166962 479360
rect 166906 479304 166962 479340
rect 186226 479340 186228 479360
rect 186228 479340 186280 479360
rect 186280 479340 186282 479360
rect 186226 479304 186282 479340
rect 205546 479340 205548 479360
rect 205548 479340 205600 479360
rect 205600 479340 205602 479360
rect 205546 479304 205602 479340
rect 224866 479340 224868 479360
rect 224868 479340 224920 479360
rect 224920 479340 224922 479360
rect 224866 479304 224922 479340
rect 244186 479340 244188 479360
rect 244188 479340 244240 479360
rect 244240 479340 244242 479360
rect 244186 479304 244242 479340
rect 99470 479168 99526 479224
rect 277398 478932 277400 478952
rect 277400 478932 277452 478952
rect 277452 478932 277454 478952
rect 3514 452376 3570 452432
rect 3514 437960 3570 438016
rect 3514 380568 3570 380624
rect 3514 366152 3570 366208
rect 3514 337456 3570 337512
rect 3514 323040 3570 323096
rect 3514 280100 3516 280120
rect 3516 280100 3568 280120
rect 3568 280100 3570 280120
rect 3514 280064 3570 280100
rect 3514 265648 3570 265704
rect 3606 251232 3662 251288
rect 3514 236952 3570 237008
rect 3514 208120 3570 208176
rect 3514 200640 3570 200696
rect 3698 200776 3754 200832
rect 3606 150728 3662 150784
rect 3882 179424 3938 179480
rect 3790 165008 3846 165064
rect 3698 136312 3754 136368
rect 3514 122032 3570 122088
rect 3514 108840 3570 108896
rect 3514 107616 3570 107672
rect 3514 80008 3570 80064
rect 3514 78920 3570 78976
rect 3422 21392 3478 21448
rect 3422 7112 3478 7168
rect 277398 478896 277454 478932
rect 277398 476720 277454 476776
rect 278686 474680 278742 474736
rect 278686 472504 278742 472560
rect 277858 470328 277914 470384
rect 278686 468288 278742 468344
rect 278686 466112 278742 466168
rect 278686 464072 278742 464128
rect 278686 461896 278742 461952
rect 278686 459720 278742 459776
rect 278686 457680 278742 457736
rect 278686 455504 278742 455560
rect 278686 453328 278742 453384
rect 278686 451308 278742 451344
rect 278686 451288 278688 451308
rect 278688 451288 278740 451308
rect 278740 451288 278742 451308
rect 278686 449112 278742 449168
rect 278686 447072 278742 447128
rect 278686 444896 278742 444952
rect 277858 442720 277914 442776
rect 278686 440680 278742 440736
rect 278686 438504 278742 438560
rect 278042 436328 278098 436384
rect 278686 434288 278742 434344
rect 278686 432112 278742 432168
rect 277674 430072 277730 430128
rect 278686 427896 278742 427952
rect 278686 425720 278742 425776
rect 278686 423700 278742 423736
rect 278686 423680 278688 423700
rect 278688 423680 278740 423700
rect 278740 423680 278742 423700
rect 278686 421504 278742 421560
rect 278686 419464 278742 419520
rect 278686 417288 278742 417344
rect 277858 415112 277914 415168
rect 278686 413072 278742 413128
rect 278686 410896 278742 410952
rect 278686 408720 278742 408776
rect 278686 406680 278742 406736
rect 278686 404504 278742 404560
rect 278410 402464 278466 402520
rect 278686 400288 278742 400344
rect 278686 398112 278742 398168
rect 278686 396092 278742 396128
rect 278686 396072 278688 396092
rect 278688 396072 278740 396092
rect 278740 396072 278742 396092
rect 278686 393896 278742 393952
rect 278318 391720 278374 391776
rect 278686 389680 278742 389736
rect 277858 387504 277914 387560
rect 277674 385464 277730 385520
rect 278686 383288 278742 383344
rect 278042 381112 278098 381168
rect 278686 379072 278742 379128
rect 278686 376896 278742 376952
rect 278410 374856 278466 374912
rect 278042 372680 278098 372736
rect 278318 370504 278374 370560
rect 278686 368500 278688 368520
rect 278688 368500 278740 368520
rect 278740 368500 278742 368520
rect 278686 368464 278742 368500
rect 278686 366288 278742 366344
rect 277858 364112 277914 364168
rect 278686 362072 278742 362128
rect 277858 359896 277914 359952
rect 278686 357856 278742 357912
rect 278686 355680 278742 355736
rect 278042 353504 278098 353560
rect 278686 351464 278742 351520
rect 278686 349288 278742 349344
rect 278686 347112 278742 347168
rect 278686 345092 278742 345128
rect 278686 345072 278688 345092
rect 278688 345072 278740 345092
rect 278740 345072 278742 345092
rect 278318 342896 278374 342952
rect 278686 340892 278688 340912
rect 278688 340892 278740 340912
rect 278740 340892 278742 340912
rect 278686 340856 278742 340892
rect 278686 338680 278742 338736
rect 277858 336504 277914 336560
rect 278686 334464 278742 334520
rect 278686 332288 278742 332344
rect 278686 330248 278742 330304
rect 278686 328072 278742 328128
rect 278042 325896 278098 325952
rect 277674 323856 277730 323912
rect 278042 321680 278098 321736
rect 278686 319504 278742 319560
rect 278686 317484 278742 317520
rect 278686 317464 278688 317484
rect 278688 317464 278740 317484
rect 278740 317464 278742 317484
rect 278686 315288 278742 315344
rect 278686 313284 278688 313304
rect 278688 313284 278740 313304
rect 278740 313284 278742 313304
rect 278686 313248 278742 313284
rect 278686 311072 278742 311128
rect 277858 308896 277914 308952
rect 278686 306856 278742 306912
rect 278686 304680 278742 304736
rect 278686 302504 278742 302560
rect 278686 300464 278742 300520
rect 278686 298288 278742 298344
rect 278686 296248 278742 296304
rect 278686 294072 278742 294128
rect 278686 291896 278742 291952
rect 278686 289876 278742 289912
rect 278686 289856 278688 289876
rect 278688 289856 278740 289876
rect 278740 289856 278742 289876
rect 278686 287680 278742 287736
rect 278686 285676 278688 285696
rect 278688 285676 278740 285696
rect 278740 285676 278742 285696
rect 278686 285640 278742 285676
rect 278686 283464 278742 283520
rect 277858 281288 277914 281344
rect 278686 279248 278742 279304
rect 278686 277072 278742 277128
rect 278042 274896 278098 274952
rect 278686 272856 278742 272912
rect 278686 270680 278742 270736
rect 278686 268640 278742 268696
rect 278042 266464 278098 266520
rect 278686 264288 278742 264344
rect 278686 262268 278742 262304
rect 278686 262248 278688 262268
rect 278688 262248 278740 262268
rect 278740 262248 278742 262268
rect 278318 260072 278374 260128
rect 277858 257896 277914 257952
rect 278686 255856 278742 255912
rect 277858 253680 277914 253736
rect 278686 251640 278742 251696
rect 278686 249464 278742 249520
rect 278042 247288 278098 247344
rect 277398 243072 277454 243128
rect 278134 245248 278190 245304
rect 278686 241032 278742 241088
rect 280158 240760 280214 240816
rect 373630 612756 373632 612776
rect 373632 612756 373684 612776
rect 373684 612756 373686 612776
rect 373630 612720 373686 612756
rect 314566 518744 314622 518800
rect 317326 518780 317328 518800
rect 317328 518780 317380 518800
rect 317380 518780 317382 518800
rect 317326 518744 317382 518780
rect 318706 518744 318762 518800
rect 321742 518744 321798 518800
rect 323122 518744 323178 518800
rect 324318 518764 324374 518800
rect 324318 518744 324320 518764
rect 324320 518744 324372 518764
rect 324372 518744 324374 518764
rect 303618 518220 303674 518256
rect 303618 518200 303620 518220
rect 303620 518200 303672 518220
rect 303672 518200 303674 518220
rect 315946 518608 316002 518664
rect 317326 518608 317382 518664
rect 320086 518628 320142 518664
rect 320086 518608 320088 518628
rect 320088 518608 320140 518628
rect 320140 518608 320142 518628
rect 316038 518472 316094 518528
rect 317510 518472 317566 518528
rect 313186 518336 313242 518392
rect 317418 518356 317474 518392
rect 317418 518336 317420 518356
rect 317420 518336 317472 518356
rect 317472 518336 317474 518356
rect 314658 518200 314714 518256
rect 312082 517928 312138 517984
rect 310334 517656 310390 517712
rect 307666 517520 307722 517576
rect 309046 517520 309102 517576
rect 310242 517520 310298 517576
rect 313278 517676 313334 517712
rect 313278 517656 313280 517676
rect 313280 517656 313332 517676
rect 313332 517656 313334 517676
rect 311714 517520 311770 517576
rect 321098 518356 321154 518392
rect 321098 518336 321100 518356
rect 321100 518336 321152 518356
rect 321152 518336 321154 518356
rect 325422 518780 325424 518800
rect 325424 518780 325476 518800
rect 325476 518780 325478 518800
rect 325422 518744 325478 518780
rect 326434 518764 326490 518800
rect 326434 518744 326436 518764
rect 326436 518744 326488 518764
rect 326488 518744 326490 518764
rect 324410 518608 324466 518664
rect 327170 518744 327226 518800
rect 328918 518744 328974 518800
rect 330114 518744 330170 518800
rect 327078 518472 327134 518528
rect 322938 518200 322994 518256
rect 318798 518064 318854 518120
rect 321834 518084 321890 518120
rect 321834 518064 321836 518084
rect 321836 518064 321888 518084
rect 321888 518064 321890 518084
rect 332322 518744 332378 518800
rect 335542 518764 335598 518800
rect 335542 518744 335544 518764
rect 335544 518744 335596 518764
rect 335596 518744 335598 518764
rect 336738 518744 336794 518800
rect 337198 518744 337254 518800
rect 339958 518744 340014 518800
rect 340510 518780 340512 518800
rect 340512 518780 340564 518800
rect 340564 518780 340566 518800
rect 340510 518744 340566 518780
rect 341614 518744 341670 518800
rect 342994 518744 343050 518800
rect 344190 518744 344246 518800
rect 345478 518764 345534 518800
rect 345478 518744 345480 518764
rect 345480 518744 345532 518764
rect 345532 518744 345534 518764
rect 331218 518608 331274 518664
rect 333426 518472 333482 518528
rect 334162 518492 334218 518528
rect 338118 518608 338174 518664
rect 334162 518472 334164 518492
rect 334164 518472 334216 518492
rect 334216 518472 334218 518492
rect 331218 517948 331274 517984
rect 331218 517928 331220 517948
rect 331220 517928 331272 517948
rect 331272 517928 331274 517948
rect 332598 517928 332654 517984
rect 320178 517812 320234 517848
rect 320178 517792 320180 517812
rect 320180 517792 320232 517812
rect 320232 517792 320234 517812
rect 333978 517792 334034 517848
rect 324318 517676 324374 517712
rect 324318 517656 324320 517676
rect 324320 517656 324372 517676
rect 324372 517656 324374 517676
rect 325698 517540 325754 517576
rect 325698 517520 325700 517540
rect 325700 517520 325752 517540
rect 325752 517520 325754 517540
rect 329838 517676 329894 517712
rect 329838 517656 329840 517676
rect 329840 517656 329892 517676
rect 329892 517656 329894 517676
rect 332598 517656 332654 517712
rect 335726 517676 335782 517712
rect 335726 517656 335728 517676
rect 335728 517656 335780 517676
rect 335780 517656 335782 517676
rect 328458 517540 328514 517576
rect 328458 517520 328460 517540
rect 328460 517520 328512 517540
rect 328512 517520 328514 517540
rect 338118 517656 338174 517712
rect 339498 517656 339554 517712
rect 336738 517540 336794 517576
rect 336738 517520 336740 517540
rect 336740 517520 336792 517540
rect 336792 517520 336794 517540
rect 339406 517520 339462 517576
rect 346490 518744 346546 518800
rect 347686 518744 347742 518800
rect 348606 518744 348662 518800
rect 342902 517656 342958 517712
rect 344282 517656 344338 517712
rect 340786 517520 340842 517576
rect 346306 517656 346362 517712
rect 348422 517656 348478 517712
rect 348974 517656 349030 517712
rect 349066 517520 349122 517576
rect 362222 479984 362278 480040
rect 369950 479984 370006 480040
rect 379702 609592 379758 609648
rect 379978 609592 380034 609648
rect 379610 549344 379666 549400
rect 379794 540912 379850 540968
rect 514850 700304 514906 700360
rect 488538 612756 488540 612776
rect 488540 612756 488592 612776
rect 488592 612756 488594 612776
rect 488538 612720 488594 612756
rect 493966 612756 493968 612776
rect 493968 612756 494020 612776
rect 494020 612756 494022 612776
rect 493966 612720 494022 612756
rect 514850 695680 514906 695736
rect 496450 609864 496506 609920
rect 416778 606056 416834 606112
rect 416778 604832 416834 604888
rect 416778 603200 416834 603256
rect 416778 601976 416834 602032
rect 416778 600480 416834 600536
rect 416778 599256 416834 599312
rect 416778 597624 416834 597680
rect 499578 549480 499634 549536
rect 499578 542000 499634 542056
rect 499578 540912 499634 540968
rect 416778 539688 416834 539744
rect 416778 538328 416834 538384
rect 425610 519696 425666 519752
rect 423678 518220 423734 518256
rect 423678 518200 423680 518220
rect 423680 518200 423732 518220
rect 423732 518200 423734 518220
rect 443182 518764 443238 518800
rect 443182 518744 443184 518764
rect 443184 518744 443236 518764
rect 443236 518744 443238 518764
rect 451278 518780 451280 518800
rect 451280 518780 451332 518800
rect 451332 518780 451334 518800
rect 451278 518744 451334 518780
rect 452566 518764 452622 518800
rect 452566 518744 452568 518764
rect 452568 518744 452620 518764
rect 452620 518744 452622 518764
rect 429290 518608 429346 518664
rect 426438 518472 426494 518528
rect 430578 518356 430634 518392
rect 430578 518336 430580 518356
rect 430580 518336 430632 518356
rect 430632 518336 430634 518356
rect 429198 518200 429254 518256
rect 362222 479712 362278 479768
rect 367098 479712 367154 479768
rect 316774 479576 316830 479632
rect 435362 518064 435418 518120
rect 435914 518084 435970 518120
rect 435914 518064 435916 518084
rect 435916 518064 435968 518084
rect 435968 518064 435970 518084
rect 432602 517792 432658 517848
rect 433890 517828 433892 517848
rect 433892 517828 433944 517848
rect 433944 517828 433946 517848
rect 433890 517792 433946 517828
rect 433246 517656 433302 517712
rect 434626 517656 434682 517712
rect 433614 482976 433670 483032
rect 433798 482976 433854 483032
rect 437294 517948 437350 517984
rect 437294 517928 437296 517948
rect 437296 517928 437348 517948
rect 437348 517928 437350 517948
rect 436006 517656 436062 517712
rect 436650 517656 436706 517712
rect 440882 517792 440938 517848
rect 437386 517656 437442 517712
rect 438674 517656 438730 517712
rect 438122 517520 438178 517576
rect 439502 517676 439558 517712
rect 439502 517656 439504 517676
rect 439504 517656 439556 517676
rect 439556 517656 439558 517676
rect 438766 517520 438822 517576
rect 440146 517520 440202 517576
rect 441526 517520 441582 517576
rect 442078 518336 442134 518392
rect 442906 517520 442962 517576
rect 445390 518472 445446 518528
rect 444286 518336 444342 518392
rect 445666 517656 445722 517712
rect 444286 517520 444342 517576
rect 445574 517520 445630 517576
rect 446586 518472 446642 518528
rect 447414 518508 447416 518528
rect 447416 518508 447468 518528
rect 447468 518508 447470 518528
rect 447414 518472 447470 518508
rect 447046 517520 447102 517576
rect 448794 518336 448850 518392
rect 449898 518356 449954 518392
rect 449898 518336 449900 518356
rect 449900 518336 449952 518356
rect 449952 518336 449954 518356
rect 453670 518744 453726 518800
rect 459558 518780 459560 518800
rect 459560 518780 459612 518800
rect 459612 518780 459614 518800
rect 459558 518744 459614 518780
rect 460938 518764 460994 518800
rect 460938 518744 460940 518764
rect 460940 518744 460992 518764
rect 460992 518744 460994 518764
rect 462318 518744 462374 518800
rect 455326 518608 455382 518664
rect 456062 518628 456118 518664
rect 456062 518608 456064 518628
rect 456064 518608 456116 518628
rect 456116 518608 456118 518628
rect 456890 518608 456946 518664
rect 458270 518608 458326 518664
rect 459558 518608 459614 518664
rect 465078 518628 465134 518664
rect 465078 518608 465080 518628
rect 465080 518608 465132 518628
rect 465132 518608 465134 518628
rect 466550 518608 466606 518664
rect 466458 518472 466514 518528
rect 463698 518336 463754 518392
rect 467838 518356 467894 518392
rect 467838 518336 467840 518356
rect 467840 518336 467892 518356
rect 467892 518336 467894 518356
rect 453946 517656 454002 517712
rect 460846 517656 460902 517712
rect 469126 517656 469182 517712
rect 448426 517520 448482 517576
rect 449806 517520 449862 517576
rect 451186 517520 451242 517576
rect 452566 517520 452622 517576
rect 453854 517520 453910 517576
rect 455326 517520 455382 517576
rect 456706 517520 456762 517576
rect 458086 517520 458142 517576
rect 459466 517520 459522 517576
rect 460754 517520 460810 517576
rect 462226 517520 462282 517576
rect 463606 517520 463662 517576
rect 464986 517520 465042 517576
rect 466366 517520 466422 517576
rect 467746 517520 467802 517576
rect 469034 517520 469090 517576
rect 463606 482432 463662 482488
rect 467746 482296 467802 482352
rect 469034 482160 469090 482216
rect 507490 482432 507546 482488
rect 514114 482296 514170 482352
rect 518530 482160 518586 482216
rect 444286 479712 444342 479768
rect 283562 479460 283618 479496
rect 283562 479440 283564 479460
rect 283564 479440 283616 479460
rect 283616 479440 283618 479460
rect 309138 479324 309194 479360
rect 466366 479576 466422 479632
rect 507122 479576 507178 479632
rect 427818 479440 427874 479496
rect 444286 479440 444342 479496
rect 473266 479460 473322 479496
rect 473266 479440 473268 479460
rect 473268 479440 473320 479460
rect 473320 479440 473322 479460
rect 492586 479440 492642 479496
rect 309138 479304 309140 479324
rect 309140 479304 309192 479324
rect 309192 479304 309194 479324
rect 321374 479304 321430 479360
rect 321558 479304 321614 479360
rect 350446 479304 350502 479360
rect 350630 479304 350686 479360
rect 427726 479304 427782 479360
rect 485686 479340 485688 479360
rect 485688 479340 485740 479360
rect 485740 479340 485742 479360
rect 485686 479304 485742 479340
rect 507122 479304 507178 479360
rect 519634 695272 519690 695328
rect 519634 686024 519690 686080
rect 519910 684256 519966 684312
rect 519910 666576 519966 666632
rect 519542 376216 519598 376272
rect 519450 372000 519506 372056
rect 519358 369688 519414 369744
rect 519358 363432 519414 363488
rect 519358 352960 519414 353016
rect 519266 346432 519322 346488
rect 519818 479032 519874 479088
rect 519818 437552 519874 437608
rect 519726 357312 519782 357368
rect 519634 344528 519690 344584
rect 520094 476176 520150 476232
rect 520094 476040 520150 476096
rect 520186 417832 520242 417888
rect 520186 414840 520242 414896
rect 520094 413616 520150 413672
rect 520002 412120 520058 412176
rect 520002 409128 520058 409184
rect 520186 406136 520242 406192
rect 520002 406000 520058 406056
rect 520002 396344 520058 396400
rect 520094 395528 520150 395584
rect 520002 393080 520058 393136
rect 520094 390632 520150 390688
rect 520462 377848 520518 377904
rect 520370 365200 520426 365256
rect 520278 358944 520334 359000
rect 519910 351056 519966 351112
rect 520830 403144 520886 403200
rect 521290 415792 521346 415848
rect 521658 459992 521714 460048
rect 521566 432520 521622 432576
rect 521474 424088 521530 424144
rect 521382 405184 521438 405240
rect 521198 379888 521254 379944
rect 521106 373632 521162 373688
rect 521014 367240 521070 367296
rect 520922 360984 520978 361040
rect 520738 354728 520794 354784
rect 520646 348336 520702 348392
rect 520554 342080 520610 342136
rect 316038 240644 316094 240680
rect 316038 240624 316040 240644
rect 316040 240624 316092 240644
rect 316092 240624 316094 240644
rect 325606 240660 325608 240680
rect 325608 240660 325660 240680
rect 325660 240660 325662 240680
rect 325606 240624 325662 240660
rect 357438 240644 357494 240680
rect 357438 240624 357440 240644
rect 357440 240624 357492 240644
rect 357492 240624 357494 240644
rect 360382 240644 360438 240680
rect 360382 240624 360384 240644
rect 360384 240624 360436 240644
rect 360436 240624 360438 240644
rect 288346 203904 288402 203960
rect 292486 204040 292542 204096
rect 289726 203768 289782 203824
rect 329378 212472 329434 212528
rect 330942 203632 330998 203688
rect 329746 203396 329748 203416
rect 329748 203396 329800 203416
rect 329800 203396 329802 203416
rect 329746 203360 329802 203396
rect 331126 203360 331182 203416
rect 328366 203224 328422 203280
rect 332506 203224 332562 203280
rect 335174 203360 335230 203416
rect 336646 220768 336702 220824
rect 336738 203360 336794 203416
rect 333886 203224 333942 203280
rect 335266 203224 335322 203280
rect 328274 203088 328330 203144
rect 332414 203088 332470 203144
rect 333794 203088 333850 203144
rect 336554 203088 336610 203144
rect 338210 203224 338266 203280
rect 340050 203496 340106 203552
rect 339590 203224 339646 203280
rect 340970 203632 341026 203688
rect 342258 203668 342260 203688
rect 342260 203668 342312 203688
rect 342312 203668 342314 203688
rect 342258 203632 342314 203668
rect 342258 203532 342260 203552
rect 342260 203532 342312 203552
rect 342312 203532 342314 203552
rect 342258 203496 342314 203532
rect 341706 203360 341762 203416
rect 335266 202952 335322 203008
rect 336646 202972 336702 203008
rect 336646 202952 336648 202972
rect 336648 202952 336700 202972
rect 336700 202952 336702 202972
rect 337934 202952 337990 203008
rect 339222 202952 339278 203008
rect 341338 202952 341394 203008
rect 343638 203496 343694 203552
rect 343638 203088 343694 203144
rect 347778 204176 347834 204232
rect 347778 203632 347834 203688
rect 349158 203632 349214 203688
rect 345570 203360 345626 203416
rect 346398 203224 346454 203280
rect 345018 203088 345074 203144
rect 349158 203260 349160 203280
rect 349160 203260 349212 203280
rect 349212 203260 349214 203280
rect 349158 203224 349214 203260
rect 351090 203124 351092 203144
rect 351092 203124 351144 203144
rect 351144 203124 351146 203144
rect 351090 203088 351146 203124
rect 355322 203904 355378 203960
rect 351918 203632 351974 203688
rect 354678 203496 354734 203552
rect 355322 203360 355378 203416
rect 357346 204176 357402 204232
rect 355966 203496 356022 203552
rect 357438 203904 357494 203960
rect 356058 203224 356114 203280
rect 357990 203088 358046 203144
rect 344926 202952 344982 203008
rect 345938 202952 345994 203008
rect 347042 202952 347098 203008
rect 348422 202952 348478 203008
rect 349434 202952 349490 203008
rect 351182 202952 351238 203008
rect 351642 202952 351698 203008
rect 353022 202952 353078 203008
rect 353298 202972 353354 203008
rect 353298 202952 353300 202972
rect 353300 202952 353352 202972
rect 353352 202952 353354 202972
rect 354586 202952 354642 203008
rect 355598 202952 355654 203008
rect 356426 202952 356482 203008
rect 362866 204176 362922 204232
rect 358726 203632 358782 203688
rect 360198 203496 360254 203552
rect 360198 203088 360254 203144
rect 364338 203360 364394 203416
rect 366822 203360 366878 203416
rect 366914 203224 366970 203280
rect 367098 204176 367154 204232
rect 368478 203260 368480 203280
rect 368480 203260 368532 203280
rect 368532 203260 368534 203280
rect 368478 203224 368534 203260
rect 371146 203224 371202 203280
rect 376574 203768 376630 203824
rect 376390 203632 376446 203688
rect 376574 203632 376630 203688
rect 375654 203224 375710 203280
rect 367006 203088 367062 203144
rect 373262 203088 373318 203144
rect 357438 202988 357440 203008
rect 357440 202988 357492 203008
rect 357492 202988 357494 203008
rect 357438 202952 357494 202988
rect 358634 202952 358690 203008
rect 358818 202952 358874 203008
rect 360014 202952 360070 203008
rect 361302 202952 361358 203008
rect 362866 202952 362922 203008
rect 363418 202952 363474 203008
rect 365074 202952 365130 203008
rect 375654 202952 375710 203008
rect 379794 182688 379850 182744
rect 297914 180240 297970 180296
rect 297914 171808 297970 171864
rect 297822 111696 297878 111752
rect 379978 123120 380034 123176
rect 380070 118088 380126 118144
rect 380530 180920 380586 180976
rect 380438 122032 380494 122088
rect 380346 120264 380402 120320
rect 380254 118632 380310 118688
rect 431774 231784 431830 231840
rect 431958 231784 432014 231840
rect 437478 203904 437534 203960
rect 442262 203768 442318 203824
rect 437478 203632 437534 203688
rect 448426 204176 448482 204232
rect 449806 204176 449862 204232
rect 449162 204076 449164 204096
rect 449164 204076 449216 204096
rect 449216 204076 449218 204096
rect 449162 204040 449218 204076
rect 450910 204040 450966 204096
rect 442262 203224 442318 203280
rect 451094 203904 451150 203960
rect 451094 203768 451150 203824
rect 451186 203632 451242 203688
rect 451094 203224 451150 203280
rect 451002 202952 451058 203008
rect 452566 204176 452622 204232
rect 453302 204176 453358 204232
rect 452014 204040 452070 204096
rect 455142 204176 455198 204232
rect 454682 204040 454738 204096
rect 453946 202988 453948 203008
rect 453948 202988 454000 203008
rect 454000 202988 454002 203008
rect 453946 202952 454002 202988
rect 456062 204040 456118 204096
rect 456706 204176 456762 204232
rect 456246 203360 456302 203416
rect 456706 203360 456762 203416
rect 457994 203904 458050 203960
rect 460846 203940 460848 203960
rect 460848 203940 460900 203960
rect 460900 203940 460902 203960
rect 460846 203904 460902 203940
rect 461582 203904 461638 203960
rect 459466 203224 459522 203280
rect 461582 203360 461638 203416
rect 462226 203224 462282 203280
rect 469126 204176 469182 204232
rect 464986 204040 465042 204096
rect 466274 204040 466330 204096
rect 470506 204176 470562 204232
rect 466366 203904 466422 203960
rect 470414 204040 470470 204096
rect 471242 203904 471298 203960
rect 463606 203360 463662 203416
rect 464710 203360 464766 203416
rect 463514 203224 463570 203280
rect 466366 203496 466422 203552
rect 467562 203380 467618 203416
rect 467562 203360 467564 203380
rect 467564 203360 467616 203380
rect 467616 203360 467618 203380
rect 469494 203360 469550 203416
rect 467746 203260 467748 203280
rect 467748 203260 467800 203280
rect 467800 203260 467802 203280
rect 467746 203224 467802 203260
rect 455326 202972 455382 203008
rect 455326 202952 455328 202972
rect 455328 202952 455380 202972
rect 455380 202952 455382 202972
rect 457902 202952 457958 203008
rect 459098 202952 459154 203008
rect 460662 202952 460718 203008
rect 461490 202952 461546 203008
rect 462410 202952 462466 203008
rect 463054 202952 463110 203008
rect 465906 202952 465962 203008
rect 467194 202952 467250 203008
rect 468482 202952 468538 203008
rect 470598 203224 470654 203280
rect 471242 203496 471298 203552
rect 471334 203224 471390 203280
rect 473910 203496 473966 203552
rect 474462 203496 474518 203552
rect 471886 203224 471942 203280
rect 472622 203224 472678 203280
rect 472898 203224 472954 203280
rect 473358 203224 473414 203280
rect 484398 204176 484454 204232
rect 475658 204040 475714 204096
rect 477498 204040 477554 204096
rect 483018 204076 483020 204096
rect 483020 204076 483072 204096
rect 483072 204076 483074 204096
rect 483018 204040 483074 204076
rect 485778 204040 485834 204096
rect 480166 203904 480222 203960
rect 474830 203224 474886 203280
rect 490194 203904 490250 203960
rect 480166 203496 480222 203552
rect 480626 203496 480682 203552
rect 477498 203360 477554 203416
rect 478878 203360 478934 203416
rect 477498 203244 477554 203280
rect 477498 203224 477500 203244
rect 477500 203224 477552 203244
rect 477552 203224 477554 203244
rect 478970 203224 479026 203280
rect 481638 203224 481694 203280
rect 484398 203532 484400 203552
rect 484400 203532 484452 203552
rect 484452 203532 484454 203552
rect 484398 203496 484454 203532
rect 471058 202952 471114 203008
rect 471794 202952 471850 203008
rect 475750 202952 475806 203008
rect 476118 202952 476174 203008
rect 477498 202952 477554 203008
rect 480534 202952 480590 203008
rect 481638 202952 481694 203008
rect 483018 202952 483074 203008
rect 448426 201320 448482 201376
rect 496450 181328 496506 181384
rect 417422 180512 417478 180568
rect 418066 171672 418122 171728
rect 380162 115776 380218 115832
rect 379978 114688 380034 114744
rect 300766 111288 300822 111344
rect 416778 111288 416834 111344
rect 303618 108996 303674 109032
rect 303618 108976 303620 108996
rect 303620 108976 303672 108996
rect 303672 108976 303674 108996
rect 307758 108996 307814 109032
rect 499762 118632 499818 118688
rect 500130 123664 500186 123720
rect 500038 122032 500094 122088
rect 499946 120808 500002 120864
rect 499854 118088 499910 118144
rect 521750 455776 521806 455832
rect 521842 453600 521898 453656
rect 521934 451560 521990 451616
rect 522026 449384 522082 449440
rect 522118 447344 522174 447400
rect 522210 443128 522266 443184
rect 522118 237088 522174 237144
rect 500314 183096 500370 183152
rect 500222 115776 500278 115832
rect 499670 115232 499726 115288
rect 307758 108976 307760 108996
rect 307760 108976 307812 108996
rect 307812 108976 307814 108996
rect 424230 108996 424286 109032
rect 424230 108976 424232 108996
rect 424232 108976 424284 108996
rect 424284 108976 424286 108996
rect 427818 108996 427874 109032
rect 427818 108976 427820 108996
rect 427820 108976 427872 108996
rect 427872 108976 427874 108996
rect 522394 440952 522450 441008
rect 522394 438912 522450 438968
rect 522302 400968 522358 401024
rect 522302 323040 522358 323096
rect 522302 316784 522358 316840
rect 522302 310428 522304 310448
rect 522304 310428 522356 310448
rect 522356 310428 522358 310448
rect 522302 310392 522358 310428
rect 522302 304136 522358 304192
rect 522302 278840 522358 278896
rect 522302 272584 522358 272640
rect 522302 249328 522358 249384
rect 522302 247288 522358 247344
rect 522302 245112 522358 245168
rect 522670 430480 522726 430536
rect 522946 445168 523002 445224
rect 522854 436736 522910 436792
rect 522946 426264 523002 426320
rect 523130 428304 523186 428360
rect 522762 422048 522818 422104
rect 522670 420044 522672 420064
rect 522672 420044 522724 420064
rect 522724 420044 522726 420064
rect 522670 420008 522726 420044
rect 522578 409400 522634 409456
rect 522486 407360 522542 407416
rect 522946 339904 523002 339960
rect 522946 337900 522948 337920
rect 522948 337900 523000 337920
rect 523000 337900 523002 337920
rect 522946 337864 523002 337900
rect 522578 335688 522634 335744
rect 522946 333648 523002 333704
rect 522578 331472 522634 331528
rect 522946 329432 523002 329488
rect 522946 327256 523002 327312
rect 522946 325216 523002 325272
rect 522670 321000 522726 321056
rect 522946 318824 523002 318880
rect 522946 314628 523002 314664
rect 522946 314608 522948 314628
rect 522948 314608 523000 314628
rect 523000 314608 523002 314628
rect 522946 312568 523002 312624
rect 522946 308352 523002 308408
rect 522946 306176 523002 306232
rect 522946 301960 523002 302016
rect 522946 299920 523002 299976
rect 522946 297880 523002 297936
rect 522946 295704 523002 295760
rect 522946 293664 523002 293720
rect 580170 697992 580226 698048
rect 542450 684392 542506 684448
rect 542542 678816 542598 678872
rect 542542 521600 542598 521656
rect 542726 521600 542782 521656
rect 542634 492768 542690 492824
rect 542542 492652 542598 492688
rect 542542 492632 542544 492652
rect 542544 492632 542596 492652
rect 542596 492632 542598 492652
rect 542358 454008 542414 454064
rect 542634 454008 542690 454064
rect 542174 434696 542230 434752
rect 542358 434696 542414 434752
rect 542174 415384 542230 415440
rect 542358 415384 542414 415440
rect 542082 394712 542138 394768
rect 542266 394712 542322 394768
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 580170 545536 580226 545592
rect 580170 533840 580226 533896
rect 580170 510312 580226 510368
rect 580170 498616 580226 498672
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 580170 451696 580226 451752
rect 580170 439864 580226 439920
rect 580170 416472 580226 416528
rect 580262 404776 580318 404832
rect 579894 392944 579950 393000
rect 579986 299104 580042 299160
rect 580354 369552 580410 369608
rect 522578 291488 522634 291544
rect 522946 289448 523002 289504
rect 580446 357856 580502 357912
rect 580538 346024 580594 346080
rect 522578 287272 522634 287328
rect 580630 322632 580686 322688
rect 522578 285232 522634 285288
rect 522486 283056 522542 283112
rect 580722 310800 580778 310856
rect 522946 281016 523002 281072
rect 522486 276800 522542 276856
rect 580170 275712 580226 275768
rect 522946 274624 523002 274680
rect 522854 270408 522910 270464
rect 522578 266192 522634 266248
rect 522762 264152 522818 264208
rect 522578 261976 522634 262032
rect 522578 259936 522634 259992
rect 522578 257760 522634 257816
rect 522486 251504 522542 251560
rect 522394 243072 522450 243128
rect 522394 240488 522450 240544
rect 522670 255720 522726 255776
rect 522946 268368 523002 268424
rect 523682 253544 523738 253600
rect 580170 263880 580226 263936
rect 579802 252184 579858 252240
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 579802 205264 579858 205320
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 89161 700770 89227 700773
rect 520590 700770 520596 700772
rect 89161 700768 520596 700770
rect 89161 700712 89166 700768
rect 89222 700712 520596 700768
rect 89161 700710 520596 700712
rect 89161 700707 89227 700710
rect 520590 700708 520596 700710
rect 520660 700708 520666 700772
rect 72969 700634 73035 700637
rect 518934 700634 518940 700636
rect 72969 700632 518940 700634
rect 72969 700576 72974 700632
rect 73030 700576 518940 700632
rect 72969 700574 518940 700576
rect 72969 700571 73035 700574
rect 518934 700572 518940 700574
rect 519004 700572 519010 700636
rect 24301 700498 24367 700501
rect 520774 700498 520780 700500
rect 24301 700496 520780 700498
rect 24301 700440 24306 700496
rect 24362 700440 520780 700496
rect 24301 700438 520780 700440
rect 24301 700435 24367 700438
rect 520774 700436 520780 700438
rect 520844 700436 520850 700500
rect 8109 700362 8175 700365
rect 514845 700362 514911 700365
rect 8109 700360 514911 700362
rect 8109 700304 8114 700360
rect 8170 700304 514850 700360
rect 514906 700304 514911 700360
rect 8109 700302 514911 700304
rect 8109 700299 8175 700302
rect 514845 700299 514911 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 514845 695738 514911 695741
rect 514845 695736 519554 695738
rect 514845 695680 514850 695736
rect 514906 695680 519554 695736
rect 514845 695678 519554 695680
rect 514845 695675 514911 695678
rect 519494 695604 519554 695678
rect 519486 695540 519492 695604
rect 519556 695540 519562 695604
rect 519486 695268 519492 695332
rect 519556 695330 519562 695332
rect 519629 695330 519695 695333
rect 519556 695328 519695 695330
rect 519556 695272 519634 695328
rect 519690 695272 519695 695328
rect 519556 695270 519695 695272
rect 519556 695268 519562 695270
rect 519629 695267 519695 695270
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 519629 686084 519695 686085
rect 519629 686082 519676 686084
rect 519584 686080 519676 686082
rect 519584 686024 519634 686080
rect 519584 686022 519676 686024
rect 519629 686020 519676 686022
rect 519740 686020 519746 686084
rect 519629 686019 519695 686020
rect 542445 684452 542511 684453
rect 519854 684388 519860 684452
rect 519924 684388 519930 684452
rect 542445 684448 542492 684452
rect 542556 684450 542562 684452
rect 542445 684392 542450 684448
rect 542445 684388 542492 684392
rect 542556 684390 542602 684450
rect 542556 684388 542562 684390
rect 519862 684317 519922 684388
rect 542445 684387 542511 684388
rect 519862 684312 519971 684317
rect 519862 684256 519910 684312
rect 519966 684256 519971 684312
rect 519862 684254 519971 684256
rect 519905 684251 519971 684254
rect -960 682274 480 682364
rect -960 682214 674 682274
rect -960 682124 480 682214
rect 614 681866 674 682214
rect 519302 681866 519308 681868
rect 614 681806 519308 681866
rect 519302 681804 519308 681806
rect 519372 681804 519378 681868
rect 542537 678876 542603 678877
rect 542486 678874 542492 678876
rect 542446 678814 542492 678874
rect 542556 678872 542603 678876
rect 542598 678816 542603 678872
rect 542486 678812 542492 678814
rect 542556 678812 542603 678816
rect 542537 678811 542603 678812
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 520958 667994 520964 667996
rect -960 667934 520964 667994
rect -960 667844 480 667934
rect 520958 667932 520964 667934
rect 521028 667932 521034 667996
rect 519905 666634 519971 666637
rect 520038 666634 520044 666636
rect 519905 666632 520044 666634
rect 519905 666576 519910 666632
rect 519966 666576 520044 666632
rect 519905 666574 520044 666576
rect 519905 666571 519971 666574
rect 520038 666572 520044 666574
rect 520108 666572 520114 666636
rect 583520 662676 584960 662916
rect 519486 659636 519492 659700
rect 519556 659698 519562 659700
rect 520038 659698 520044 659700
rect 519556 659638 520044 659698
rect 519556 659636 519562 659638
rect 520038 659636 520044 659638
rect 520108 659636 520114 659700
rect -960 653578 480 653668
rect 3325 653578 3391 653581
rect -960 653576 3391 653578
rect -960 653520 3330 653576
rect 3386 653520 3391 653576
rect -960 653518 3391 653520
rect -960 653428 480 653518
rect 3325 653515 3391 653518
rect 3325 652898 3391 652901
rect 519486 652898 519492 652900
rect 3325 652896 519492 652898
rect 3325 652840 3330 652896
rect 3386 652840 519492 652896
rect 3325 652838 519492 652840
rect 3325 652835 3391 652838
rect 519486 652836 519492 652838
rect 519556 652836 519562 652900
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 519118 644540 519124 644604
rect 519188 644602 519194 644604
rect 519854 644602 519860 644604
rect 519188 644542 519860 644602
rect 519188 644540 519194 644542
rect 519854 644540 519860 644542
rect 519924 644540 519930 644604
rect 519118 644404 519124 644468
rect 519188 644466 519194 644468
rect 519670 644466 519676 644468
rect 519188 644406 519676 644466
rect 519188 644404 519194 644406
rect 519670 644404 519676 644406
rect 519740 644404 519746 644468
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 519118 634884 519124 634948
rect 519188 634946 519194 634948
rect 519670 634946 519676 634948
rect 519188 634886 519676 634946
rect 519188 634884 519194 634886
rect 519670 634884 519676 634886
rect 519740 634884 519746 634948
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect 519118 625092 519124 625156
rect 519188 625154 519194 625156
rect 519854 625154 519860 625156
rect 519188 625094 519860 625154
rect 519188 625092 519194 625094
rect 519854 625092 519860 625094
rect 519924 625092 519930 625156
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 3417 623794 3483 623797
rect 519670 623794 519676 623796
rect 3417 623792 519676 623794
rect 3417 623736 3422 623792
rect 3478 623736 519676 623792
rect 3417 623734 519676 623736
rect 3417 623731 3483 623734
rect 519670 623732 519676 623734
rect 519740 623732 519746 623796
rect 583520 615756 584960 615996
rect 519118 615572 519124 615636
rect 519188 615634 519194 615636
rect 519854 615634 519860 615636
rect 519188 615574 519860 615634
rect 519188 615572 519194 615574
rect 519854 615572 519860 615574
rect 519924 615572 519930 615636
rect 373625 612780 373691 612781
rect 373574 612716 373580 612780
rect 373644 612778 373691 612780
rect 488533 612780 488599 612781
rect 493961 612780 494027 612781
rect 373644 612776 373736 612778
rect 373686 612720 373736 612776
rect 373644 612718 373736 612720
rect 488533 612776 488580 612780
rect 488644 612778 488650 612780
rect 493910 612778 493916 612780
rect 488533 612720 488538 612776
rect 373644 612716 373691 612718
rect 373625 612715 373691 612716
rect 488533 612716 488580 612720
rect 488644 612718 488690 612778
rect 493870 612718 493916 612778
rect 493980 612776 494027 612780
rect 494022 612720 494027 612776
rect 488644 612716 488650 612718
rect 493910 612716 493916 612718
rect 493980 612716 494027 612720
rect 488533 612715 488599 612716
rect 493961 612715 494027 612716
rect 369158 610948 369164 611012
rect 369228 611010 369234 611012
rect 373022 611010 373028 611012
rect 369228 610950 373028 611010
rect 369228 610948 369234 610950
rect 373022 610948 373028 610950
rect 373092 610948 373098 611012
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 496445 609922 496511 609925
rect 496445 609920 496554 609922
rect 496445 609864 496450 609920
rect 496506 609864 496554 609920
rect 496445 609859 496554 609864
rect 377292 609653 377874 609713
rect 496494 609683 496554 609859
rect 377814 609650 377874 609653
rect 379697 609650 379763 609653
rect 379973 609650 380039 609653
rect 377814 609648 380039 609650
rect 377814 609592 379702 609648
rect 379758 609592 379978 609648
rect 380034 609592 380039 609648
rect 377814 609590 380039 609592
rect 379697 609587 379763 609590
rect 379973 609587 380039 609590
rect 298001 606658 298067 606661
rect 298001 606656 299490 606658
rect 298001 606600 298006 606656
rect 298062 606617 299490 606656
rect 298062 606600 300012 606617
rect 298001 606598 300012 606600
rect 298001 606595 298067 606598
rect 299430 606557 300012 606598
rect 416773 606114 416839 606117
rect 420134 606114 420194 606587
rect 416773 606112 420194 606114
rect 416773 606056 416778 606112
rect 416834 606056 420194 606112
rect 416773 606054 420194 606056
rect 416773 606051 416839 606054
rect 519118 605780 519124 605844
rect 519188 605842 519194 605844
rect 519854 605842 519860 605844
rect 519188 605782 519860 605842
rect 519188 605780 519194 605782
rect 519854 605780 519860 605782
rect 519924 605780 519930 605844
rect 297909 605434 297975 605437
rect 299430 605434 300012 605489
rect 297909 605432 300012 605434
rect 297909 605376 297914 605432
rect 297970 605429 300012 605432
rect 297970 605376 299490 605429
rect 297909 605374 299490 605376
rect 297909 605371 297975 605374
rect 416773 604890 416839 604893
rect 420134 604890 420194 605459
rect 416773 604888 420194 604890
rect 416773 604832 416778 604888
rect 416834 604832 420194 604888
rect 416773 604830 420194 604832
rect 416773 604827 416839 604830
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect 297817 603802 297883 603805
rect 297817 603800 299490 603802
rect 297817 603744 297822 603800
rect 297878 603789 299490 603800
rect 297878 603744 300012 603789
rect 297817 603742 300012 603744
rect 297817 603739 297883 603742
rect 299430 603729 300012 603742
rect 416773 603258 416839 603261
rect 420134 603258 420194 603759
rect 416773 603256 420194 603258
rect 416773 603200 416778 603256
rect 416834 603200 420194 603256
rect 416773 603198 420194 603200
rect 416773 603195 416839 603198
rect 299430 602601 300012 602661
rect 297725 602578 297791 602581
rect 299430 602578 299490 602601
rect 297725 602576 299490 602578
rect 297725 602520 297730 602576
rect 297786 602520 299490 602576
rect 297725 602518 299490 602520
rect 297725 602515 297791 602518
rect 416773 602034 416839 602037
rect 420134 602034 420194 602631
rect 416773 602032 420194 602034
rect 416773 601976 416778 602032
rect 416834 601976 420194 602032
rect 416773 601974 420194 601976
rect 416773 601971 416839 601974
rect 297633 600946 297699 600949
rect 299430 600946 300012 600961
rect 297633 600944 300012 600946
rect 297633 600888 297638 600944
rect 297694 600901 300012 600944
rect 297694 600888 299490 600901
rect 297633 600886 299490 600888
rect 297633 600883 297699 600886
rect 416773 600538 416839 600541
rect 420134 600538 420194 600931
rect 416773 600536 420194 600538
rect 416773 600480 416778 600536
rect 416834 600480 420194 600536
rect 416773 600478 420194 600480
rect 416773 600475 416839 600478
rect 297541 599858 297607 599861
rect 297541 599856 299490 599858
rect 297541 599800 297546 599856
rect 297602 599833 299490 599856
rect 297602 599800 300012 599833
rect 297541 599798 300012 599800
rect 297541 599795 297607 599798
rect 299430 599773 300012 599798
rect 416773 599314 416839 599317
rect 420134 599314 420194 599803
rect 416773 599312 420194 599314
rect 416773 599256 416778 599312
rect 416834 599256 420194 599312
rect 416773 599254 420194 599256
rect 416773 599251 416839 599254
rect 297449 598090 297515 598093
rect 299430 598090 300012 598133
rect 297449 598088 300012 598090
rect 297449 598032 297454 598088
rect 297510 598073 300012 598088
rect 297510 598032 299490 598073
rect 297449 598030 299490 598032
rect 297449 598027 297515 598030
rect 416773 597682 416839 597685
rect 420134 597682 420194 598103
rect 416773 597680 420194 597682
rect 416773 597624 416778 597680
rect 416834 597624 420194 597680
rect 416773 597622 420194 597624
rect 416773 597619 416839 597622
rect 519118 596260 519124 596324
rect 519188 596322 519194 596324
rect 519854 596322 519860 596324
rect 519188 596262 519860 596322
rect 519188 596260 519194 596262
rect 519854 596260 519860 596262
rect 519924 596260 519930 596324
rect -960 596050 480 596140
rect 3509 596050 3575 596053
rect -960 596048 3575 596050
rect -960 595992 3514 596048
rect 3570 595992 3575 596048
rect -960 595990 3575 595992
rect -960 595900 480 595990
rect 3509 595987 3575 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect 519118 586332 519124 586396
rect 519188 586394 519194 586396
rect 519854 586394 519860 586396
rect 519188 586334 519860 586394
rect 519188 586332 519194 586334
rect 519854 586332 519860 586334
rect 519924 586332 519930 586396
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 519118 576812 519124 576876
rect 519188 576874 519194 576876
rect 519854 576874 519860 576876
rect 519188 576814 519860 576874
rect 519188 576812 519194 576814
rect 519854 576812 519860 576814
rect 519924 576812 519930 576876
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3601 567354 3667 567357
rect -960 567352 3667 567354
rect -960 567296 3606 567352
rect 3662 567296 3667 567352
rect -960 567294 3667 567296
rect -960 567204 480 567294
rect 3601 567291 3667 567294
rect 519118 567020 519124 567084
rect 519188 567082 519194 567084
rect 519854 567082 519860 567084
rect 519188 567022 519860 567082
rect 519188 567020 519194 567022
rect 519854 567020 519860 567022
rect 519924 567020 519930 567084
rect 519118 557500 519124 557564
rect 519188 557562 519194 557564
rect 519854 557562 519860 557564
rect 519188 557502 519860 557562
rect 519188 557500 519194 557502
rect 519854 557500 519860 557502
rect 519924 557500 519930 557564
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3693 553074 3759 553077
rect -960 553072 3759 553074
rect -960 553016 3698 553072
rect 3754 553016 3759 553072
rect -960 553014 3759 553016
rect -960 552924 480 553014
rect 3693 553011 3759 553014
rect 499573 549538 499639 549541
rect 497782 549536 499639 549538
rect 497782 549480 499578 549536
rect 499634 549480 499639 549536
rect 497782 549478 499639 549480
rect 497782 549442 497842 549478
rect 499573 549475 499639 549478
rect 377108 549412 377874 549442
rect 497076 549412 497842 549442
rect 377078 549402 377874 549412
rect 379605 549402 379671 549405
rect 377078 549400 379671 549402
rect 377078 549382 379610 549400
rect 377078 540958 377138 549382
rect 377814 549344 379610 549382
rect 379666 549344 379671 549400
rect 377814 549342 379671 549344
rect 379605 549339 379671 549342
rect 497046 549382 497842 549412
rect 497046 547906 497106 549382
rect 497046 547846 497290 547906
rect 497230 542058 497290 547846
rect 519118 547708 519124 547772
rect 519188 547770 519194 547772
rect 519854 547770 519860 547772
rect 519188 547710 519860 547770
rect 519188 547708 519194 547710
rect 519854 547708 519860 547710
rect 519924 547708 519930 547772
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 499573 542058 499639 542061
rect 497230 542056 499639 542058
rect 497230 542000 499578 542056
rect 499634 542000 499639 542056
rect 497230 541998 499639 542000
rect 499573 541995 499639 541998
rect 379789 540970 379855 540973
rect 499573 540970 499639 540973
rect 377446 540968 379855 540970
rect 377446 540958 379794 540968
rect 377078 540928 379794 540958
rect 377108 540912 379794 540928
rect 379850 540912 379855 540968
rect 377108 540910 379855 540912
rect 497230 540968 499639 540970
rect 497230 540912 499578 540968
rect 499634 540912 499639 540968
rect 497230 540910 499639 540912
rect 377108 540898 377506 540910
rect 379789 540907 379855 540910
rect 499573 540907 499639 540910
rect 297357 540290 297423 540293
rect 297357 540288 299490 540290
rect 297357 540232 297362 540288
rect 297418 540285 299490 540288
rect 297418 540232 300012 540285
rect 297357 540230 300012 540232
rect 297357 540227 297423 540230
rect 299430 540225 300012 540230
rect 416773 539746 416839 539749
rect 420134 539746 420194 540255
rect 416773 539744 420194 539746
rect 416773 539688 416778 539744
rect 416834 539688 420194 539744
rect 416773 539686 420194 539688
rect 416773 539683 416839 539686
rect -960 538658 480 538748
rect 3785 538658 3851 538661
rect -960 538656 3851 538658
rect -960 538600 3790 538656
rect 3846 538600 3851 538656
rect -960 538598 3851 538600
rect -960 538508 480 538598
rect 3785 538595 3851 538598
rect 299430 538525 300012 538585
rect 297265 538522 297331 538525
rect 299430 538522 299490 538525
rect 297265 538520 299490 538522
rect 297265 538464 297270 538520
rect 297326 538464 299490 538520
rect 297265 538462 299490 538464
rect 297265 538459 297331 538462
rect 416773 538386 416839 538389
rect 420134 538386 420194 538555
rect 416773 538384 420194 538386
rect 416773 538328 416778 538384
rect 416834 538328 420194 538384
rect 416773 538326 420194 538328
rect 416773 538323 416839 538326
rect 519118 538188 519124 538252
rect 519188 538250 519194 538252
rect 519854 538250 519860 538252
rect 519188 538190 519860 538250
rect 519188 538188 519194 538190
rect 519854 538188 519860 538190
rect 519924 538188 519930 538252
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 519118 528396 519124 528460
rect 519188 528458 519194 528460
rect 519854 528458 519860 528460
rect 519188 528398 519860 528458
rect 519188 528396 519194 528398
rect 519854 528396 519860 528398
rect 519924 528396 519930 528460
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 542537 521658 542603 521661
rect 542721 521658 542787 521661
rect 542537 521656 542787 521658
rect 542537 521600 542542 521656
rect 542598 521600 542726 521656
rect 542782 521600 542787 521656
rect 542537 521598 542787 521600
rect 542537 521595 542603 521598
rect 542721 521595 542787 521598
rect 425605 519754 425671 519757
rect 427962 519754 427968 519756
rect 425605 519752 427968 519754
rect 425605 519696 425610 519752
rect 425666 519696 427968 519752
rect 425605 519694 427968 519696
rect 425605 519691 425671 519694
rect 427962 519692 427968 519694
rect 428032 519692 428038 519756
rect 519118 518876 519124 518940
rect 519188 518938 519194 518940
rect 519854 518938 519860 518940
rect 519188 518878 519860 518938
rect 519188 518876 519194 518878
rect 519854 518876 519860 518878
rect 519924 518876 519930 518940
rect 313774 518740 313780 518804
rect 313844 518802 313850 518804
rect 314561 518802 314627 518805
rect 313844 518800 314627 518802
rect 313844 518744 314566 518800
rect 314622 518744 314627 518800
rect 313844 518742 314627 518744
rect 313844 518740 313850 518742
rect 314561 518739 314627 518742
rect 316166 518740 316172 518804
rect 316236 518802 316242 518804
rect 317321 518802 317387 518805
rect 316236 518800 317387 518802
rect 316236 518744 317326 518800
rect 317382 518744 317387 518800
rect 316236 518742 317387 518744
rect 316236 518740 316242 518742
rect 317321 518739 317387 518742
rect 318558 518740 318564 518804
rect 318628 518802 318634 518804
rect 318701 518802 318767 518805
rect 321737 518804 321803 518805
rect 321686 518802 321692 518804
rect 318628 518800 318767 518802
rect 318628 518744 318706 518800
rect 318762 518744 318767 518800
rect 318628 518742 318767 518744
rect 321646 518742 321692 518802
rect 321756 518800 321803 518804
rect 321798 518744 321803 518800
rect 318628 518740 318634 518742
rect 318701 518739 318767 518742
rect 321686 518740 321692 518742
rect 321756 518740 321803 518744
rect 321737 518739 321803 518740
rect 323117 518804 323183 518805
rect 323117 518800 323164 518804
rect 323228 518802 323234 518804
rect 324313 518802 324379 518805
rect 324446 518802 324452 518804
rect 323117 518744 323122 518800
rect 323117 518740 323164 518744
rect 323228 518742 323274 518802
rect 324313 518800 324452 518802
rect 324313 518744 324318 518800
rect 324374 518744 324452 518800
rect 324313 518742 324452 518744
rect 323228 518740 323234 518742
rect 323117 518739 323183 518740
rect 324313 518739 324379 518742
rect 324446 518740 324452 518742
rect 324516 518740 324522 518804
rect 325182 518740 325188 518804
rect 325252 518802 325258 518804
rect 325417 518802 325483 518805
rect 325252 518800 325483 518802
rect 325252 518744 325422 518800
rect 325478 518744 325483 518800
rect 325252 518742 325483 518744
rect 325252 518740 325258 518742
rect 325417 518739 325483 518742
rect 326429 518804 326495 518805
rect 327165 518804 327231 518805
rect 328913 518804 328979 518805
rect 326429 518800 326476 518804
rect 326540 518802 326546 518804
rect 326429 518744 326434 518800
rect 326429 518740 326476 518744
rect 326540 518742 326586 518802
rect 327165 518800 327212 518804
rect 327276 518802 327282 518804
rect 328862 518802 328868 518804
rect 327165 518744 327170 518800
rect 326540 518740 326546 518742
rect 327165 518740 327212 518744
rect 327276 518742 327322 518802
rect 328822 518742 328868 518802
rect 328932 518800 328979 518804
rect 328974 518744 328979 518800
rect 327276 518740 327282 518742
rect 328862 518740 328868 518742
rect 328932 518740 328979 518744
rect 326429 518739 326495 518740
rect 327165 518739 327231 518740
rect 328913 518739 328979 518740
rect 330109 518804 330175 518805
rect 332317 518804 332383 518805
rect 335537 518804 335603 518805
rect 330109 518800 330156 518804
rect 330220 518802 330226 518804
rect 330109 518744 330114 518800
rect 330109 518740 330156 518744
rect 330220 518742 330266 518802
rect 332317 518800 332364 518804
rect 332428 518802 332434 518804
rect 335486 518802 335492 518804
rect 332317 518744 332322 518800
rect 330220 518740 330226 518742
rect 332317 518740 332364 518744
rect 332428 518742 332474 518802
rect 335446 518742 335492 518802
rect 335556 518800 335603 518804
rect 335598 518744 335603 518800
rect 332428 518740 332434 518742
rect 335486 518740 335492 518742
rect 335556 518740 335603 518744
rect 330109 518739 330175 518740
rect 332317 518739 332383 518740
rect 335537 518739 335603 518740
rect 336733 518802 336799 518805
rect 337193 518804 337259 518805
rect 337142 518802 337148 518804
rect 336733 518800 337148 518802
rect 337212 518800 337259 518804
rect 336733 518744 336738 518800
rect 336794 518744 337148 518800
rect 337254 518744 337259 518800
rect 336733 518742 337148 518744
rect 336733 518739 336799 518742
rect 337142 518740 337148 518742
rect 337212 518740 337259 518744
rect 339350 518740 339356 518804
rect 339420 518802 339426 518804
rect 339953 518802 340019 518805
rect 340505 518804 340571 518805
rect 341609 518804 341675 518805
rect 340454 518802 340460 518804
rect 339420 518800 340019 518802
rect 339420 518744 339958 518800
rect 340014 518744 340019 518800
rect 339420 518742 340019 518744
rect 340414 518742 340460 518802
rect 340524 518800 340571 518804
rect 341558 518802 341564 518804
rect 340566 518744 340571 518800
rect 339420 518740 339426 518742
rect 337193 518739 337259 518740
rect 339953 518739 340019 518742
rect 340454 518740 340460 518742
rect 340524 518740 340571 518744
rect 341518 518742 341564 518802
rect 341628 518800 341675 518804
rect 341670 518744 341675 518800
rect 341558 518740 341564 518742
rect 341628 518740 341675 518744
rect 340505 518739 340571 518740
rect 341609 518739 341675 518740
rect 342989 518804 343055 518805
rect 344185 518804 344251 518805
rect 345473 518804 345539 518805
rect 342989 518800 343036 518804
rect 343100 518802 343106 518804
rect 344134 518802 344140 518804
rect 342989 518744 342994 518800
rect 342989 518740 343036 518744
rect 343100 518742 343146 518802
rect 344094 518742 344140 518802
rect 344204 518800 344251 518804
rect 345422 518802 345428 518804
rect 344246 518744 344251 518800
rect 343100 518740 343106 518742
rect 344134 518740 344140 518742
rect 344204 518740 344251 518744
rect 345382 518742 345428 518802
rect 345492 518800 345539 518804
rect 345534 518744 345539 518800
rect 345422 518740 345428 518742
rect 345492 518740 345539 518744
rect 342989 518739 343055 518740
rect 344185 518739 344251 518740
rect 345473 518739 345539 518740
rect 346485 518804 346551 518805
rect 347681 518804 347747 518805
rect 348601 518804 348667 518805
rect 443177 518804 443243 518805
rect 451273 518804 451339 518805
rect 452561 518804 452627 518805
rect 453665 518804 453731 518805
rect 346485 518800 346532 518804
rect 346596 518802 346602 518804
rect 347630 518802 347636 518804
rect 346485 518744 346490 518800
rect 346485 518740 346532 518744
rect 346596 518742 346642 518802
rect 347590 518742 347636 518802
rect 347700 518800 347747 518804
rect 348550 518802 348556 518804
rect 347742 518744 347747 518800
rect 346596 518740 346602 518742
rect 347630 518740 347636 518742
rect 347700 518740 347747 518744
rect 348510 518742 348556 518802
rect 348620 518800 348667 518804
rect 443126 518802 443132 518804
rect 348662 518744 348667 518800
rect 348550 518740 348556 518742
rect 348620 518740 348667 518744
rect 443086 518742 443132 518802
rect 443196 518800 443243 518804
rect 443238 518744 443243 518800
rect 443126 518740 443132 518742
rect 443196 518740 443243 518744
rect 451222 518740 451228 518804
rect 451292 518802 451339 518804
rect 452510 518802 452516 518804
rect 451292 518800 451384 518802
rect 451334 518744 451384 518800
rect 451292 518742 451384 518744
rect 452470 518742 452516 518802
rect 452580 518800 452627 518804
rect 453614 518802 453620 518804
rect 452622 518744 452627 518800
rect 451292 518740 451339 518742
rect 452510 518740 452516 518742
rect 452580 518740 452627 518744
rect 453574 518742 453620 518802
rect 453684 518800 453731 518804
rect 453726 518744 453731 518800
rect 453614 518740 453620 518742
rect 453684 518740 453731 518744
rect 346485 518739 346551 518740
rect 347681 518739 347747 518740
rect 348601 518739 348667 518740
rect 443177 518739 443243 518740
rect 451273 518739 451339 518740
rect 452561 518739 452627 518740
rect 453665 518739 453731 518740
rect 459553 518802 459619 518805
rect 460422 518802 460428 518804
rect 459553 518800 460428 518802
rect 459553 518744 459558 518800
rect 459614 518744 460428 518800
rect 459553 518742 460428 518744
rect 459553 518739 459619 518742
rect 460422 518740 460428 518742
rect 460492 518740 460498 518804
rect 460933 518802 460999 518805
rect 461158 518802 461164 518804
rect 460933 518800 461164 518802
rect 460933 518744 460938 518800
rect 460994 518744 461164 518800
rect 460933 518742 461164 518744
rect 460933 518739 460999 518742
rect 461158 518740 461164 518742
rect 461228 518740 461234 518804
rect 462313 518802 462379 518805
rect 462446 518802 462452 518804
rect 462313 518800 462452 518802
rect 462313 518744 462318 518800
rect 462374 518744 462452 518800
rect 462313 518742 462452 518744
rect 462313 518739 462379 518742
rect 462446 518740 462452 518742
rect 462516 518740 462522 518804
rect 314694 518604 314700 518668
rect 314764 518666 314770 518668
rect 315941 518666 316007 518669
rect 317321 518668 317387 518669
rect 314764 518664 316007 518666
rect 314764 518608 315946 518664
rect 316002 518608 316007 518664
rect 314764 518606 316007 518608
rect 314764 518604 314770 518606
rect 315941 518603 316007 518606
rect 317270 518604 317276 518668
rect 317340 518666 317387 518668
rect 317340 518664 317432 518666
rect 317382 518608 317432 518664
rect 317340 518606 317432 518608
rect 317340 518604 317387 518606
rect 319662 518604 319668 518668
rect 319732 518666 319738 518668
rect 320081 518666 320147 518669
rect 319732 518664 320147 518666
rect 319732 518608 320086 518664
rect 320142 518608 320147 518664
rect 319732 518606 320147 518608
rect 319732 518604 319738 518606
rect 317321 518603 317387 518604
rect 320081 518603 320147 518606
rect 324262 518604 324268 518668
rect 324332 518666 324338 518668
rect 324405 518666 324471 518669
rect 324332 518664 324471 518666
rect 324332 518608 324410 518664
rect 324466 518608 324471 518664
rect 324332 518606 324471 518608
rect 324332 518604 324338 518606
rect 324405 518603 324471 518606
rect 331213 518668 331279 518669
rect 338113 518668 338179 518669
rect 331213 518664 331260 518668
rect 331324 518666 331330 518668
rect 338062 518666 338068 518668
rect 331213 518608 331218 518664
rect 331213 518604 331260 518608
rect 331324 518606 331370 518666
rect 338022 518606 338068 518666
rect 338132 518664 338179 518668
rect 338174 518608 338179 518664
rect 331324 518604 331330 518606
rect 338062 518604 338068 518606
rect 338132 518604 338179 518608
rect 331213 518603 331279 518604
rect 338113 518603 338179 518604
rect 429285 518666 429351 518669
rect 429694 518666 429700 518668
rect 429285 518664 429700 518666
rect 429285 518608 429290 518664
rect 429346 518608 429700 518664
rect 429285 518606 429700 518608
rect 429285 518603 429351 518606
rect 429694 518604 429700 518606
rect 429764 518604 429770 518668
rect 454718 518604 454724 518668
rect 454788 518666 454794 518668
rect 455321 518666 455387 518669
rect 456057 518668 456123 518669
rect 456006 518666 456012 518668
rect 454788 518664 455387 518666
rect 454788 518608 455326 518664
rect 455382 518608 455387 518664
rect 454788 518606 455387 518608
rect 455966 518606 456012 518666
rect 456076 518664 456123 518668
rect 456118 518608 456123 518664
rect 454788 518604 454794 518606
rect 455321 518603 455387 518606
rect 456006 518604 456012 518606
rect 456076 518604 456123 518608
rect 456057 518603 456123 518604
rect 456885 518666 456951 518669
rect 457110 518666 457116 518668
rect 456885 518664 457116 518666
rect 456885 518608 456890 518664
rect 456946 518608 457116 518664
rect 456885 518606 457116 518608
rect 456885 518603 456951 518606
rect 457110 518604 457116 518606
rect 457180 518604 457186 518668
rect 458265 518666 458331 518669
rect 459553 518668 459619 518669
rect 458398 518666 458404 518668
rect 458265 518664 458404 518666
rect 458265 518608 458270 518664
rect 458326 518608 458404 518664
rect 458265 518606 458404 518608
rect 458265 518603 458331 518606
rect 458398 518604 458404 518606
rect 458468 518604 458474 518668
rect 459502 518666 459508 518668
rect 459462 518606 459508 518666
rect 459572 518664 459619 518668
rect 459614 518608 459619 518664
rect 459502 518604 459508 518606
rect 459572 518604 459619 518608
rect 459553 518603 459619 518604
rect 465073 518666 465139 518669
rect 465206 518666 465212 518668
rect 465073 518664 465212 518666
rect 465073 518608 465078 518664
rect 465134 518608 465212 518664
rect 465073 518606 465212 518608
rect 465073 518603 465139 518606
rect 465206 518604 465212 518606
rect 465276 518604 465282 518668
rect 466545 518666 466611 518669
rect 467414 518666 467420 518668
rect 466545 518664 467420 518666
rect 466545 518608 466550 518664
rect 466606 518608 467420 518664
rect 466545 518606 467420 518608
rect 466545 518603 466611 518606
rect 467414 518604 467420 518606
rect 467484 518604 467490 518668
rect 316033 518530 316099 518533
rect 316534 518530 316540 518532
rect 316033 518528 316540 518530
rect 316033 518472 316038 518528
rect 316094 518472 316540 518528
rect 316033 518470 316540 518472
rect 316033 518467 316099 518470
rect 316534 518468 316540 518470
rect 316604 518468 316610 518532
rect 317505 518530 317571 518533
rect 318558 518530 318564 518532
rect 317505 518528 318564 518530
rect 317505 518472 317510 518528
rect 317566 518472 318564 518528
rect 317505 518470 318564 518472
rect 317505 518467 317571 518470
rect 318558 518468 318564 518470
rect 318628 518468 318634 518532
rect 327073 518530 327139 518533
rect 333421 518532 333487 518533
rect 334157 518532 334223 518533
rect 327942 518530 327948 518532
rect 327073 518528 327948 518530
rect 327073 518472 327078 518528
rect 327134 518472 327948 518528
rect 327073 518470 327948 518472
rect 327073 518467 327139 518470
rect 327942 518468 327948 518470
rect 328012 518468 328018 518532
rect 333421 518528 333468 518532
rect 333532 518530 333538 518532
rect 333421 518472 333426 518528
rect 333421 518468 333468 518472
rect 333532 518470 333578 518530
rect 334157 518528 334204 518532
rect 334268 518530 334274 518532
rect 426433 518530 426499 518533
rect 445385 518532 445451 518533
rect 426566 518530 426572 518532
rect 334157 518472 334162 518528
rect 333532 518468 333538 518470
rect 334157 518468 334204 518472
rect 334268 518470 334314 518530
rect 426433 518528 426572 518530
rect 426433 518472 426438 518528
rect 426494 518472 426572 518528
rect 426433 518470 426572 518472
rect 334268 518468 334274 518470
rect 333421 518467 333487 518468
rect 334157 518467 334223 518468
rect 426433 518467 426499 518470
rect 426566 518468 426572 518470
rect 426636 518468 426642 518532
rect 445334 518530 445340 518532
rect 445294 518470 445340 518530
rect 445404 518528 445451 518532
rect 445446 518472 445451 518528
rect 445334 518468 445340 518470
rect 445404 518468 445451 518472
rect 445385 518467 445451 518468
rect 446581 518532 446647 518533
rect 446581 518528 446628 518532
rect 446692 518530 446698 518532
rect 447409 518530 447475 518533
rect 466453 518532 466519 518533
rect 447726 518530 447732 518532
rect 446581 518472 446586 518528
rect 446581 518468 446628 518472
rect 446692 518470 446738 518530
rect 447409 518528 447732 518530
rect 447409 518472 447414 518528
rect 447470 518472 447732 518528
rect 447409 518470 447732 518472
rect 446692 518468 446698 518470
rect 446581 518467 446647 518468
rect 447409 518467 447475 518470
rect 447726 518468 447732 518470
rect 447796 518468 447802 518532
rect 466453 518530 466500 518532
rect 466408 518528 466500 518530
rect 466408 518472 466458 518528
rect 466408 518470 466500 518472
rect 466453 518468 466500 518470
rect 466564 518468 466570 518532
rect 466453 518467 466519 518468
rect 312486 518332 312492 518396
rect 312556 518394 312562 518396
rect 313181 518394 313247 518397
rect 317413 518396 317479 518397
rect 317413 518394 317460 518396
rect 312556 518392 313247 518394
rect 312556 518336 313186 518392
rect 313242 518336 313247 518392
rect 312556 518334 313247 518336
rect 317368 518392 317460 518394
rect 317368 518336 317418 518392
rect 317368 518334 317460 518336
rect 312556 518332 312562 518334
rect 313181 518331 313247 518334
rect 317413 518332 317460 518334
rect 317524 518332 317530 518396
rect 320766 518332 320772 518396
rect 320836 518394 320842 518396
rect 321093 518394 321159 518397
rect 320836 518392 321159 518394
rect 320836 518336 321098 518392
rect 321154 518336 321159 518392
rect 320836 518334 321159 518336
rect 320836 518332 320842 518334
rect 317413 518331 317479 518332
rect 321093 518331 321159 518334
rect 430573 518394 430639 518397
rect 442073 518396 442139 518397
rect 430798 518394 430804 518396
rect 430573 518392 430804 518394
rect 430573 518336 430578 518392
rect 430634 518336 430804 518392
rect 430573 518334 430804 518336
rect 430573 518331 430639 518334
rect 430798 518332 430804 518334
rect 430868 518332 430874 518396
rect 442022 518394 442028 518396
rect 441982 518334 442028 518394
rect 442092 518392 442139 518396
rect 442134 518336 442139 518392
rect 442022 518332 442028 518334
rect 442092 518332 442139 518336
rect 444046 518332 444052 518396
rect 444116 518394 444122 518396
rect 444281 518394 444347 518397
rect 444116 518392 444347 518394
rect 444116 518336 444286 518392
rect 444342 518336 444347 518392
rect 444116 518334 444347 518336
rect 444116 518332 444122 518334
rect 442073 518331 442139 518332
rect 444281 518331 444347 518334
rect 448789 518396 448855 518397
rect 449893 518396 449959 518397
rect 448789 518392 448836 518396
rect 448900 518394 448906 518396
rect 448789 518336 448794 518392
rect 448789 518332 448836 518336
rect 448900 518334 448946 518394
rect 449893 518392 449940 518396
rect 450004 518394 450010 518396
rect 463693 518394 463759 518397
rect 463918 518394 463924 518396
rect 449893 518336 449898 518392
rect 448900 518332 448906 518334
rect 449893 518332 449940 518336
rect 450004 518334 450050 518394
rect 463693 518392 463924 518394
rect 463693 518336 463698 518392
rect 463754 518336 463924 518392
rect 463693 518334 463924 518336
rect 450004 518332 450010 518334
rect 448789 518331 448855 518332
rect 449893 518331 449959 518332
rect 463693 518331 463759 518334
rect 463918 518332 463924 518334
rect 463988 518332 463994 518396
rect 467833 518394 467899 518397
rect 468518 518394 468524 518396
rect 467833 518392 468524 518394
rect 467833 518336 467838 518392
rect 467894 518336 468524 518392
rect 467833 518334 468524 518336
rect 467833 518331 467899 518334
rect 468518 518332 468524 518334
rect 468588 518332 468594 518396
rect 303613 518260 303679 518261
rect 303613 518256 303660 518260
rect 303724 518258 303730 518260
rect 314653 518258 314719 518261
rect 315062 518258 315068 518260
rect 303613 518200 303618 518256
rect 303613 518196 303660 518200
rect 303724 518198 303770 518258
rect 314653 518256 315068 518258
rect 314653 518200 314658 518256
rect 314714 518200 315068 518256
rect 314653 518198 315068 518200
rect 303724 518196 303730 518198
rect 303613 518195 303679 518196
rect 314653 518195 314719 518198
rect 315062 518196 315068 518198
rect 315132 518196 315138 518260
rect 322933 518258 322999 518261
rect 323526 518258 323532 518260
rect 322933 518256 323532 518258
rect 322933 518200 322938 518256
rect 322994 518200 323532 518256
rect 322933 518198 323532 518200
rect 322933 518195 322999 518198
rect 323526 518196 323532 518198
rect 323596 518196 323602 518260
rect 423673 518258 423739 518261
rect 429193 518260 429259 518261
rect 423806 518258 423812 518260
rect 423673 518256 423812 518258
rect 423673 518200 423678 518256
rect 423734 518200 423812 518256
rect 423673 518198 423812 518200
rect 423673 518195 423739 518198
rect 423806 518196 423812 518198
rect 423876 518196 423882 518260
rect 429142 518196 429148 518260
rect 429212 518258 429259 518260
rect 429212 518256 429304 518258
rect 429254 518200 429304 518256
rect 429212 518198 429304 518200
rect 429212 518196 429259 518198
rect 429193 518195 429259 518196
rect 318793 518122 318859 518125
rect 320030 518122 320036 518124
rect 318793 518120 320036 518122
rect 318793 518064 318798 518120
rect 318854 518064 320036 518120
rect 318793 518062 320036 518064
rect 318793 518059 318859 518062
rect 320030 518060 320036 518062
rect 320100 518060 320106 518124
rect 321829 518122 321895 518125
rect 322054 518122 322060 518124
rect 321829 518120 322060 518122
rect 321829 518064 321834 518120
rect 321890 518064 322060 518120
rect 321829 518062 322060 518064
rect 321829 518059 321895 518062
rect 322054 518060 322060 518062
rect 322124 518060 322130 518124
rect 435030 518060 435036 518124
rect 435100 518122 435106 518124
rect 435357 518122 435423 518125
rect 435909 518122 435975 518125
rect 435100 518120 435975 518122
rect 435100 518064 435362 518120
rect 435418 518064 435914 518120
rect 435970 518064 435975 518120
rect 435100 518062 435975 518064
rect 435100 518060 435106 518062
rect 435357 518059 435423 518062
rect 435909 518059 435975 518062
rect 312077 517986 312143 517989
rect 312670 517986 312676 517988
rect 312077 517984 312676 517986
rect 312077 517928 312082 517984
rect 312138 517928 312676 517984
rect 312077 517926 312676 517928
rect 312077 517923 312143 517926
rect 312670 517924 312676 517926
rect 312740 517924 312746 517988
rect 331213 517986 331279 517989
rect 331438 517986 331444 517988
rect 331213 517984 331444 517986
rect 331213 517928 331218 517984
rect 331274 517928 331444 517984
rect 331213 517926 331444 517928
rect 331213 517923 331279 517926
rect 331438 517924 331444 517926
rect 331508 517924 331514 517988
rect 332593 517986 332659 517989
rect 437289 517988 437355 517989
rect 332726 517986 332732 517988
rect 332593 517984 332732 517986
rect 332593 517928 332598 517984
rect 332654 517928 332732 517984
rect 332593 517926 332732 517928
rect 332593 517923 332659 517926
rect 332726 517924 332732 517926
rect 332796 517924 332802 517988
rect 437238 517924 437244 517988
rect 437308 517986 437355 517988
rect 437308 517984 437400 517986
rect 437350 517928 437400 517984
rect 437308 517926 437400 517928
rect 437308 517924 437355 517926
rect 437289 517923 437355 517924
rect 320173 517850 320239 517853
rect 320950 517850 320956 517852
rect 320173 517848 320956 517850
rect 320173 517792 320178 517848
rect 320234 517792 320956 517848
rect 320173 517790 320956 517792
rect 320173 517787 320239 517790
rect 320950 517788 320956 517790
rect 321020 517788 321026 517852
rect 333973 517850 334039 517853
rect 432597 517852 432663 517853
rect 334934 517850 334940 517852
rect 333973 517848 334940 517850
rect 333973 517792 333978 517848
rect 334034 517792 334940 517848
rect 333973 517790 334940 517792
rect 333973 517787 334039 517790
rect 334934 517788 334940 517790
rect 335004 517788 335010 517852
rect 432597 517850 432644 517852
rect 432552 517848 432644 517850
rect 432552 517792 432602 517848
rect 432552 517790 432644 517792
rect 432597 517788 432644 517790
rect 432708 517788 432714 517852
rect 433742 517788 433748 517852
rect 433812 517850 433818 517852
rect 433885 517850 433951 517853
rect 433812 517848 433951 517850
rect 433812 517792 433890 517848
rect 433946 517792 433951 517848
rect 433812 517790 433951 517792
rect 433812 517788 433818 517790
rect 432597 517787 432663 517788
rect 433885 517787 433951 517790
rect 440734 517788 440740 517852
rect 440804 517850 440810 517852
rect 440877 517850 440943 517853
rect 440804 517848 440943 517850
rect 440804 517792 440882 517848
rect 440938 517792 440943 517848
rect 440804 517790 440943 517792
rect 440804 517788 440810 517790
rect 440877 517787 440943 517790
rect 309726 517652 309732 517716
rect 309796 517714 309802 517716
rect 310329 517714 310395 517717
rect 309796 517712 310395 517714
rect 309796 517656 310334 517712
rect 310390 517656 310395 517712
rect 309796 517654 310395 517656
rect 309796 517652 309802 517654
rect 310329 517651 310395 517654
rect 313273 517714 313339 517717
rect 313958 517714 313964 517716
rect 313273 517712 313964 517714
rect 313273 517656 313278 517712
rect 313334 517656 313964 517712
rect 313273 517654 313964 517656
rect 313273 517651 313339 517654
rect 313958 517652 313964 517654
rect 314028 517652 314034 517716
rect 324313 517714 324379 517717
rect 325550 517714 325556 517716
rect 324313 517712 325556 517714
rect 324313 517656 324318 517712
rect 324374 517656 325556 517712
rect 324313 517654 325556 517656
rect 324313 517651 324379 517654
rect 325550 517652 325556 517654
rect 325620 517652 325626 517716
rect 329833 517714 329899 517717
rect 330334 517714 330340 517716
rect 329833 517712 330340 517714
rect 329833 517656 329838 517712
rect 329894 517656 330340 517712
rect 329833 517654 330340 517656
rect 329833 517651 329899 517654
rect 330334 517652 330340 517654
rect 330404 517652 330410 517716
rect 332593 517714 332659 517717
rect 333830 517714 333836 517716
rect 332593 517712 333836 517714
rect 332593 517656 332598 517712
rect 332654 517656 333836 517712
rect 332593 517654 333836 517656
rect 332593 517651 332659 517654
rect 333830 517652 333836 517654
rect 333900 517652 333906 517716
rect 335721 517714 335787 517717
rect 336038 517714 336044 517716
rect 335721 517712 336044 517714
rect 335721 517656 335726 517712
rect 335782 517656 336044 517712
rect 335721 517654 336044 517656
rect 335721 517651 335787 517654
rect 336038 517652 336044 517654
rect 336108 517652 336114 517716
rect 338113 517714 338179 517717
rect 339493 517716 339559 517717
rect 338430 517714 338436 517716
rect 338113 517712 338436 517714
rect 338113 517656 338118 517712
rect 338174 517656 338436 517712
rect 338113 517654 338436 517656
rect 338113 517651 338179 517654
rect 338430 517652 338436 517654
rect 338500 517652 338506 517716
rect 339493 517714 339540 517716
rect 339448 517712 339540 517714
rect 339448 517656 339498 517712
rect 339448 517654 339540 517656
rect 339493 517652 339540 517654
rect 339604 517652 339610 517716
rect 342897 517714 342963 517717
rect 344277 517716 344343 517717
rect 343398 517714 343404 517716
rect 342897 517712 343404 517714
rect 342897 517656 342902 517712
rect 342958 517656 343404 517712
rect 342897 517654 343404 517656
rect 339493 517651 339559 517652
rect 342897 517651 342963 517654
rect 343398 517652 343404 517654
rect 343468 517652 343474 517716
rect 344277 517714 344324 517716
rect 344232 517712 344324 517714
rect 344232 517656 344282 517712
rect 344232 517654 344324 517656
rect 344277 517652 344324 517654
rect 344388 517652 344394 517716
rect 345790 517652 345796 517716
rect 345860 517714 345866 517716
rect 346301 517714 346367 517717
rect 345860 517712 346367 517714
rect 345860 517656 346306 517712
rect 346362 517656 346367 517712
rect 345860 517654 346367 517656
rect 345860 517652 345866 517654
rect 344277 517651 344343 517652
rect 346301 517651 346367 517654
rect 347262 517652 347268 517716
rect 347332 517714 347338 517716
rect 348417 517714 348483 517717
rect 348969 517716 349035 517717
rect 347332 517712 348483 517714
rect 347332 517656 348422 517712
rect 348478 517656 348483 517712
rect 347332 517654 348483 517656
rect 347332 517652 347338 517654
rect 348417 517651 348483 517654
rect 348918 517652 348924 517716
rect 348988 517714 349035 517716
rect 348988 517712 349080 517714
rect 349030 517656 349080 517712
rect 348988 517654 349080 517656
rect 348988 517652 349035 517654
rect 433006 517652 433012 517716
rect 433076 517714 433082 517716
rect 433241 517714 433307 517717
rect 433076 517712 433307 517714
rect 433076 517656 433246 517712
rect 433302 517656 433307 517712
rect 433076 517654 433307 517656
rect 433076 517652 433082 517654
rect 348969 517651 349035 517652
rect 433241 517651 433307 517654
rect 433926 517652 433932 517716
rect 433996 517714 434002 517716
rect 434621 517714 434687 517717
rect 433996 517712 434687 517714
rect 433996 517656 434626 517712
rect 434682 517656 434687 517712
rect 433996 517654 434687 517656
rect 433996 517652 434002 517654
rect 434621 517651 434687 517654
rect 435766 517652 435772 517716
rect 435836 517714 435842 517716
rect 436001 517714 436067 517717
rect 435836 517712 436067 517714
rect 435836 517656 436006 517712
rect 436062 517656 436067 517712
rect 435836 517654 436067 517656
rect 435836 517652 435842 517654
rect 436001 517651 436067 517654
rect 436134 517652 436140 517716
rect 436204 517714 436210 517716
rect 436645 517714 436711 517717
rect 436204 517712 436711 517714
rect 436204 517656 436650 517712
rect 436706 517656 436711 517712
rect 436204 517654 436711 517656
rect 436204 517652 436210 517654
rect 436645 517651 436711 517654
rect 436870 517652 436876 517716
rect 436940 517714 436946 517716
rect 437381 517714 437447 517717
rect 436940 517712 437447 517714
rect 436940 517656 437386 517712
rect 437442 517656 437447 517712
rect 436940 517654 437447 517656
rect 436940 517652 436946 517654
rect 437381 517651 437447 517654
rect 437974 517652 437980 517716
rect 438044 517714 438050 517716
rect 438669 517714 438735 517717
rect 438044 517712 438735 517714
rect 438044 517656 438674 517712
rect 438730 517656 438735 517712
rect 438044 517654 438735 517656
rect 438044 517652 438050 517654
rect 438669 517651 438735 517654
rect 439497 517714 439563 517717
rect 439630 517714 439636 517716
rect 439497 517712 439636 517714
rect 439497 517656 439502 517712
rect 439558 517656 439636 517712
rect 439497 517654 439636 517656
rect 439497 517651 439563 517654
rect 439630 517652 439636 517654
rect 439700 517652 439706 517716
rect 444966 517652 444972 517716
rect 445036 517714 445042 517716
rect 445661 517714 445727 517717
rect 445036 517712 445727 517714
rect 445036 517656 445666 517712
rect 445722 517656 445727 517712
rect 445036 517654 445727 517656
rect 445036 517652 445042 517654
rect 445661 517651 445727 517654
rect 453246 517652 453252 517716
rect 453316 517714 453322 517716
rect 453941 517714 454007 517717
rect 453316 517712 454007 517714
rect 453316 517656 453946 517712
rect 454002 517656 454007 517712
rect 453316 517654 454007 517656
rect 453316 517652 453322 517654
rect 453941 517651 454007 517654
rect 460238 517652 460244 517716
rect 460308 517714 460314 517716
rect 460841 517714 460907 517717
rect 460308 517712 460907 517714
rect 460308 517656 460846 517712
rect 460902 517656 460907 517712
rect 460308 517654 460907 517656
rect 460308 517652 460314 517654
rect 460841 517651 460907 517654
rect 468334 517652 468340 517716
rect 468404 517714 468410 517716
rect 469121 517714 469187 517717
rect 468404 517712 469187 517714
rect 468404 517656 469126 517712
rect 469182 517656 469187 517712
rect 468404 517654 469187 517656
rect 468404 517652 468410 517654
rect 469121 517651 469187 517654
rect 307334 517516 307340 517580
rect 307404 517578 307410 517580
rect 307661 517578 307727 517581
rect 307404 517576 307727 517578
rect 307404 517520 307666 517576
rect 307722 517520 307727 517576
rect 307404 517518 307727 517520
rect 307404 517516 307410 517518
rect 307661 517515 307727 517518
rect 308622 517516 308628 517580
rect 308692 517578 308698 517580
rect 309041 517578 309107 517581
rect 310237 517580 310303 517581
rect 310237 517578 310284 517580
rect 308692 517576 309107 517578
rect 308692 517520 309046 517576
rect 309102 517520 309107 517576
rect 308692 517518 309107 517520
rect 310192 517576 310284 517578
rect 310192 517520 310242 517576
rect 310192 517518 310284 517520
rect 308692 517516 308698 517518
rect 309041 517515 309107 517518
rect 310237 517516 310284 517518
rect 310348 517516 310354 517580
rect 311566 517516 311572 517580
rect 311636 517578 311642 517580
rect 311709 517578 311775 517581
rect 311636 517576 311775 517578
rect 311636 517520 311714 517576
rect 311770 517520 311775 517576
rect 311636 517518 311775 517520
rect 311636 517516 311642 517518
rect 310237 517515 310303 517516
rect 311709 517515 311775 517518
rect 325693 517578 325759 517581
rect 326654 517578 326660 517580
rect 325693 517576 326660 517578
rect 325693 517520 325698 517576
rect 325754 517520 326660 517576
rect 325693 517518 326660 517520
rect 325693 517515 325759 517518
rect 326654 517516 326660 517518
rect 326724 517516 326730 517580
rect 328453 517578 328519 517581
rect 329046 517578 329052 517580
rect 328453 517576 329052 517578
rect 328453 517520 328458 517576
rect 328514 517520 329052 517576
rect 328453 517518 329052 517520
rect 328453 517515 328519 517518
rect 329046 517516 329052 517518
rect 329116 517516 329122 517580
rect 336733 517578 336799 517581
rect 337326 517578 337332 517580
rect 336733 517576 337332 517578
rect 336733 517520 336738 517576
rect 336794 517520 337332 517576
rect 336733 517518 337332 517520
rect 336733 517515 336799 517518
rect 337326 517516 337332 517518
rect 337396 517516 337402 517580
rect 339401 517578 339467 517581
rect 340638 517578 340644 517580
rect 339401 517576 340644 517578
rect 339401 517520 339406 517576
rect 339462 517520 340644 517576
rect 339401 517518 340644 517520
rect 339401 517515 339467 517518
rect 340638 517516 340644 517518
rect 340708 517516 340714 517580
rect 340781 517578 340847 517581
rect 341926 517578 341932 517580
rect 340781 517576 341932 517578
rect 340781 517520 340786 517576
rect 340842 517520 341932 517576
rect 340781 517518 341932 517520
rect 340781 517515 340847 517518
rect 341926 517516 341932 517518
rect 341996 517516 342002 517580
rect 348366 517516 348372 517580
rect 348436 517578 348442 517580
rect 349061 517578 349127 517581
rect 348436 517576 349127 517578
rect 348436 517520 349066 517576
rect 349122 517520 349127 517576
rect 348436 517518 349127 517520
rect 348436 517516 348442 517518
rect 349061 517515 349127 517518
rect 438117 517578 438183 517581
rect 438761 517580 438827 517581
rect 438342 517578 438348 517580
rect 438117 517576 438348 517578
rect 438117 517520 438122 517576
rect 438178 517520 438348 517576
rect 438117 517518 438348 517520
rect 438117 517515 438183 517518
rect 438342 517516 438348 517518
rect 438412 517516 438418 517580
rect 438710 517578 438716 517580
rect 438670 517518 438716 517578
rect 438780 517576 438827 517580
rect 438822 517520 438827 517576
rect 438710 517516 438716 517518
rect 438780 517516 438827 517520
rect 439998 517516 440004 517580
rect 440068 517578 440074 517580
rect 440141 517578 440207 517581
rect 441521 517580 441587 517581
rect 441470 517578 441476 517580
rect 440068 517576 440207 517578
rect 440068 517520 440146 517576
rect 440202 517520 440207 517576
rect 440068 517518 440207 517520
rect 441430 517518 441476 517578
rect 441540 517576 441587 517580
rect 441582 517520 441587 517576
rect 440068 517516 440074 517518
rect 438761 517515 438827 517516
rect 440141 517515 440207 517518
rect 441470 517516 441476 517518
rect 441540 517516 441587 517520
rect 442758 517516 442764 517580
rect 442828 517578 442834 517580
rect 442901 517578 442967 517581
rect 442828 517576 442967 517578
rect 442828 517520 442906 517576
rect 442962 517520 442967 517576
rect 442828 517518 442967 517520
rect 442828 517516 442834 517518
rect 441521 517515 441587 517516
rect 442901 517515 442967 517518
rect 443862 517516 443868 517580
rect 443932 517578 443938 517580
rect 444281 517578 444347 517581
rect 445569 517580 445635 517581
rect 447041 517580 447107 517581
rect 445518 517578 445524 517580
rect 443932 517576 444347 517578
rect 443932 517520 444286 517576
rect 444342 517520 444347 517576
rect 443932 517518 444347 517520
rect 445478 517518 445524 517578
rect 445588 517576 445635 517580
rect 446990 517578 446996 517580
rect 445630 517520 445635 517576
rect 443932 517516 443938 517518
rect 444281 517515 444347 517518
rect 445518 517516 445524 517518
rect 445588 517516 445635 517520
rect 446950 517518 446996 517578
rect 447060 517576 447107 517580
rect 447102 517520 447107 517576
rect 446990 517516 446996 517518
rect 447060 517516 447107 517520
rect 448278 517516 448284 517580
rect 448348 517578 448354 517580
rect 448421 517578 448487 517581
rect 449801 517580 449867 517581
rect 449750 517578 449756 517580
rect 448348 517576 448487 517578
rect 448348 517520 448426 517576
rect 448482 517520 448487 517576
rect 448348 517518 448487 517520
rect 449710 517518 449756 517578
rect 449820 517576 449867 517580
rect 449862 517520 449867 517576
rect 448348 517516 448354 517518
rect 445569 517515 445635 517516
rect 447041 517515 447107 517516
rect 448421 517515 448487 517518
rect 449750 517516 449756 517518
rect 449820 517516 449867 517520
rect 450854 517516 450860 517580
rect 450924 517578 450930 517580
rect 451181 517578 451247 517581
rect 450924 517576 451247 517578
rect 450924 517520 451186 517576
rect 451242 517520 451247 517576
rect 450924 517518 451247 517520
rect 450924 517516 450930 517518
rect 449801 517515 449867 517516
rect 451181 517515 451247 517518
rect 451958 517516 451964 517580
rect 452028 517578 452034 517580
rect 452561 517578 452627 517581
rect 453849 517580 453915 517581
rect 455321 517580 455387 517581
rect 453798 517578 453804 517580
rect 452028 517576 452627 517578
rect 452028 517520 452566 517576
rect 452622 517520 452627 517576
rect 452028 517518 452627 517520
rect 453758 517518 453804 517578
rect 453868 517576 453915 517580
rect 455270 517578 455276 517580
rect 453910 517520 453915 517576
rect 452028 517516 452034 517518
rect 452561 517515 452627 517518
rect 453798 517516 453804 517518
rect 453868 517516 453915 517520
rect 455230 517518 455276 517578
rect 455340 517576 455387 517580
rect 455382 517520 455387 517576
rect 455270 517516 455276 517518
rect 455340 517516 455387 517520
rect 456374 517516 456380 517580
rect 456444 517578 456450 517580
rect 456701 517578 456767 517581
rect 456444 517576 456767 517578
rect 456444 517520 456706 517576
rect 456762 517520 456767 517576
rect 456444 517518 456767 517520
rect 456444 517516 456450 517518
rect 453849 517515 453915 517516
rect 455321 517515 455387 517516
rect 456701 517515 456767 517518
rect 457846 517516 457852 517580
rect 457916 517578 457922 517580
rect 458081 517578 458147 517581
rect 457916 517576 458147 517578
rect 457916 517520 458086 517576
rect 458142 517520 458147 517576
rect 457916 517518 458147 517520
rect 457916 517516 457922 517518
rect 458081 517515 458147 517518
rect 459134 517516 459140 517580
rect 459204 517578 459210 517580
rect 459461 517578 459527 517581
rect 460749 517580 460815 517581
rect 460749 517578 460796 517580
rect 459204 517576 459527 517578
rect 459204 517520 459466 517576
rect 459522 517520 459527 517576
rect 459204 517518 459527 517520
rect 460704 517576 460796 517578
rect 460704 517520 460754 517576
rect 460704 517518 460796 517520
rect 459204 517516 459210 517518
rect 459461 517515 459527 517518
rect 460749 517516 460796 517518
rect 460860 517516 460866 517580
rect 462078 517516 462084 517580
rect 462148 517578 462154 517580
rect 462221 517578 462287 517581
rect 463601 517580 463667 517581
rect 463550 517578 463556 517580
rect 462148 517576 462287 517578
rect 462148 517520 462226 517576
rect 462282 517520 462287 517576
rect 462148 517518 462287 517520
rect 463510 517518 463556 517578
rect 463620 517576 463667 517580
rect 463662 517520 463667 517576
rect 462148 517516 462154 517518
rect 460749 517515 460815 517516
rect 462221 517515 462287 517518
rect 463550 517516 463556 517518
rect 463620 517516 463667 517520
rect 464838 517516 464844 517580
rect 464908 517578 464914 517580
rect 464981 517578 465047 517581
rect 464908 517576 465047 517578
rect 464908 517520 464986 517576
rect 465042 517520 465047 517576
rect 464908 517518 465047 517520
rect 464908 517516 464914 517518
rect 463601 517515 463667 517516
rect 464981 517515 465047 517518
rect 466126 517516 466132 517580
rect 466196 517578 466202 517580
rect 466361 517578 466427 517581
rect 466196 517576 466427 517578
rect 466196 517520 466366 517576
rect 466422 517520 466427 517576
rect 466196 517518 466427 517520
rect 466196 517516 466202 517518
rect 466361 517515 466427 517518
rect 467230 517516 467236 517580
rect 467300 517578 467306 517580
rect 467741 517578 467807 517581
rect 469029 517580 469095 517581
rect 469029 517578 469076 517580
rect 467300 517576 467807 517578
rect 467300 517520 467746 517576
rect 467802 517520 467807 517576
rect 467300 517518 467807 517520
rect 468984 517576 469076 517578
rect 468984 517520 469034 517576
rect 468984 517518 469076 517520
rect 467300 517516 467306 517518
rect 467741 517515 467807 517518
rect 469029 517516 469076 517518
rect 469140 517516 469146 517580
rect 469029 517515 469095 517516
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3325 509962 3391 509965
rect -960 509960 3391 509962
rect -960 509904 3330 509960
rect 3386 509904 3391 509960
rect -960 509902 3391 509904
rect -960 509812 480 509902
rect 3325 509899 3391 509902
rect 519118 509084 519124 509148
rect 519188 509146 519194 509148
rect 519854 509146 519860 509148
rect 519188 509086 519860 509146
rect 519188 509084 519194 509086
rect 519854 509084 519860 509086
rect 519924 509084 519930 509148
rect 519118 499564 519124 499628
rect 519188 499626 519194 499628
rect 519854 499626 519860 499628
rect 519188 499566 519860 499626
rect 519188 499564 519194 499566
rect 519854 499564 519860 499566
rect 519924 499564 519930 499628
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3417 495546 3483 495549
rect -960 495544 3483 495546
rect -960 495488 3422 495544
rect 3478 495488 3483 495544
rect -960 495486 3483 495488
rect -960 495396 480 495486
rect 3417 495483 3483 495486
rect 542629 492826 542695 492829
rect 542494 492824 542695 492826
rect 542494 492768 542634 492824
rect 542690 492768 542695 492824
rect 542494 492766 542695 492768
rect 542494 492693 542554 492766
rect 542629 492763 542695 492766
rect 542494 492688 542603 492693
rect 542494 492632 542542 492688
rect 542598 492632 542603 492688
rect 542494 492630 542603 492632
rect 542537 492627 542603 492630
rect 519118 489772 519124 489836
rect 519188 489834 519194 489836
rect 519854 489834 519860 489836
rect 519188 489774 519860 489834
rect 519188 489772 519194 489774
rect 519854 489772 519860 489774
rect 519924 489772 519930 489836
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 433609 483034 433675 483037
rect 433793 483034 433859 483037
rect 433609 483032 433859 483034
rect 433609 482976 433614 483032
rect 433670 482976 433798 483032
rect 433854 482976 433859 483032
rect 433609 482974 433859 482976
rect 433609 482971 433675 482974
rect 433793 482971 433859 482974
rect 463601 482490 463667 482493
rect 507485 482490 507551 482493
rect 463601 482488 507551 482490
rect 463601 482432 463606 482488
rect 463662 482432 507490 482488
rect 507546 482432 507551 482488
rect 463601 482430 507551 482432
rect 463601 482427 463667 482430
rect 507485 482427 507551 482430
rect 467741 482354 467807 482357
rect 514109 482354 514175 482357
rect 467741 482352 514175 482354
rect 467741 482296 467746 482352
rect 467802 482296 514114 482352
rect 514170 482296 514175 482352
rect 467741 482294 514175 482296
rect 467741 482291 467807 482294
rect 514109 482291 514175 482294
rect 469029 482218 469095 482221
rect 518525 482218 518591 482221
rect 469029 482216 518591 482218
rect 469029 482160 469034 482216
rect 469090 482160 518530 482216
rect 518586 482160 518591 482216
rect 469029 482158 518591 482160
rect 469029 482155 469095 482158
rect 518525 482155 518591 482158
rect -960 481130 480 481220
rect 2957 481130 3023 481133
rect -960 481128 3023 481130
rect -960 481072 2962 481128
rect 3018 481072 3023 481128
rect -960 481070 3023 481072
rect -960 480980 480 481070
rect 2957 481067 3023 481070
rect 357382 479980 357388 480044
rect 357452 480042 357458 480044
rect 362217 480042 362283 480045
rect 357452 480040 362283 480042
rect 357452 479984 362222 480040
rect 362278 479984 362283 480040
rect 357452 479982 362283 479984
rect 357452 479980 357458 479982
rect 362217 479979 362283 479982
rect 369945 480042 370011 480045
rect 376702 480042 376708 480044
rect 369945 480040 376708 480042
rect 369945 479984 369950 480040
rect 370006 479984 376708 480040
rect 369945 479982 376708 479984
rect 369945 479979 370011 479982
rect 376702 479980 376708 479982
rect 376772 479980 376778 480044
rect 67582 479844 67588 479908
rect 67652 479906 67658 479908
rect 71313 479906 71379 479909
rect 67652 479904 71379 479906
rect 67652 479848 71318 479904
rect 71374 479848 71379 479904
rect 67652 479846 71379 479848
rect 67652 479844 67658 479846
rect 71313 479843 71379 479846
rect 362217 479770 362283 479773
rect 367093 479770 367159 479773
rect 362217 479768 367159 479770
rect 362217 479712 362222 479768
rect 362278 479712 367098 479768
rect 367154 479712 367159 479768
rect 362217 479710 367159 479712
rect 362217 479707 362283 479710
rect 367093 479707 367159 479710
rect 434662 479708 434668 479772
rect 434732 479770 434738 479772
rect 444281 479770 444347 479773
rect 434732 479768 444347 479770
rect 434732 479712 444286 479768
rect 444342 479712 444347 479768
rect 434732 479710 444347 479712
rect 434732 479708 434738 479710
rect 444281 479707 444347 479710
rect 446998 479710 463802 479770
rect 61837 479634 61903 479637
rect 67582 479634 67588 479636
rect 61837 479632 67588 479634
rect 61837 479576 61842 479632
rect 61898 479576 67588 479632
rect 61837 479574 67588 479576
rect 61837 479571 61903 479574
rect 67582 479572 67588 479574
rect 67652 479572 67658 479636
rect 71313 479634 71379 479637
rect 71313 479632 77218 479634
rect 71313 479576 71318 479632
rect 71374 479576 77218 479632
rect 71313 479574 77218 479576
rect 71313 479571 71379 479574
rect 50981 479498 51047 479501
rect 41462 479496 51047 479498
rect 41462 479440 50986 479496
rect 51042 479440 51047 479496
rect 41462 479438 51047 479440
rect 77158 479498 77218 479574
rect 96662 479540 96906 479600
rect 106222 479572 106228 479636
rect 106292 479634 106298 479636
rect 108941 479634 109007 479637
rect 106292 479632 109007 479634
rect 106292 479576 108946 479632
rect 109002 479576 109007 479632
rect 106292 479574 109007 479576
rect 106292 479572 106298 479574
rect 108941 479571 109007 479574
rect 109125 479634 109191 479637
rect 316769 479634 316835 479637
rect 318742 479634 318748 479636
rect 109125 479632 118802 479634
rect 109125 479576 109130 479632
rect 109186 479576 118802 479632
rect 109125 479574 118802 479576
rect 109125 479571 109191 479574
rect 77158 479438 77402 479498
rect 41321 479362 41387 479365
rect 41462 479362 41522 479438
rect 50981 479435 51047 479438
rect 41321 479360 41522 479362
rect 41321 479304 41326 479360
rect 41382 479304 41522 479360
rect 41321 479302 41522 479304
rect 57789 479362 57855 479365
rect 57973 479362 58039 479365
rect 77342 479364 77402 479438
rect 77518 479436 77524 479500
rect 77588 479498 77594 479500
rect 86902 479498 86908 479500
rect 77588 479438 86908 479498
rect 77588 479436 77594 479438
rect 86902 479436 86908 479438
rect 86972 479436 86978 479500
rect 96470 479436 96476 479500
rect 96540 479498 96546 479500
rect 96662 479498 96722 479540
rect 96540 479438 96722 479498
rect 96846 479498 96906 479540
rect 99373 479498 99439 479501
rect 96846 479496 99439 479498
rect 96846 479440 99378 479496
rect 99434 479440 99439 479496
rect 96846 479438 99439 479440
rect 96540 479436 96546 479438
rect 99373 479435 99439 479438
rect 57789 479360 58039 479362
rect 57789 479304 57794 479360
rect 57850 479304 57978 479360
rect 58034 479304 58039 479360
rect 57789 479302 58039 479304
rect 41321 479299 41387 479302
rect 57789 479299 57855 479302
rect 57973 479299 58039 479302
rect 77334 479300 77340 479364
rect 77404 479300 77410 479364
rect 118742 479362 118802 479574
rect 292438 479574 302434 479634
rect 135161 479498 135227 479501
rect 154481 479498 154547 479501
rect 173801 479498 173867 479501
rect 193121 479498 193187 479501
rect 212441 479498 212507 479501
rect 231761 479498 231827 479501
rect 251081 479498 251147 479501
rect 278773 479498 278839 479501
rect 135161 479496 138122 479498
rect 135161 479440 135166 479496
rect 135222 479440 138122 479496
rect 135161 479438 138122 479440
rect 135161 479435 135227 479438
rect 128261 479362 128327 479365
rect 118742 479360 128327 479362
rect 118742 479304 128266 479360
rect 128322 479304 128327 479360
rect 118742 479302 128327 479304
rect 138062 479362 138122 479438
rect 154481 479496 157442 479498
rect 154481 479440 154486 479496
rect 154542 479440 157442 479496
rect 154481 479438 157442 479440
rect 154481 479435 154547 479438
rect 147581 479362 147647 479365
rect 138062 479360 147647 479362
rect 138062 479304 147586 479360
rect 147642 479304 147647 479360
rect 138062 479302 147647 479304
rect 157382 479362 157442 479438
rect 173801 479496 176762 479498
rect 173801 479440 173806 479496
rect 173862 479440 176762 479496
rect 173801 479438 176762 479440
rect 173801 479435 173867 479438
rect 166901 479362 166967 479365
rect 157382 479360 166967 479362
rect 157382 479304 166906 479360
rect 166962 479304 166967 479360
rect 157382 479302 166967 479304
rect 176702 479362 176762 479438
rect 193121 479496 196082 479498
rect 193121 479440 193126 479496
rect 193182 479440 196082 479496
rect 193121 479438 196082 479440
rect 193121 479435 193187 479438
rect 186221 479362 186287 479365
rect 176702 479360 186287 479362
rect 176702 479304 186226 479360
rect 186282 479304 186287 479360
rect 176702 479302 186287 479304
rect 196022 479362 196082 479438
rect 212441 479496 215402 479498
rect 212441 479440 212446 479496
rect 212502 479440 215402 479496
rect 212441 479438 215402 479440
rect 212441 479435 212507 479438
rect 205541 479362 205607 479365
rect 196022 479360 205607 479362
rect 196022 479304 205546 479360
rect 205602 479304 205607 479360
rect 196022 479302 205607 479304
rect 215342 479362 215402 479438
rect 231761 479496 234722 479498
rect 231761 479440 231766 479496
rect 231822 479440 234722 479496
rect 231761 479438 234722 479440
rect 231761 479435 231827 479438
rect 224861 479362 224927 479365
rect 215342 479360 224927 479362
rect 215342 479304 224866 479360
rect 224922 479304 224927 479360
rect 215342 479302 224927 479304
rect 234662 479362 234722 479438
rect 251081 479496 254042 479498
rect 251081 479440 251086 479496
rect 251142 479440 254042 479496
rect 251081 479438 254042 479440
rect 251081 479435 251147 479438
rect 244181 479362 244247 479365
rect 234662 479360 244247 479362
rect 234662 479304 244186 479360
rect 244242 479304 244247 479360
rect 234662 479302 244247 479304
rect 253982 479362 254042 479438
rect 270542 479496 278839 479498
rect 270542 479440 278778 479496
rect 278834 479440 278839 479496
rect 270542 479438 278839 479440
rect 253982 479302 263426 479362
rect 128261 479299 128327 479302
rect 147581 479299 147647 479302
rect 166901 479299 166967 479302
rect 186221 479299 186287 479302
rect 205541 479299 205607 479302
rect 224861 479299 224927 479302
rect 244181 479299 244247 479302
rect 86902 479164 86908 479228
rect 86972 479226 86978 479228
rect 96470 479226 96476 479228
rect 86972 479166 96476 479226
rect 86972 479164 86978 479166
rect 96470 479164 96476 479166
rect 96540 479164 96546 479228
rect 99465 479226 99531 479229
rect 106222 479226 106228 479228
rect 99465 479224 106228 479226
rect 99465 479168 99470 479224
rect 99526 479168 106228 479224
rect 99465 479166 106228 479168
rect 99465 479163 99531 479166
rect 106222 479164 106228 479166
rect 106292 479164 106298 479228
rect 263366 479090 263426 479302
rect 269062 479300 269068 479364
rect 269132 479362 269138 479364
rect 270542 479362 270602 479438
rect 278773 479435 278839 479438
rect 283557 479498 283623 479501
rect 292438 479498 292498 479574
rect 283557 479496 292498 479498
rect 283557 479440 283562 479496
rect 283618 479440 292498 479496
rect 283557 479438 292498 479440
rect 283557 479435 283623 479438
rect 269132 479302 270602 479362
rect 302374 479362 302434 479574
rect 316769 479632 318748 479634
rect 316769 479576 316774 479632
rect 316830 479576 318748 479632
rect 316769 479574 318748 479576
rect 316769 479571 316835 479574
rect 318742 479572 318748 479574
rect 318812 479572 318818 479636
rect 339726 479574 347698 479634
rect 309133 479362 309199 479365
rect 302374 479360 309199 479362
rect 302374 479304 309138 479360
rect 309194 479304 309199 479360
rect 302374 479302 309199 479304
rect 269132 479300 269138 479302
rect 309133 479299 309199 479302
rect 318742 479300 318748 479364
rect 318812 479362 318818 479364
rect 321369 479362 321435 479365
rect 318812 479360 321435 479362
rect 318812 479304 321374 479360
rect 321430 479304 321435 479360
rect 318812 479302 321435 479304
rect 318812 479300 318818 479302
rect 321369 479299 321435 479302
rect 321553 479362 321619 479365
rect 339726 479362 339786 479574
rect 321553 479360 321754 479362
rect 321553 479304 321558 479360
rect 321614 479304 321754 479360
rect 321553 479302 321754 479304
rect 321553 479299 321619 479302
rect 321694 479226 321754 479302
rect 331262 479302 339786 479362
rect 331262 479226 331322 479302
rect 321694 479166 331322 479226
rect 347638 479226 347698 479574
rect 376702 479572 376708 479636
rect 376772 479634 376778 479636
rect 376772 479574 389282 479634
rect 376772 479572 376778 479574
rect 389222 479498 389282 479574
rect 415350 479574 424978 479634
rect 389222 479438 398850 479498
rect 350441 479362 350507 479365
rect 347822 479360 350507 479362
rect 347822 479304 350446 479360
rect 350502 479304 350507 479360
rect 347822 479302 350507 479304
rect 347822 479226 347882 479302
rect 350441 479299 350507 479302
rect 350625 479362 350691 479365
rect 357382 479362 357388 479364
rect 350625 479360 357388 479362
rect 350625 479304 350630 479360
rect 350686 479304 357388 479360
rect 350625 479302 357388 479304
rect 350625 479299 350691 479302
rect 357382 479300 357388 479302
rect 357452 479300 357458 479364
rect 347638 479166 347882 479226
rect 398790 479226 398850 479438
rect 415350 479362 415410 479574
rect 408542 479302 415410 479362
rect 408542 479226 408602 479302
rect 398790 479166 408602 479226
rect 424918 479226 424978 479574
rect 427813 479498 427879 479501
rect 434662 479498 434668 479500
rect 427813 479496 434668 479498
rect 427813 479440 427818 479496
rect 427874 479440 434668 479496
rect 427813 479438 434668 479440
rect 427813 479435 427879 479438
rect 434662 479436 434668 479438
rect 434732 479436 434738 479500
rect 444281 479498 444347 479501
rect 446998 479498 447058 479710
rect 463742 479634 463802 479710
rect 466361 479634 466427 479637
rect 463742 479632 466427 479634
rect 463742 479576 466366 479632
rect 466422 479576 466427 479632
rect 463742 479574 466427 479576
rect 466361 479571 466427 479574
rect 507117 479634 507183 479637
rect 511942 479634 511948 479636
rect 507117 479632 511948 479634
rect 507117 479576 507122 479632
rect 507178 479576 511948 479632
rect 507117 479574 511948 479576
rect 507117 479571 507183 479574
rect 511942 479572 511948 479574
rect 512012 479572 512018 479636
rect 519118 479572 519124 479636
rect 519188 479634 519194 479636
rect 519854 479634 519860 479636
rect 519188 479574 519860 479634
rect 519188 479572 519194 479574
rect 519854 479572 519860 479574
rect 519924 479572 519930 479636
rect 444281 479496 447058 479498
rect 444281 479440 444286 479496
rect 444342 479440 447058 479496
rect 444281 479438 447058 479440
rect 473261 479498 473327 479501
rect 492581 479498 492647 479501
rect 473261 479496 476130 479498
rect 473261 479440 473266 479496
rect 473322 479440 476130 479496
rect 473261 479438 476130 479440
rect 444281 479435 444347 479438
rect 473261 479435 473327 479438
rect 427721 479362 427787 479365
rect 427678 479360 427787 479362
rect 427678 479304 427726 479360
rect 427782 479304 427787 479360
rect 427678 479299 427787 479304
rect 427678 479226 427738 479299
rect 424918 479166 427738 479226
rect 476070 479226 476130 479438
rect 492581 479496 495450 479498
rect 492581 479440 492586 479496
rect 492642 479440 495450 479496
rect 492581 479438 495450 479440
rect 492581 479435 492647 479438
rect 485681 479362 485747 479365
rect 483062 479360 485747 479362
rect 483062 479304 485686 479360
rect 485742 479304 485747 479360
rect 483062 479302 485747 479304
rect 483062 479226 483122 479302
rect 485681 479299 485747 479302
rect 476070 479166 483122 479226
rect 495390 479226 495450 479438
rect 507117 479362 507183 479365
rect 502382 479360 507183 479362
rect 502382 479304 507122 479360
rect 507178 479304 507183 479360
rect 502382 479302 507183 479304
rect 502382 479226 502442 479302
rect 507117 479299 507183 479302
rect 511942 479300 511948 479364
rect 512012 479362 512018 479364
rect 519854 479362 519860 479364
rect 512012 479302 519860 479362
rect 512012 479300 512018 479302
rect 519854 479300 519860 479302
rect 519924 479300 519930 479364
rect 495390 479166 502442 479226
rect 269062 479090 269068 479092
rect 263366 479030 269068 479090
rect 269062 479028 269068 479030
rect 269132 479028 269138 479092
rect 519813 479090 519879 479093
rect 519813 479088 519922 479090
rect 519813 479032 519818 479088
rect 519874 479032 519922 479088
rect 519813 479027 519922 479032
rect 277393 478954 277459 478957
rect 277393 478952 280140 478954
rect 277393 478896 277398 478952
rect 277454 478896 280140 478952
rect 519862 478924 519922 479027
rect 277393 478894 280140 478896
rect 277393 478891 277459 478894
rect 522798 476914 522804 476916
rect 519892 476854 522804 476914
rect 522798 476852 522804 476854
rect 522868 476852 522874 476916
rect 277393 476778 277459 476781
rect 277393 476776 280140 476778
rect 277393 476720 277398 476776
rect 277454 476720 280140 476776
rect 277393 476718 280140 476720
rect 277393 476715 277459 476718
rect 520089 476234 520155 476237
rect 520406 476234 520412 476236
rect 520089 476232 520412 476234
rect 520089 476176 520094 476232
rect 520150 476176 520412 476232
rect 520089 476174 520412 476176
rect 520089 476171 520155 476174
rect 520406 476172 520412 476174
rect 520476 476172 520482 476236
rect 520089 476098 520155 476101
rect 520406 476098 520412 476100
rect 520089 476096 520412 476098
rect 520089 476040 520094 476096
rect 520150 476040 520412 476096
rect 520089 476038 520412 476040
rect 520089 476035 520155 476038
rect 520406 476036 520412 476038
rect 520476 476036 520482 476100
rect 519302 475764 519308 475828
rect 519372 475764 519378 475828
rect 519486 475764 519492 475828
rect 519556 475764 519562 475828
rect 519670 475764 519676 475828
rect 519740 475764 519746 475828
rect 519854 475764 519860 475828
rect 519924 475764 519930 475828
rect 519310 475556 519370 475764
rect 519494 475556 519554 475764
rect 519678 475556 519738 475764
rect 519862 475556 519922 475764
rect 519302 475492 519308 475556
rect 519372 475492 519378 475556
rect 519486 475492 519492 475556
rect 519556 475492 519562 475556
rect 519670 475492 519676 475556
rect 519740 475492 519746 475556
rect 519854 475492 519860 475556
rect 519924 475492 519930 475556
rect 583520 474996 584960 475236
rect 278681 474738 278747 474741
rect 521694 474738 521700 474740
rect 278681 474736 280140 474738
rect 278681 474680 278686 474736
rect 278742 474680 280140 474736
rect 278681 474678 280140 474680
rect 519892 474678 521700 474738
rect 278681 474675 278747 474678
rect 521694 474676 521700 474678
rect 521764 474676 521770 474740
rect 520222 472698 520228 472700
rect 519892 472638 520228 472698
rect 520222 472636 520228 472638
rect 520292 472636 520298 472700
rect 278681 472562 278747 472565
rect 278681 472560 280140 472562
rect 278681 472504 278686 472560
rect 278742 472504 280140 472560
rect 278681 472502 280140 472504
rect 278681 472499 278747 472502
rect 521878 470522 521884 470524
rect 519892 470462 521884 470522
rect 521878 470460 521884 470462
rect 521948 470460 521954 470524
rect 277853 470386 277919 470389
rect 277853 470384 280140 470386
rect 277853 470328 277858 470384
rect 277914 470328 280140 470384
rect 277853 470326 280140 470328
rect 277853 470323 277919 470326
rect 519302 468692 519308 468756
rect 519372 468754 519378 468756
rect 521326 468754 521332 468756
rect 519372 468694 521332 468754
rect 519372 468692 519378 468694
rect 521326 468692 521332 468694
rect 521396 468692 521402 468756
rect 519486 468556 519492 468620
rect 519556 468618 519562 468620
rect 521142 468618 521148 468620
rect 519556 468558 521148 468618
rect 519556 468556 519562 468558
rect 521142 468556 521148 468558
rect 521212 468556 521218 468620
rect 522062 468482 522068 468484
rect 519892 468422 522068 468482
rect 522062 468420 522068 468422
rect 522132 468420 522138 468484
rect 278681 468346 278747 468349
rect 278681 468344 280140 468346
rect 278681 468288 278686 468344
rect 278742 468288 280140 468344
rect 278681 468286 280140 468288
rect 278681 468283 278747 468286
rect -960 466700 480 466940
rect 519854 466516 519860 466580
rect 519924 466578 519930 466580
rect 519924 466518 520842 466578
rect 519924 466516 519930 466518
rect 519670 466380 519676 466444
rect 519740 466442 519746 466444
rect 519740 466382 520658 466442
rect 519740 466380 519746 466382
rect 520406 466306 520412 466308
rect 519892 466246 520412 466306
rect 520406 466244 520412 466246
rect 520476 466244 520482 466308
rect 278681 466170 278747 466173
rect 278681 466168 280140 466170
rect 278681 466112 278686 466168
rect 278742 466112 280140 466168
rect 278681 466110 280140 466112
rect 278681 466107 278747 466110
rect 519670 465972 519676 466036
rect 519740 466034 519746 466036
rect 520598 466034 520658 466382
rect 519740 465974 520658 466034
rect 519740 465972 519746 465974
rect 519854 465836 519860 465900
rect 519924 465898 519930 465900
rect 520782 465898 520842 466518
rect 519924 465838 520842 465898
rect 519924 465836 519930 465838
rect 519486 465564 519492 465628
rect 519556 465626 519562 465628
rect 521142 465626 521148 465628
rect 519556 465566 521148 465626
rect 519556 465564 519562 465566
rect 521142 465564 521148 465566
rect 521212 465564 521218 465628
rect 519302 465428 519308 465492
rect 519372 465490 519378 465492
rect 521326 465490 521332 465492
rect 519372 465430 521332 465490
rect 519372 465428 519378 465430
rect 521326 465428 521332 465430
rect 521396 465428 521402 465492
rect 522246 464266 522252 464268
rect 519892 464206 522252 464266
rect 522246 464204 522252 464206
rect 522316 464204 522322 464268
rect 278681 464130 278747 464133
rect 278681 464128 280140 464130
rect 278681 464072 278686 464128
rect 278742 464072 280140 464128
rect 278681 464070 280140 464072
rect 278681 464067 278747 464070
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 522430 462090 522436 462092
rect 519892 462030 522436 462090
rect 522430 462028 522436 462030
rect 522500 462028 522506 462092
rect 278681 461954 278747 461957
rect 278681 461952 280140 461954
rect 278681 461896 278686 461952
rect 278742 461896 280140 461952
rect 278681 461894 280140 461896
rect 278681 461891 278747 461894
rect 521653 460050 521719 460053
rect 519892 460048 521719 460050
rect 519892 459992 521658 460048
rect 521714 459992 521719 460048
rect 519892 459990 521719 459992
rect 521653 459987 521719 459990
rect 278681 459778 278747 459781
rect 278681 459776 280140 459778
rect 278681 459720 278686 459776
rect 278742 459720 280140 459776
rect 278681 459718 280140 459720
rect 278681 459715 278747 459718
rect 522614 457874 522620 457876
rect 519892 457814 522620 457874
rect 522614 457812 522620 457814
rect 522684 457812 522690 457876
rect 278681 457738 278747 457741
rect 278681 457736 280140 457738
rect 278681 457680 278686 457736
rect 278742 457680 280140 457736
rect 278681 457678 280140 457680
rect 278681 457675 278747 457678
rect 521745 455834 521811 455837
rect 519892 455832 521811 455834
rect 519892 455776 521750 455832
rect 521806 455776 521811 455832
rect 519892 455774 521811 455776
rect 521745 455771 521811 455774
rect 278681 455562 278747 455565
rect 278681 455560 280140 455562
rect 278681 455504 278686 455560
rect 278742 455504 280140 455560
rect 278681 455502 280140 455504
rect 278681 455499 278747 455502
rect 542353 454066 542419 454069
rect 542629 454066 542695 454069
rect 542353 454064 542695 454066
rect 542353 454008 542358 454064
rect 542414 454008 542634 454064
rect 542690 454008 542695 454064
rect 542353 454006 542695 454008
rect 542353 454003 542419 454006
rect 542629 454003 542695 454006
rect 521837 453658 521903 453661
rect 519892 453656 521903 453658
rect 519892 453600 521842 453656
rect 521898 453600 521903 453656
rect 519892 453598 521903 453600
rect 521837 453595 521903 453598
rect 278681 453386 278747 453389
rect 278681 453384 280140 453386
rect 278681 453328 278686 453384
rect 278742 453328 280140 453384
rect 278681 453326 280140 453328
rect 278681 453323 278747 453326
rect 519486 452644 519492 452708
rect 519556 452644 519562 452708
rect 519670 452644 519676 452708
rect 519740 452644 519746 452708
rect 519854 452644 519860 452708
rect 519924 452644 519930 452708
rect -960 452434 480 452524
rect 3509 452434 3575 452437
rect 519494 452436 519554 452644
rect 519678 452436 519738 452644
rect 519862 452436 519922 452644
rect -960 452432 3575 452434
rect -960 452376 3514 452432
rect 3570 452376 3575 452432
rect -960 452374 3575 452376
rect -960 452284 480 452374
rect 3509 452371 3575 452374
rect 519486 452372 519492 452436
rect 519556 452372 519562 452436
rect 519670 452372 519676 452436
rect 519740 452372 519746 452436
rect 519854 452372 519860 452436
rect 519924 452372 519930 452436
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 521929 451618 521995 451621
rect 519892 451616 521995 451618
rect 519892 451560 521934 451616
rect 521990 451560 521995 451616
rect 583520 451604 584960 451694
rect 519892 451558 521995 451560
rect 521929 451555 521995 451558
rect 278681 451346 278747 451349
rect 278681 451344 280140 451346
rect 278681 451288 278686 451344
rect 278742 451288 280140 451344
rect 278681 451286 280140 451288
rect 278681 451283 278747 451286
rect 522021 449442 522087 449445
rect 519892 449440 522087 449442
rect 519892 449384 522026 449440
rect 522082 449384 522087 449440
rect 519892 449382 522087 449384
rect 522021 449379 522087 449382
rect 278681 449170 278747 449173
rect 278681 449168 280140 449170
rect 278681 449112 278686 449168
rect 278742 449112 280140 449168
rect 278681 449110 280140 449112
rect 278681 449107 278747 449110
rect 522113 447402 522179 447405
rect 519892 447400 522179 447402
rect 519892 447344 522118 447400
rect 522174 447344 522179 447400
rect 519892 447342 522179 447344
rect 522113 447339 522179 447342
rect 278681 447130 278747 447133
rect 278681 447128 280140 447130
rect 278681 447072 278686 447128
rect 278742 447072 280140 447128
rect 278681 447070 280140 447072
rect 278681 447067 278747 447070
rect 522941 445226 523007 445229
rect 519892 445224 523007 445226
rect 519892 445168 522946 445224
rect 523002 445168 523007 445224
rect 519892 445166 523007 445168
rect 522941 445163 523007 445166
rect 278681 444954 278747 444957
rect 278681 444952 280140 444954
rect 278681 444896 278686 444952
rect 278742 444896 280140 444952
rect 278681 444894 280140 444896
rect 278681 444891 278747 444894
rect 522205 443186 522271 443189
rect 519892 443184 522271 443186
rect 519892 443128 522210 443184
rect 522266 443128 522271 443184
rect 519892 443126 522271 443128
rect 522205 443123 522271 443126
rect 277853 442778 277919 442781
rect 277853 442776 280140 442778
rect 277853 442720 277858 442776
rect 277914 442720 280140 442776
rect 277853 442718 280140 442720
rect 277853 442715 277919 442718
rect 522389 441010 522455 441013
rect 519892 441008 522455 441010
rect 519892 440952 522394 441008
rect 522450 440952 522455 441008
rect 519892 440950 522455 440952
rect 522389 440947 522455 440950
rect 278681 440738 278747 440741
rect 278681 440736 280140 440738
rect 278681 440680 278686 440736
rect 278742 440680 280140 440736
rect 278681 440678 280140 440680
rect 278681 440675 278747 440678
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect 522389 438970 522455 438973
rect 519892 438968 522455 438970
rect 519892 438912 522394 438968
rect 522450 438912 522455 438968
rect 519892 438910 522455 438912
rect 522389 438907 522455 438910
rect 278681 438562 278747 438565
rect 278681 438560 280140 438562
rect 278681 438504 278686 438560
rect 278742 438504 280140 438560
rect 278681 438502 280140 438504
rect 278681 438499 278747 438502
rect -960 438018 480 438108
rect 3509 438018 3575 438021
rect -960 438016 3575 438018
rect -960 437960 3514 438016
rect 3570 437960 3575 438016
rect -960 437958 3575 437960
rect -960 437868 480 437958
rect 3509 437955 3575 437958
rect 520038 437684 520044 437748
rect 520108 437746 520114 437748
rect 521142 437746 521148 437748
rect 520108 437686 521148 437746
rect 520108 437684 520114 437686
rect 521142 437684 521148 437686
rect 521212 437684 521218 437748
rect 519813 437610 519879 437613
rect 520038 437610 520044 437612
rect 519813 437608 520044 437610
rect 519813 437552 519818 437608
rect 519874 437552 520044 437608
rect 519813 437550 520044 437552
rect 519813 437547 519879 437550
rect 520038 437548 520044 437550
rect 520108 437548 520114 437612
rect 522849 436794 522915 436797
rect 519892 436792 522915 436794
rect 519892 436736 522854 436792
rect 522910 436736 522915 436792
rect 519892 436734 522915 436736
rect 522849 436731 522915 436734
rect 278037 436386 278103 436389
rect 278037 436384 280140 436386
rect 278037 436328 278042 436384
rect 278098 436328 280140 436384
rect 278037 436326 280140 436328
rect 278037 436323 278103 436326
rect 520038 435298 520044 435300
rect 519862 435238 520044 435298
rect 519862 434724 519922 435238
rect 520038 435236 520044 435238
rect 520108 435236 520114 435300
rect 520038 435100 520044 435164
rect 520108 435162 520114 435164
rect 521142 435162 521148 435164
rect 520108 435102 521148 435162
rect 520108 435100 520114 435102
rect 521142 435100 521148 435102
rect 521212 435100 521218 435164
rect 542169 434754 542235 434757
rect 542353 434754 542419 434757
rect 542169 434752 542419 434754
rect 542169 434696 542174 434752
rect 542230 434696 542358 434752
rect 542414 434696 542419 434752
rect 542169 434694 542419 434696
rect 542169 434691 542235 434694
rect 542353 434691 542419 434694
rect 278681 434346 278747 434349
rect 278681 434344 280140 434346
rect 278681 434288 278686 434344
rect 278742 434288 280140 434344
rect 278681 434286 280140 434288
rect 278681 434283 278747 434286
rect 521561 432578 521627 432581
rect 519892 432576 521627 432578
rect 519892 432520 521566 432576
rect 521622 432520 521627 432576
rect 519892 432518 521627 432520
rect 521561 432515 521627 432518
rect 278681 432170 278747 432173
rect 278681 432168 280140 432170
rect 278681 432112 278686 432168
rect 278742 432112 280140 432168
rect 278681 432110 280140 432112
rect 278681 432107 278747 432110
rect 522665 430538 522731 430541
rect 519892 430536 522731 430538
rect 519892 430480 522670 430536
rect 522726 430480 522731 430536
rect 519892 430478 522731 430480
rect 522665 430475 522731 430478
rect 277669 430130 277735 430133
rect 277669 430128 280140 430130
rect 277669 430072 277674 430128
rect 277730 430072 280140 430128
rect 277669 430070 280140 430072
rect 277669 430067 277735 430070
rect 520038 429796 520044 429860
rect 520108 429858 520114 429860
rect 521142 429858 521148 429860
rect 520108 429798 521148 429858
rect 520108 429796 520114 429798
rect 521142 429796 521148 429798
rect 521212 429796 521218 429860
rect 519670 429660 519676 429724
rect 519740 429722 519746 429724
rect 520038 429722 520044 429724
rect 519740 429662 520044 429722
rect 519740 429660 519746 429662
rect 520038 429660 520044 429662
rect 520108 429660 520114 429724
rect 519862 428438 520474 428498
rect 519862 428332 519922 428438
rect 520414 428362 520474 428438
rect 523125 428362 523191 428365
rect 520414 428360 523191 428362
rect 520414 428304 523130 428360
rect 523186 428304 523191 428360
rect 520414 428302 523191 428304
rect 523125 428299 523191 428302
rect 520038 428090 520044 428092
rect 519678 428030 520044 428090
rect 278681 427954 278747 427957
rect 519678 427956 519738 428030
rect 520038 428028 520044 428030
rect 520108 428028 520114 428092
rect 583520 428076 584960 428316
rect 278681 427952 280140 427954
rect 278681 427896 278686 427952
rect 278742 427896 280140 427952
rect 278681 427894 280140 427896
rect 278681 427891 278747 427894
rect 519670 427892 519676 427956
rect 519740 427892 519746 427956
rect 522941 426322 523007 426325
rect 519892 426320 523007 426322
rect 519892 426264 522946 426320
rect 523002 426264 523007 426320
rect 519892 426262 523007 426264
rect 522941 426259 523007 426262
rect 278681 425778 278747 425781
rect 278681 425776 280140 425778
rect 278681 425720 278686 425776
rect 278742 425720 280140 425776
rect 278681 425718 280140 425720
rect 278681 425715 278747 425718
rect 520038 425036 520044 425100
rect 520108 425098 520114 425100
rect 521142 425098 521148 425100
rect 520108 425038 521148 425098
rect 520108 425036 520114 425038
rect 521142 425036 521148 425038
rect 521212 425036 521218 425100
rect 521469 424146 521535 424149
rect 519892 424144 521535 424146
rect 519892 424088 521474 424144
rect 521530 424088 521535 424144
rect 519892 424086 521535 424088
rect 521469 424083 521535 424086
rect -960 423738 480 423828
rect 3233 423738 3299 423741
rect -960 423736 3299 423738
rect -960 423680 3238 423736
rect 3294 423680 3299 423736
rect -960 423678 3299 423680
rect -960 423588 480 423678
rect 3233 423675 3299 423678
rect 278681 423738 278747 423741
rect 278681 423736 280140 423738
rect 278681 423680 278686 423736
rect 278742 423680 280140 423736
rect 278681 423678 280140 423680
rect 278681 423675 278747 423678
rect 522757 422106 522823 422109
rect 519892 422104 522823 422106
rect 519892 422048 522762 422104
rect 522818 422048 522823 422104
rect 519892 422046 522823 422048
rect 522757 422043 522823 422046
rect 278681 421562 278747 421565
rect 278681 421560 280140 421562
rect 278681 421504 278686 421560
rect 278742 421504 280140 421560
rect 278681 421502 280140 421504
rect 278681 421499 278747 421502
rect 522665 420066 522731 420069
rect 519892 420064 522731 420066
rect 519892 420008 522670 420064
rect 522726 420008 522731 420064
rect 519892 420006 522731 420008
rect 522665 420003 522731 420006
rect 278681 419522 278747 419525
rect 278681 419520 280140 419522
rect 278681 419464 278686 419520
rect 278742 419464 280140 419520
rect 278681 419462 280140 419464
rect 278681 419459 278747 419462
rect 520181 417890 520247 417893
rect 519892 417888 520247 417890
rect 519892 417832 520186 417888
rect 520242 417832 520247 417888
rect 519892 417830 520247 417832
rect 520181 417827 520247 417830
rect 278681 417346 278747 417349
rect 278681 417344 280140 417346
rect 278681 417288 278686 417344
rect 278742 417288 280140 417344
rect 278681 417286 280140 417288
rect 278681 417283 278747 417286
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 521285 415850 521351 415853
rect 519892 415848 521351 415850
rect 519892 415792 521290 415848
rect 521346 415792 521351 415848
rect 519892 415790 521351 415792
rect 521285 415787 521351 415790
rect 519302 415516 519308 415580
rect 519372 415516 519378 415580
rect 277853 415170 277919 415173
rect 277853 415168 280140 415170
rect 277853 415112 277858 415168
rect 277914 415112 280140 415168
rect 277853 415110 280140 415112
rect 277853 415107 277919 415110
rect 519310 415036 519370 415516
rect 542169 415442 542235 415445
rect 542353 415442 542419 415445
rect 542169 415440 542419 415442
rect 542169 415384 542174 415440
rect 542230 415384 542358 415440
rect 542414 415384 542419 415440
rect 542169 415382 542419 415384
rect 542169 415379 542235 415382
rect 542353 415379 542419 415382
rect 519486 415244 519492 415308
rect 519556 415306 519562 415308
rect 519556 415246 519738 415306
rect 519556 415244 519562 415246
rect 519302 414972 519308 415036
rect 519372 414972 519378 415036
rect 519678 414898 519738 415246
rect 519854 415244 519860 415308
rect 519924 415244 519930 415308
rect 519862 415036 519922 415244
rect 519854 414972 519860 415036
rect 519924 414972 519930 415036
rect 520181 414898 520247 414901
rect 519678 414896 520247 414898
rect 519678 414840 520186 414896
rect 520242 414840 520247 414896
rect 519678 414838 520247 414840
rect 520181 414835 520247 414838
rect 520089 413674 520155 413677
rect 519892 413672 520155 413674
rect 519892 413616 520094 413672
rect 520150 413616 520155 413672
rect 519892 413614 520155 413616
rect 520089 413611 520155 413614
rect 278681 413130 278747 413133
rect 278681 413128 280140 413130
rect 278681 413072 278686 413128
rect 278742 413072 280140 413128
rect 278681 413070 280140 413072
rect 278681 413067 278747 413070
rect 519997 412178 520063 412181
rect 519862 412176 520063 412178
rect 519862 412120 520002 412176
rect 520058 412120 520063 412176
rect 519862 412118 520063 412120
rect 519862 411604 519922 412118
rect 519997 412115 520063 412118
rect 278681 410954 278747 410957
rect 278681 410952 280140 410954
rect 278681 410896 278686 410952
rect 278742 410896 280140 410952
rect 278681 410894 280140 410896
rect 278681 410891 278747 410894
rect 522573 409458 522639 409461
rect 519892 409456 522639 409458
rect -960 409172 480 409412
rect 519892 409400 522578 409456
rect 522634 409400 522639 409456
rect 519892 409398 522639 409400
rect 522573 409395 522639 409398
rect 519302 409124 519308 409188
rect 519372 409186 519378 409188
rect 519997 409186 520063 409189
rect 519372 409184 520063 409186
rect 519372 409128 520002 409184
rect 520058 409128 520063 409184
rect 519372 409126 520063 409128
rect 519372 409124 519378 409126
rect 519997 409123 520063 409126
rect 278681 408778 278747 408781
rect 519670 408778 519676 408780
rect 278681 408776 280140 408778
rect 278681 408720 278686 408776
rect 278742 408720 280140 408776
rect 278681 408718 280140 408720
rect 519310 408718 519676 408778
rect 278681 408715 278747 408718
rect 519310 408370 519370 408718
rect 519670 408716 519676 408718
rect 519740 408716 519746 408780
rect 519670 408370 519676 408372
rect 519310 408310 519676 408370
rect 519670 408308 519676 408310
rect 519740 408308 519746 408372
rect 522481 407418 522547 407421
rect 519892 407416 522547 407418
rect 519892 407360 522486 407416
rect 522542 407360 522547 407416
rect 519892 407358 522547 407360
rect 522481 407355 522547 407358
rect 519302 406948 519308 407012
rect 519372 407010 519378 407012
rect 520038 407010 520044 407012
rect 519372 406950 520044 407010
rect 519372 406948 519378 406950
rect 520038 406948 520044 406950
rect 520108 406948 520114 407012
rect 278681 406738 278747 406741
rect 278681 406736 280140 406738
rect 278681 406680 278686 406736
rect 278742 406680 280140 406736
rect 278681 406678 280140 406680
rect 278681 406675 278747 406678
rect 519486 406330 519492 406332
rect 519310 406270 519492 406330
rect 519310 406196 519370 406270
rect 519486 406268 519492 406270
rect 519556 406268 519562 406332
rect 519302 406132 519308 406196
rect 519372 406132 519378 406196
rect 519486 406132 519492 406196
rect 519556 406194 519562 406196
rect 520181 406194 520247 406197
rect 519556 406192 520247 406194
rect 519556 406136 520186 406192
rect 520242 406136 520247 406192
rect 519556 406134 520247 406136
rect 519556 406132 519562 406134
rect 520181 406131 520247 406134
rect 519302 405996 519308 406060
rect 519372 406058 519378 406060
rect 519997 406058 520063 406061
rect 519372 406056 520063 406058
rect 519372 406000 520002 406056
rect 520058 406000 520063 406056
rect 519372 405998 520063 406000
rect 519372 405996 519378 405998
rect 519997 405995 520063 405998
rect 521377 405242 521443 405245
rect 519892 405240 521443 405242
rect 519892 405184 521382 405240
rect 521438 405184 521443 405240
rect 519892 405182 521443 405184
rect 521377 405179 521443 405182
rect 580257 404834 580323 404837
rect 583520 404834 584960 404924
rect 580257 404832 584960 404834
rect 580257 404776 580262 404832
rect 580318 404776 584960 404832
rect 580257 404774 584960 404776
rect 580257 404771 580323 404774
rect 583520 404684 584960 404774
rect 278681 404562 278747 404565
rect 278681 404560 280140 404562
rect 278681 404504 278686 404560
rect 278742 404504 280140 404560
rect 278681 404502 280140 404504
rect 278681 404499 278747 404502
rect 520825 403202 520891 403205
rect 519892 403200 520891 403202
rect 519892 403144 520830 403200
rect 520886 403144 520891 403200
rect 519892 403142 520891 403144
rect 520825 403139 520891 403142
rect 278405 402522 278471 402525
rect 278405 402520 280140 402522
rect 278405 402464 278410 402520
rect 278466 402464 280140 402520
rect 278405 402462 280140 402464
rect 278405 402459 278471 402462
rect 522297 401026 522363 401029
rect 519892 401024 522363 401026
rect 519892 400968 522302 401024
rect 522358 400968 522363 401024
rect 519892 400966 522363 400968
rect 522297 400963 522363 400966
rect 278681 400346 278747 400349
rect 278681 400344 280140 400346
rect 278681 400288 278686 400344
rect 278742 400288 280140 400344
rect 278681 400286 280140 400288
rect 278681 400283 278747 400286
rect 519670 399468 519676 399532
rect 519740 399468 519746 399532
rect 519678 398956 519738 399468
rect 278681 398170 278747 398173
rect 278681 398168 280140 398170
rect 278681 398112 278686 398168
rect 278742 398112 280140 398168
rect 278681 398110 280140 398112
rect 278681 398107 278747 398110
rect 520958 396810 520964 396812
rect 519892 396750 520964 396810
rect 520958 396748 520964 396750
rect 521028 396748 521034 396812
rect 519302 396340 519308 396404
rect 519372 396402 519378 396404
rect 519997 396402 520063 396405
rect 519372 396400 520063 396402
rect 519372 396344 520002 396400
rect 520058 396344 520063 396400
rect 519372 396342 520063 396344
rect 519372 396340 519378 396342
rect 519997 396339 520063 396342
rect 278681 396130 278747 396133
rect 278681 396128 280140 396130
rect 278681 396072 278686 396128
rect 278742 396072 280140 396128
rect 278681 396070 280140 396072
rect 278681 396067 278747 396070
rect 519302 395524 519308 395588
rect 519372 395586 519378 395588
rect 520089 395586 520155 395589
rect 519372 395584 520155 395586
rect 519372 395528 520094 395584
rect 520150 395528 520155 395584
rect 519372 395526 520155 395528
rect 519372 395524 519378 395526
rect 520089 395523 520155 395526
rect 519486 395252 519492 395316
rect 519556 395252 519562 395316
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 519494 394740 519554 395252
rect 542077 394770 542143 394773
rect 542261 394770 542327 394773
rect 542077 394768 542327 394770
rect 542077 394712 542082 394768
rect 542138 394712 542266 394768
rect 542322 394712 542327 394768
rect 542077 394710 542327 394712
rect 542077 394707 542143 394710
rect 542261 394707 542327 394710
rect 278681 393954 278747 393957
rect 278681 393952 280140 393954
rect 278681 393896 278686 393952
rect 278742 393896 280140 393952
rect 278681 393894 280140 393896
rect 278681 393891 278747 393894
rect 519302 393348 519308 393412
rect 519372 393410 519378 393412
rect 519670 393410 519676 393412
rect 519372 393350 519676 393410
rect 519372 393348 519378 393350
rect 519670 393348 519676 393350
rect 519740 393348 519746 393412
rect 519997 393138 520063 393141
rect 519862 393136 520063 393138
rect 519862 393080 520002 393136
rect 520058 393080 520063 393136
rect 519862 393078 520063 393080
rect 519862 392564 519922 393078
rect 519997 393075 520063 393078
rect 579889 393002 579955 393005
rect 583520 393002 584960 393092
rect 579889 393000 584960 393002
rect 579889 392944 579894 393000
rect 579950 392944 584960 393000
rect 579889 392942 584960 392944
rect 579889 392939 579955 392942
rect 583520 392852 584960 392942
rect 278313 391778 278379 391781
rect 278313 391776 280140 391778
rect 278313 391720 278318 391776
rect 278374 391720 280140 391776
rect 278313 391718 280140 391720
rect 278313 391715 278379 391718
rect 519302 390628 519308 390692
rect 519372 390690 519378 390692
rect 520089 390690 520155 390693
rect 519372 390688 520155 390690
rect 519372 390632 520094 390688
rect 520150 390632 520155 390688
rect 519372 390630 520155 390632
rect 519372 390628 519378 390630
rect 520089 390627 520155 390630
rect 520774 390554 520780 390556
rect 519892 390494 520780 390554
rect 520774 390492 520780 390494
rect 520844 390492 520850 390556
rect 278681 389738 278747 389741
rect 278681 389736 280140 389738
rect 278681 389680 278686 389736
rect 278742 389680 280140 389736
rect 278681 389678 280140 389680
rect 278681 389675 278747 389678
rect 519670 388860 519676 388924
rect 519740 388860 519746 388924
rect 519678 388348 519738 388860
rect 277853 387562 277919 387565
rect 277853 387560 280140 387562
rect 277853 387504 277858 387560
rect 277914 387504 280140 387560
rect 277853 387502 280140 387504
rect 277853 387499 277919 387502
rect 519862 386068 519922 386308
rect 519854 386004 519860 386068
rect 519924 386004 519930 386068
rect 277669 385522 277735 385525
rect 277669 385520 280140 385522
rect 277669 385464 277674 385520
rect 277730 385464 280140 385520
rect 277669 385462 280140 385464
rect 277669 385459 277735 385462
rect 520590 384162 520596 384164
rect 519892 384102 520596 384162
rect 520590 384100 520596 384102
rect 520660 384100 520666 384164
rect 278681 383346 278747 383349
rect 278681 383344 280140 383346
rect 278681 383288 278686 383344
rect 278742 383288 280140 383344
rect 278681 383286 280140 383288
rect 278681 383283 278747 383286
rect 519302 382196 519308 382260
rect 519372 382196 519378 382260
rect 519310 382092 519370 382196
rect 278037 381170 278103 381173
rect 278037 381168 280140 381170
rect 278037 381112 278042 381168
rect 278098 381112 280140 381168
rect 583520 381156 584960 381396
rect 278037 381110 280140 381112
rect 278037 381107 278103 381110
rect -960 380626 480 380716
rect 3509 380626 3575 380629
rect -960 380624 3575 380626
rect -960 380568 3514 380624
rect 3570 380568 3575 380624
rect -960 380566 3575 380568
rect -960 380476 480 380566
rect 3509 380563 3575 380566
rect 521193 379946 521259 379949
rect 519892 379944 521259 379946
rect 519892 379888 521198 379944
rect 521254 379888 521259 379944
rect 519892 379886 521259 379888
rect 521193 379883 521259 379886
rect 278681 379130 278747 379133
rect 278681 379128 280140 379130
rect 278681 379072 278686 379128
rect 278742 379072 280140 379128
rect 278681 379070 280140 379072
rect 278681 379067 278747 379070
rect 520457 377906 520523 377909
rect 519892 377904 520523 377906
rect 519892 377848 520462 377904
rect 520518 377848 520523 377904
rect 519892 377846 520523 377848
rect 520457 377843 520523 377846
rect 278681 376954 278747 376957
rect 278681 376952 280140 376954
rect 278681 376896 278686 376952
rect 278742 376896 280140 376952
rect 278681 376894 280140 376896
rect 278681 376891 278747 376894
rect 519537 376274 519603 376277
rect 519494 376272 519603 376274
rect 519494 376216 519542 376272
rect 519598 376216 519603 376272
rect 519494 376211 519603 376216
rect 519494 375700 519554 376211
rect 278405 374914 278471 374917
rect 278405 374912 280140 374914
rect 278405 374856 278410 374912
rect 278466 374856 280140 374912
rect 278405 374854 280140 374856
rect 278405 374851 278471 374854
rect 521101 373690 521167 373693
rect 519892 373688 521167 373690
rect 519892 373632 521106 373688
rect 521162 373632 521167 373688
rect 519892 373630 521167 373632
rect 521101 373627 521167 373630
rect 278037 372738 278103 372741
rect 278037 372736 280140 372738
rect 278037 372680 278042 372736
rect 278098 372680 280140 372736
rect 278037 372678 280140 372680
rect 278037 372675 278103 372678
rect 519445 372058 519511 372061
rect 519445 372056 519554 372058
rect 519445 372000 519450 372056
rect 519506 372000 519554 372056
rect 519445 371995 519554 372000
rect 519494 371484 519554 371995
rect 278313 370562 278379 370565
rect 278313 370560 280140 370562
rect 278313 370504 278318 370560
rect 278374 370504 280140 370560
rect 278313 370502 280140 370504
rect 278313 370499 278379 370502
rect 519353 369746 519419 369749
rect 519310 369744 519419 369746
rect 519310 369688 519358 369744
rect 519414 369688 519419 369744
rect 519310 369683 519419 369688
rect 519310 369444 519370 369683
rect 580349 369610 580415 369613
rect 583520 369610 584960 369700
rect 580349 369608 584960 369610
rect 580349 369552 580354 369608
rect 580410 369552 584960 369608
rect 580349 369550 584960 369552
rect 580349 369547 580415 369550
rect 583520 369460 584960 369550
rect 278681 368522 278747 368525
rect 278681 368520 280140 368522
rect 278681 368464 278686 368520
rect 278742 368464 280140 368520
rect 278681 368462 280140 368464
rect 278681 368459 278747 368462
rect 521009 367298 521075 367301
rect 519892 367296 521075 367298
rect 519892 367240 521014 367296
rect 521070 367240 521075 367296
rect 519892 367238 521075 367240
rect 521009 367235 521075 367238
rect 278681 366346 278747 366349
rect 278681 366344 280140 366346
rect -960 366210 480 366300
rect 278681 366288 278686 366344
rect 278742 366288 280140 366344
rect 278681 366286 280140 366288
rect 278681 366283 278747 366286
rect 3509 366210 3575 366213
rect -960 366208 3575 366210
rect -960 366152 3514 366208
rect 3570 366152 3575 366208
rect -960 366150 3575 366152
rect -960 366060 480 366150
rect 3509 366147 3575 366150
rect 520365 365258 520431 365261
rect 519892 365256 520431 365258
rect 519892 365200 520370 365256
rect 520426 365200 520431 365256
rect 519892 365198 520431 365200
rect 520365 365195 520431 365198
rect 277853 364170 277919 364173
rect 277853 364168 280140 364170
rect 277853 364112 277858 364168
rect 277914 364112 280140 364168
rect 277853 364110 280140 364112
rect 277853 364107 277919 364110
rect 519353 363490 519419 363493
rect 519310 363488 519419 363490
rect 519310 363432 519358 363488
rect 519414 363432 519419 363488
rect 519310 363427 519419 363432
rect 519310 363052 519370 363427
rect 278681 362130 278747 362133
rect 278681 362128 280140 362130
rect 278681 362072 278686 362128
rect 278742 362072 280140 362128
rect 278681 362070 280140 362072
rect 278681 362067 278747 362070
rect 520917 361042 520983 361045
rect 519892 361040 520983 361042
rect 519892 360984 520922 361040
rect 520978 360984 520983 361040
rect 519892 360982 520983 360984
rect 520917 360979 520983 360982
rect 277853 359954 277919 359957
rect 277853 359952 280140 359954
rect 277853 359896 277858 359952
rect 277914 359896 280140 359952
rect 277853 359894 280140 359896
rect 277853 359891 277919 359894
rect 520273 359002 520339 359005
rect 519892 359000 520339 359002
rect 519892 358944 520278 359000
rect 520334 358944 520339 359000
rect 519892 358942 520339 358944
rect 520273 358939 520339 358942
rect 278681 357914 278747 357917
rect 580441 357914 580507 357917
rect 583520 357914 584960 358004
rect 278681 357912 280140 357914
rect 278681 357856 278686 357912
rect 278742 357856 280140 357912
rect 278681 357854 280140 357856
rect 580441 357912 584960 357914
rect 580441 357856 580446 357912
rect 580502 357856 584960 357912
rect 580441 357854 584960 357856
rect 278681 357851 278747 357854
rect 580441 357851 580507 357854
rect 583520 357764 584960 357854
rect 519721 357370 519787 357373
rect 519678 357368 519787 357370
rect 519678 357312 519726 357368
rect 519782 357312 519787 357368
rect 519678 357307 519787 357312
rect 519678 356796 519738 357307
rect 278681 355738 278747 355741
rect 278681 355736 280140 355738
rect 278681 355680 278686 355736
rect 278742 355680 280140 355736
rect 278681 355678 280140 355680
rect 278681 355675 278747 355678
rect 520733 354786 520799 354789
rect 519892 354784 520799 354786
rect 519892 354728 520738 354784
rect 520794 354728 520799 354784
rect 519892 354726 520799 354728
rect 520733 354723 520799 354726
rect 278037 353562 278103 353565
rect 278037 353560 280140 353562
rect 278037 353504 278042 353560
rect 278098 353504 280140 353560
rect 278037 353502 280140 353504
rect 278037 353499 278103 353502
rect 519353 353018 519419 353021
rect 519310 353016 519419 353018
rect 519310 352960 519358 353016
rect 519414 352960 519419 353016
rect 519310 352955 519419 352960
rect 519310 352580 519370 352955
rect -960 351780 480 352020
rect 278681 351522 278747 351525
rect 278681 351520 280140 351522
rect 278681 351464 278686 351520
rect 278742 351464 280140 351520
rect 278681 351462 280140 351464
rect 278681 351459 278747 351462
rect 519905 351114 519971 351117
rect 519862 351112 519971 351114
rect 519862 351056 519910 351112
rect 519966 351056 519971 351112
rect 519862 351051 519971 351056
rect 519862 350540 519922 351051
rect 278681 349346 278747 349349
rect 278681 349344 280140 349346
rect 278681 349288 278686 349344
rect 278742 349288 280140 349344
rect 278681 349286 280140 349288
rect 278681 349283 278747 349286
rect 520641 348394 520707 348397
rect 519892 348392 520707 348394
rect 519892 348336 520646 348392
rect 520702 348336 520707 348392
rect 519892 348334 520707 348336
rect 520641 348331 520707 348334
rect 278681 347170 278747 347173
rect 278681 347168 280140 347170
rect 278681 347112 278686 347168
rect 278742 347112 280140 347168
rect 278681 347110 280140 347112
rect 278681 347107 278747 347110
rect 519261 346490 519327 346493
rect 519261 346488 519370 346490
rect 519261 346432 519266 346488
rect 519322 346432 519370 346488
rect 519261 346427 519370 346432
rect 519310 346324 519370 346427
rect 580533 346082 580599 346085
rect 583520 346082 584960 346172
rect 580533 346080 584960 346082
rect 580533 346024 580538 346080
rect 580594 346024 584960 346080
rect 580533 346022 584960 346024
rect 580533 346019 580599 346022
rect 583520 345932 584960 346022
rect 278681 345130 278747 345133
rect 278681 345128 280140 345130
rect 278681 345072 278686 345128
rect 278742 345072 280140 345128
rect 278681 345070 280140 345072
rect 278681 345067 278747 345070
rect 519629 344586 519695 344589
rect 519629 344584 519738 344586
rect 519629 344528 519634 344584
rect 519690 344528 519738 344584
rect 519629 344523 519738 344528
rect 519678 344148 519738 344523
rect 278313 342954 278379 342957
rect 278313 342952 280140 342954
rect 278313 342896 278318 342952
rect 278374 342896 280140 342952
rect 278313 342894 280140 342896
rect 278313 342891 278379 342894
rect 520549 342138 520615 342141
rect 519892 342136 520615 342138
rect 519892 342080 520554 342136
rect 520610 342080 520615 342136
rect 519892 342078 520615 342080
rect 520549 342075 520615 342078
rect 278681 340914 278747 340917
rect 278681 340912 280140 340914
rect 278681 340856 278686 340912
rect 278742 340856 280140 340912
rect 278681 340854 280140 340856
rect 278681 340851 278747 340854
rect 522941 339962 523007 339965
rect 519892 339960 523007 339962
rect 519892 339904 522946 339960
rect 523002 339904 523007 339960
rect 519892 339902 523007 339904
rect 522941 339899 523007 339902
rect 278681 338738 278747 338741
rect 278681 338736 280140 338738
rect 278681 338680 278686 338736
rect 278742 338680 280140 338736
rect 278681 338678 280140 338680
rect 278681 338675 278747 338678
rect 522941 337922 523007 337925
rect 519892 337920 523007 337922
rect 519892 337864 522946 337920
rect 523002 337864 523007 337920
rect 519892 337862 523007 337864
rect 522941 337859 523007 337862
rect -960 337514 480 337604
rect 3509 337514 3575 337517
rect -960 337512 3575 337514
rect -960 337456 3514 337512
rect 3570 337456 3575 337512
rect -960 337454 3575 337456
rect -960 337364 480 337454
rect 3509 337451 3575 337454
rect 277853 336562 277919 336565
rect 277853 336560 280140 336562
rect 277853 336504 277858 336560
rect 277914 336504 280140 336560
rect 277853 336502 280140 336504
rect 277853 336499 277919 336502
rect 522573 335746 522639 335749
rect 519892 335744 522639 335746
rect 519892 335688 522578 335744
rect 522634 335688 522639 335744
rect 519892 335686 522639 335688
rect 522573 335683 522639 335686
rect 278681 334522 278747 334525
rect 278681 334520 280140 334522
rect 278681 334464 278686 334520
rect 278742 334464 280140 334520
rect 278681 334462 280140 334464
rect 278681 334459 278747 334462
rect 583520 334236 584960 334476
rect 522941 333706 523007 333709
rect 519892 333704 523007 333706
rect 519892 333648 522946 333704
rect 523002 333648 523007 333704
rect 519892 333646 523007 333648
rect 522941 333643 523007 333646
rect 278681 332346 278747 332349
rect 278681 332344 280140 332346
rect 278681 332288 278686 332344
rect 278742 332288 280140 332344
rect 278681 332286 280140 332288
rect 278681 332283 278747 332286
rect 522573 331530 522639 331533
rect 519892 331528 522639 331530
rect 519892 331472 522578 331528
rect 522634 331472 522639 331528
rect 519892 331470 522639 331472
rect 522573 331467 522639 331470
rect 278681 330306 278747 330309
rect 278681 330304 280140 330306
rect 278681 330248 278686 330304
rect 278742 330248 280140 330304
rect 278681 330246 280140 330248
rect 278681 330243 278747 330246
rect 522941 329490 523007 329493
rect 519892 329488 523007 329490
rect 519892 329432 522946 329488
rect 523002 329432 523007 329488
rect 519892 329430 523007 329432
rect 522941 329427 523007 329430
rect 278681 328130 278747 328133
rect 278681 328128 280140 328130
rect 278681 328072 278686 328128
rect 278742 328072 280140 328128
rect 278681 328070 280140 328072
rect 278681 328067 278747 328070
rect 522941 327314 523007 327317
rect 519892 327312 523007 327314
rect 519892 327256 522946 327312
rect 523002 327256 523007 327312
rect 519892 327254 523007 327256
rect 522941 327251 523007 327254
rect 278037 325954 278103 325957
rect 278037 325952 280140 325954
rect 278037 325896 278042 325952
rect 278098 325896 280140 325952
rect 278037 325894 280140 325896
rect 278037 325891 278103 325894
rect 522941 325274 523007 325277
rect 519892 325272 523007 325274
rect 519892 325216 522946 325272
rect 523002 325216 523007 325272
rect 519892 325214 523007 325216
rect 522941 325211 523007 325214
rect 277669 323914 277735 323917
rect 277669 323912 280140 323914
rect 277669 323856 277674 323912
rect 277730 323856 280140 323912
rect 277669 323854 280140 323856
rect 277669 323851 277735 323854
rect -960 323098 480 323188
rect 3509 323098 3575 323101
rect 522297 323098 522363 323101
rect -960 323096 3575 323098
rect -960 323040 3514 323096
rect 3570 323040 3575 323096
rect -960 323038 3575 323040
rect 519892 323096 522363 323098
rect 519892 323040 522302 323096
rect 522358 323040 522363 323096
rect 519892 323038 522363 323040
rect -960 322948 480 323038
rect 3509 323035 3575 323038
rect 522297 323035 522363 323038
rect 580625 322690 580691 322693
rect 583520 322690 584960 322780
rect 580625 322688 584960 322690
rect 580625 322632 580630 322688
rect 580686 322632 584960 322688
rect 580625 322630 584960 322632
rect 580625 322627 580691 322630
rect 583520 322540 584960 322630
rect 278037 321738 278103 321741
rect 278037 321736 280140 321738
rect 278037 321680 278042 321736
rect 278098 321680 280140 321736
rect 278037 321678 280140 321680
rect 278037 321675 278103 321678
rect 522665 321058 522731 321061
rect 519892 321056 522731 321058
rect 519892 321000 522670 321056
rect 522726 321000 522731 321056
rect 519892 320998 522731 321000
rect 522665 320995 522731 320998
rect 278681 319562 278747 319565
rect 278681 319560 280140 319562
rect 278681 319504 278686 319560
rect 278742 319504 280140 319560
rect 278681 319502 280140 319504
rect 278681 319499 278747 319502
rect 522941 318882 523007 318885
rect 519892 318880 523007 318882
rect 519892 318824 522946 318880
rect 523002 318824 523007 318880
rect 519892 318822 523007 318824
rect 522941 318819 523007 318822
rect 278681 317522 278747 317525
rect 278681 317520 280140 317522
rect 278681 317464 278686 317520
rect 278742 317464 280140 317520
rect 278681 317462 280140 317464
rect 278681 317459 278747 317462
rect 522297 316842 522363 316845
rect 519892 316840 522363 316842
rect 519892 316784 522302 316840
rect 522358 316784 522363 316840
rect 519892 316782 522363 316784
rect 522297 316779 522363 316782
rect 278681 315346 278747 315349
rect 278681 315344 280140 315346
rect 278681 315288 278686 315344
rect 278742 315288 280140 315344
rect 278681 315286 280140 315288
rect 278681 315283 278747 315286
rect 522941 314666 523007 314669
rect 519892 314664 523007 314666
rect 519892 314608 522946 314664
rect 523002 314608 523007 314664
rect 519892 314606 523007 314608
rect 522941 314603 523007 314606
rect 278681 313306 278747 313309
rect 278681 313304 280140 313306
rect 278681 313248 278686 313304
rect 278742 313248 280140 313304
rect 278681 313246 280140 313248
rect 278681 313243 278747 313246
rect 522941 312626 523007 312629
rect 519892 312624 523007 312626
rect 519892 312568 522946 312624
rect 523002 312568 523007 312624
rect 519892 312566 523007 312568
rect 522941 312563 523007 312566
rect 278681 311130 278747 311133
rect 278681 311128 280140 311130
rect 278681 311072 278686 311128
rect 278742 311072 280140 311128
rect 278681 311070 280140 311072
rect 278681 311067 278747 311070
rect 580717 310858 580783 310861
rect 583520 310858 584960 310948
rect 580717 310856 584960 310858
rect 580717 310800 580722 310856
rect 580778 310800 584960 310856
rect 580717 310798 584960 310800
rect 580717 310795 580783 310798
rect 583520 310708 584960 310798
rect 522297 310450 522363 310453
rect 519892 310448 522363 310450
rect 519892 310392 522302 310448
rect 522358 310392 522363 310448
rect 519892 310390 522363 310392
rect 522297 310387 522363 310390
rect 277853 308954 277919 308957
rect 277853 308952 280140 308954
rect -960 308818 480 308908
rect 277853 308896 277858 308952
rect 277914 308896 280140 308952
rect 277853 308894 280140 308896
rect 277853 308891 277919 308894
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 522941 308410 523007 308413
rect 519892 308408 523007 308410
rect 519892 308352 522946 308408
rect 523002 308352 523007 308408
rect 519892 308350 523007 308352
rect 522941 308347 523007 308350
rect 278681 306914 278747 306917
rect 278681 306912 280140 306914
rect 278681 306856 278686 306912
rect 278742 306856 280140 306912
rect 278681 306854 280140 306856
rect 278681 306851 278747 306854
rect 522941 306234 523007 306237
rect 519892 306232 523007 306234
rect 519892 306176 522946 306232
rect 523002 306176 523007 306232
rect 519892 306174 523007 306176
rect 522941 306171 523007 306174
rect 278681 304738 278747 304741
rect 278681 304736 280140 304738
rect 278681 304680 278686 304736
rect 278742 304680 280140 304736
rect 278681 304678 280140 304680
rect 278681 304675 278747 304678
rect 522297 304194 522363 304197
rect 519892 304192 522363 304194
rect 519892 304136 522302 304192
rect 522358 304136 522363 304192
rect 519892 304134 522363 304136
rect 522297 304131 522363 304134
rect 278681 302562 278747 302565
rect 278681 302560 280140 302562
rect 278681 302504 278686 302560
rect 278742 302504 280140 302560
rect 278681 302502 280140 302504
rect 278681 302499 278747 302502
rect 522941 302018 523007 302021
rect 519892 302016 523007 302018
rect 519892 301960 522946 302016
rect 523002 301960 523007 302016
rect 519892 301958 523007 301960
rect 522941 301955 523007 301958
rect 278681 300522 278747 300525
rect 278681 300520 280140 300522
rect 278681 300464 278686 300520
rect 278742 300464 280140 300520
rect 278681 300462 280140 300464
rect 278681 300459 278747 300462
rect 522941 299978 523007 299981
rect 519892 299976 523007 299978
rect 519892 299920 522946 299976
rect 523002 299920 523007 299976
rect 519892 299918 523007 299920
rect 522941 299915 523007 299918
rect 579981 299162 580047 299165
rect 583520 299162 584960 299252
rect 579981 299160 584960 299162
rect 579981 299104 579986 299160
rect 580042 299104 584960 299160
rect 579981 299102 584960 299104
rect 579981 299099 580047 299102
rect 583520 299012 584960 299102
rect 278681 298346 278747 298349
rect 278681 298344 280140 298346
rect 278681 298288 278686 298344
rect 278742 298288 280140 298344
rect 278681 298286 280140 298288
rect 278681 298283 278747 298286
rect 522941 297938 523007 297941
rect 519892 297936 523007 297938
rect 519892 297880 522946 297936
rect 523002 297880 523007 297936
rect 519892 297878 523007 297880
rect 522941 297875 523007 297878
rect 278681 296306 278747 296309
rect 278681 296304 280140 296306
rect 278681 296248 278686 296304
rect 278742 296248 280140 296304
rect 278681 296246 280140 296248
rect 278681 296243 278747 296246
rect 522941 295762 523007 295765
rect 519892 295760 523007 295762
rect 519892 295704 522946 295760
rect 523002 295704 523007 295760
rect 519892 295702 523007 295704
rect 522941 295699 523007 295702
rect -960 294402 480 294492
rect 3049 294402 3115 294405
rect -960 294400 3115 294402
rect -960 294344 3054 294400
rect 3110 294344 3115 294400
rect -960 294342 3115 294344
rect -960 294252 480 294342
rect 3049 294339 3115 294342
rect 278681 294130 278747 294133
rect 278681 294128 280140 294130
rect 278681 294072 278686 294128
rect 278742 294072 280140 294128
rect 278681 294070 280140 294072
rect 278681 294067 278747 294070
rect 522941 293722 523007 293725
rect 519892 293720 523007 293722
rect 519892 293664 522946 293720
rect 523002 293664 523007 293720
rect 519892 293662 523007 293664
rect 522941 293659 523007 293662
rect 278681 291954 278747 291957
rect 278681 291952 280140 291954
rect 278681 291896 278686 291952
rect 278742 291896 280140 291952
rect 278681 291894 280140 291896
rect 278681 291891 278747 291894
rect 522573 291546 522639 291549
rect 519892 291544 522639 291546
rect 519892 291488 522578 291544
rect 522634 291488 522639 291544
rect 519892 291486 522639 291488
rect 522573 291483 522639 291486
rect 278681 289914 278747 289917
rect 278681 289912 280140 289914
rect 278681 289856 278686 289912
rect 278742 289856 280140 289912
rect 278681 289854 280140 289856
rect 278681 289851 278747 289854
rect 522941 289506 523007 289509
rect 519892 289504 523007 289506
rect 519892 289448 522946 289504
rect 523002 289448 523007 289504
rect 519892 289446 523007 289448
rect 522941 289443 523007 289446
rect 278681 287738 278747 287741
rect 278681 287736 280140 287738
rect 278681 287680 278686 287736
rect 278742 287680 280140 287736
rect 278681 287678 280140 287680
rect 278681 287675 278747 287678
rect 522573 287330 522639 287333
rect 519892 287328 522639 287330
rect 519892 287272 522578 287328
rect 522634 287272 522639 287328
rect 583520 287316 584960 287556
rect 519892 287270 522639 287272
rect 522573 287267 522639 287270
rect 278681 285698 278747 285701
rect 278681 285696 280140 285698
rect 278681 285640 278686 285696
rect 278742 285640 280140 285696
rect 278681 285638 280140 285640
rect 278681 285635 278747 285638
rect 522573 285290 522639 285293
rect 519892 285288 522639 285290
rect 519892 285232 522578 285288
rect 522634 285232 522639 285288
rect 519892 285230 522639 285232
rect 522573 285227 522639 285230
rect 278681 283522 278747 283525
rect 278681 283520 280140 283522
rect 278681 283464 278686 283520
rect 278742 283464 280140 283520
rect 278681 283462 280140 283464
rect 278681 283459 278747 283462
rect 522481 283114 522547 283117
rect 519892 283112 522547 283114
rect 519892 283056 522486 283112
rect 522542 283056 522547 283112
rect 519892 283054 522547 283056
rect 522481 283051 522547 283054
rect 277853 281346 277919 281349
rect 277853 281344 280140 281346
rect 277853 281288 277858 281344
rect 277914 281288 280140 281344
rect 277853 281286 280140 281288
rect 277853 281283 277919 281286
rect 522941 281074 523007 281077
rect 519892 281072 523007 281074
rect 519892 281016 522946 281072
rect 523002 281016 523007 281072
rect 519892 281014 523007 281016
rect 522941 281011 523007 281014
rect -960 280122 480 280212
rect 3509 280122 3575 280125
rect -960 280120 3575 280122
rect -960 280064 3514 280120
rect 3570 280064 3575 280120
rect -960 280062 3575 280064
rect -960 279972 480 280062
rect 3509 280059 3575 280062
rect 278681 279306 278747 279309
rect 278681 279304 280140 279306
rect 278681 279248 278686 279304
rect 278742 279248 280140 279304
rect 278681 279246 280140 279248
rect 278681 279243 278747 279246
rect 522297 278898 522363 278901
rect 519892 278896 522363 278898
rect 519892 278840 522302 278896
rect 522358 278840 522363 278896
rect 519892 278838 522363 278840
rect 522297 278835 522363 278838
rect 278681 277130 278747 277133
rect 278681 277128 280140 277130
rect 278681 277072 278686 277128
rect 278742 277072 280140 277128
rect 278681 277070 280140 277072
rect 278681 277067 278747 277070
rect 522481 276858 522547 276861
rect 519892 276856 522547 276858
rect 519892 276800 522486 276856
rect 522542 276800 522547 276856
rect 519892 276798 522547 276800
rect 522481 276795 522547 276798
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 278037 274954 278103 274957
rect 278037 274952 280140 274954
rect 278037 274896 278042 274952
rect 278098 274896 280140 274952
rect 278037 274894 280140 274896
rect 278037 274891 278103 274894
rect 522941 274682 523007 274685
rect 519892 274680 523007 274682
rect 519892 274624 522946 274680
rect 523002 274624 523007 274680
rect 519892 274622 523007 274624
rect 522941 274619 523007 274622
rect 278681 272914 278747 272917
rect 278681 272912 280140 272914
rect 278681 272856 278686 272912
rect 278742 272856 280140 272912
rect 278681 272854 280140 272856
rect 278681 272851 278747 272854
rect 522297 272642 522363 272645
rect 519892 272640 522363 272642
rect 519892 272584 522302 272640
rect 522358 272584 522363 272640
rect 519892 272582 522363 272584
rect 522297 272579 522363 272582
rect 278681 270738 278747 270741
rect 278681 270736 280140 270738
rect 278681 270680 278686 270736
rect 278742 270680 280140 270736
rect 278681 270678 280140 270680
rect 278681 270675 278747 270678
rect 522849 270466 522915 270469
rect 519892 270464 522915 270466
rect 519892 270408 522854 270464
rect 522910 270408 522915 270464
rect 519892 270406 522915 270408
rect 522849 270403 522915 270406
rect 278681 268698 278747 268701
rect 278681 268696 280140 268698
rect 278681 268640 278686 268696
rect 278742 268640 280140 268696
rect 278681 268638 280140 268640
rect 278681 268635 278747 268638
rect 522941 268426 523007 268429
rect 519892 268424 523007 268426
rect 519892 268368 522946 268424
rect 523002 268368 523007 268424
rect 519892 268366 523007 268368
rect 522941 268363 523007 268366
rect 278037 266522 278103 266525
rect 278037 266520 280140 266522
rect 278037 266464 278042 266520
rect 278098 266464 280140 266520
rect 278037 266462 280140 266464
rect 278037 266459 278103 266462
rect 522573 266250 522639 266253
rect 519892 266248 522639 266250
rect 519892 266192 522578 266248
rect 522634 266192 522639 266248
rect 519892 266190 522639 266192
rect 522573 266187 522639 266190
rect -960 265706 480 265796
rect 3509 265706 3575 265709
rect -960 265704 3575 265706
rect -960 265648 3514 265704
rect 3570 265648 3575 265704
rect -960 265646 3575 265648
rect -960 265556 480 265646
rect 3509 265643 3575 265646
rect 278681 264346 278747 264349
rect 278681 264344 280140 264346
rect 278681 264288 278686 264344
rect 278742 264288 280140 264344
rect 278681 264286 280140 264288
rect 278681 264283 278747 264286
rect 522757 264210 522823 264213
rect 519892 264208 522823 264210
rect 519892 264152 522762 264208
rect 522818 264152 522823 264208
rect 519892 264150 522823 264152
rect 522757 264147 522823 264150
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 278681 262306 278747 262309
rect 278681 262304 280140 262306
rect 278681 262248 278686 262304
rect 278742 262248 280140 262304
rect 278681 262246 280140 262248
rect 278681 262243 278747 262246
rect 522573 262034 522639 262037
rect 519892 262032 522639 262034
rect 519892 261976 522578 262032
rect 522634 261976 522639 262032
rect 519892 261974 522639 261976
rect 522573 261971 522639 261974
rect 278313 260130 278379 260133
rect 278313 260128 280140 260130
rect 278313 260072 278318 260128
rect 278374 260072 280140 260128
rect 278313 260070 280140 260072
rect 278313 260067 278379 260070
rect 522573 259994 522639 259997
rect 519892 259992 522639 259994
rect 519892 259936 522578 259992
rect 522634 259936 522639 259992
rect 519892 259934 522639 259936
rect 522573 259931 522639 259934
rect 277853 257954 277919 257957
rect 277853 257952 280140 257954
rect 277853 257896 277858 257952
rect 277914 257896 280140 257952
rect 277853 257894 280140 257896
rect 277853 257891 277919 257894
rect 522573 257818 522639 257821
rect 519892 257816 522639 257818
rect 519892 257760 522578 257816
rect 522634 257760 522639 257816
rect 519892 257758 522639 257760
rect 522573 257755 522639 257758
rect 278681 255914 278747 255917
rect 278681 255912 280140 255914
rect 278681 255856 278686 255912
rect 278742 255856 280140 255912
rect 278681 255854 280140 255856
rect 278681 255851 278747 255854
rect 522665 255778 522731 255781
rect 519892 255776 522731 255778
rect 519892 255720 522670 255776
rect 522726 255720 522731 255776
rect 519892 255718 522731 255720
rect 522665 255715 522731 255718
rect 277853 253738 277919 253741
rect 277853 253736 280140 253738
rect 277853 253680 277858 253736
rect 277914 253680 280140 253736
rect 277853 253678 280140 253680
rect 277853 253675 277919 253678
rect 523677 253602 523743 253605
rect 519892 253600 523743 253602
rect 519892 253544 523682 253600
rect 523738 253544 523743 253600
rect 519892 253542 523743 253544
rect 523677 253539 523743 253542
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect 278681 251698 278747 251701
rect 278681 251696 280140 251698
rect 278681 251640 278686 251696
rect 278742 251640 280140 251696
rect 278681 251638 280140 251640
rect 278681 251635 278747 251638
rect 522481 251562 522547 251565
rect 519892 251560 522547 251562
rect 519892 251504 522486 251560
rect 522542 251504 522547 251560
rect 519892 251502 522547 251504
rect 522481 251499 522547 251502
rect -960 251290 480 251380
rect 3601 251290 3667 251293
rect -960 251288 3667 251290
rect -960 251232 3606 251288
rect 3662 251232 3667 251288
rect -960 251230 3667 251232
rect -960 251140 480 251230
rect 3601 251227 3667 251230
rect 278681 249522 278747 249525
rect 278681 249520 280140 249522
rect 278681 249464 278686 249520
rect 278742 249464 280140 249520
rect 278681 249462 280140 249464
rect 278681 249459 278747 249462
rect 522297 249386 522363 249389
rect 519892 249384 522363 249386
rect 519892 249328 522302 249384
rect 522358 249328 522363 249384
rect 519892 249326 522363 249328
rect 522297 249323 522363 249326
rect 278037 247346 278103 247349
rect 522297 247346 522363 247349
rect 278037 247344 280140 247346
rect 278037 247288 278042 247344
rect 278098 247288 280140 247344
rect 278037 247286 280140 247288
rect 519892 247344 522363 247346
rect 519892 247288 522302 247344
rect 522358 247288 522363 247344
rect 519892 247286 522363 247288
rect 278037 247283 278103 247286
rect 522297 247283 522363 247286
rect 278129 245306 278195 245309
rect 278129 245304 280140 245306
rect 278129 245248 278134 245304
rect 278190 245248 280140 245304
rect 278129 245246 280140 245248
rect 278129 245243 278195 245246
rect 522297 245170 522363 245173
rect 519892 245168 522363 245170
rect 519892 245112 522302 245168
rect 522358 245112 522363 245168
rect 519892 245110 522363 245112
rect 522297 245107 522363 245110
rect 277393 243130 277459 243133
rect 522389 243130 522455 243133
rect 277393 243128 280140 243130
rect 277393 243072 277398 243128
rect 277454 243072 280140 243128
rect 277393 243070 280140 243072
rect 519892 243128 522455 243130
rect 519892 243072 522394 243128
rect 522450 243072 522455 243128
rect 519892 243070 522455 243072
rect 277393 243067 277459 243070
rect 522389 243067 522455 243070
rect 278681 241090 278747 241093
rect 278681 241088 280140 241090
rect 278681 241032 278686 241088
rect 278742 241060 280140 241088
rect 278742 241032 280170 241060
rect 278681 241030 280170 241032
rect 278681 241027 278747 241030
rect 280110 240821 280170 241030
rect 280110 240816 280219 240821
rect 280110 240760 280158 240816
rect 280214 240760 280219 240816
rect 280110 240758 280219 240760
rect 280153 240755 280219 240758
rect 316033 240682 316099 240685
rect 325601 240682 325667 240685
rect 316033 240680 325667 240682
rect 316033 240624 316038 240680
rect 316094 240624 325606 240680
rect 325662 240624 325667 240680
rect 316033 240622 325667 240624
rect 316033 240619 316099 240622
rect 325601 240619 325667 240622
rect 357433 240682 357499 240685
rect 360377 240682 360443 240685
rect 357433 240680 360443 240682
rect 357433 240624 357438 240680
rect 357494 240624 360382 240680
rect 360438 240624 360443 240680
rect 357433 240622 360443 240624
rect 357433 240619 357499 240622
rect 360377 240619 360443 240622
rect 519862 240546 519922 241060
rect 522389 240546 522455 240549
rect 519862 240544 522455 240546
rect 519862 240488 522394 240544
rect 522450 240488 522455 240544
rect 519862 240486 522455 240488
rect 522389 240483 522455 240486
rect 583520 240396 584960 240636
rect 522113 237146 522179 237149
rect 522798 237146 522804 237148
rect 522113 237144 522804 237146
rect -960 237010 480 237100
rect 522113 237088 522118 237144
rect 522174 237088 522804 237144
rect 522113 237086 522804 237088
rect 522113 237083 522179 237086
rect 522798 237084 522804 237086
rect 522868 237084 522874 237148
rect 3509 237010 3575 237013
rect -960 237008 3575 237010
rect -960 236952 3514 237008
rect 3570 236952 3575 237008
rect -960 236950 3575 236952
rect -960 236860 480 236950
rect 3509 236947 3575 236950
rect 431769 231842 431835 231845
rect 431953 231842 432019 231845
rect 431769 231840 432019 231842
rect 431769 231784 431774 231840
rect 431830 231784 431958 231840
rect 432014 231784 432019 231840
rect 431769 231782 432019 231784
rect 431769 231779 431835 231782
rect 431953 231779 432019 231782
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 336406 220764 336412 220828
rect 336476 220826 336482 220828
rect 336641 220826 336707 220829
rect 336476 220824 336707 220826
rect 336476 220768 336646 220824
rect 336702 220768 336707 220824
rect 336476 220766 336707 220768
rect 336476 220764 336482 220766
rect 336641 220763 336707 220766
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 329373 212532 329439 212533
rect 329373 212530 329420 212532
rect 329328 212528 329420 212530
rect 329328 212472 329378 212528
rect 329328 212470 329420 212472
rect 329373 212468 329420 212470
rect 329484 212468 329490 212532
rect 329373 212467 329439 212468
rect -960 208178 480 208268
rect 3509 208178 3575 208181
rect -960 208176 3575 208178
rect -960 208120 3514 208176
rect 3570 208120 3575 208176
rect -960 208118 3575 208120
rect -960 208028 480 208118
rect 3509 208115 3575 208118
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 347773 204232 347839 204237
rect 347773 204176 347778 204232
rect 347834 204176 347839 204232
rect 347773 204171 347839 204176
rect 357341 204234 357407 204237
rect 362861 204234 362927 204237
rect 367093 204234 367159 204237
rect 357341 204232 357818 204234
rect 357341 204176 357346 204232
rect 357402 204176 357818 204232
rect 357341 204174 357818 204176
rect 357341 204171 357407 204174
rect 292481 204098 292547 204101
rect 347776 204098 347836 204171
rect 292481 204096 347836 204098
rect 292481 204040 292486 204096
rect 292542 204040 347836 204096
rect 292481 204038 347836 204040
rect 292481 204035 292547 204038
rect 288341 203962 288407 203965
rect 355317 203962 355383 203965
rect 357433 203964 357499 203965
rect 288341 203960 355383 203962
rect 288341 203904 288346 203960
rect 288402 203904 355322 203960
rect 355378 203904 355383 203960
rect 288341 203902 355383 203904
rect 288341 203899 288407 203902
rect 355317 203899 355383 203902
rect 357382 203900 357388 203964
rect 357452 203962 357499 203964
rect 357758 203962 357818 204174
rect 362861 204232 367159 204234
rect 362861 204176 362866 204232
rect 362922 204176 367098 204232
rect 367154 204176 367159 204232
rect 362861 204174 367159 204176
rect 362861 204171 362927 204174
rect 367093 204171 367159 204174
rect 448278 204172 448284 204236
rect 448348 204234 448354 204236
rect 448421 204234 448487 204237
rect 448348 204232 448487 204234
rect 448348 204176 448426 204232
rect 448482 204176 448487 204232
rect 448348 204174 448487 204176
rect 448348 204172 448354 204174
rect 448421 204171 448487 204174
rect 449382 204172 449388 204236
rect 449452 204234 449458 204236
rect 449801 204234 449867 204237
rect 449452 204232 449867 204234
rect 449452 204176 449806 204232
rect 449862 204176 449867 204232
rect 449452 204174 449867 204176
rect 449452 204172 449458 204174
rect 449801 204171 449867 204174
rect 451774 204172 451780 204236
rect 451844 204234 451850 204236
rect 452561 204234 452627 204237
rect 453297 204236 453363 204237
rect 453246 204234 453252 204236
rect 451844 204232 452627 204234
rect 451844 204176 452566 204232
rect 452622 204176 452627 204232
rect 451844 204174 452627 204176
rect 453206 204174 453252 204234
rect 453316 204232 453363 204236
rect 453358 204176 453363 204232
rect 451844 204172 451850 204174
rect 452561 204171 452627 204174
rect 453246 204172 453252 204174
rect 453316 204172 453363 204176
rect 454166 204172 454172 204236
rect 454236 204234 454242 204236
rect 455137 204234 455203 204237
rect 454236 204232 455203 204234
rect 454236 204176 455142 204232
rect 455198 204176 455203 204232
rect 454236 204174 455203 204176
rect 454236 204172 454242 204174
rect 453297 204171 453363 204172
rect 455137 204171 455203 204174
rect 456374 204172 456380 204236
rect 456444 204234 456450 204236
rect 456701 204234 456767 204237
rect 456444 204232 456767 204234
rect 456444 204176 456706 204232
rect 456762 204176 456767 204232
rect 456444 204174 456767 204176
rect 456444 204172 456450 204174
rect 456701 204171 456767 204174
rect 468150 204172 468156 204236
rect 468220 204234 468226 204236
rect 469121 204234 469187 204237
rect 468220 204232 469187 204234
rect 468220 204176 469126 204232
rect 469182 204176 469187 204232
rect 468220 204174 469187 204176
rect 468220 204172 468226 204174
rect 469121 204171 469187 204174
rect 470358 204172 470364 204236
rect 470428 204234 470434 204236
rect 470501 204234 470567 204237
rect 484393 204236 484459 204237
rect 470428 204232 470567 204234
rect 470428 204176 470506 204232
rect 470562 204176 470567 204232
rect 470428 204174 470567 204176
rect 470428 204172 470434 204174
rect 470501 204171 470567 204174
rect 484342 204172 484348 204236
rect 484412 204234 484459 204236
rect 484412 204232 484504 204234
rect 484454 204176 484504 204232
rect 484412 204174 484504 204176
rect 484412 204172 484459 204174
rect 484393 204171 484459 204172
rect 449157 204098 449223 204101
rect 450905 204100 450971 204101
rect 449566 204098 449572 204100
rect 449157 204096 449572 204098
rect 449157 204040 449162 204096
rect 449218 204040 449572 204096
rect 449157 204038 449572 204040
rect 449157 204035 449223 204038
rect 449566 204036 449572 204038
rect 449636 204036 449642 204100
rect 450854 204036 450860 204100
rect 450924 204098 450971 204100
rect 452009 204098 452075 204101
rect 452142 204098 452148 204100
rect 450924 204096 451016 204098
rect 450966 204040 451016 204096
rect 450924 204038 451016 204040
rect 452009 204096 452148 204098
rect 452009 204040 452014 204096
rect 452070 204040 452148 204096
rect 452009 204038 452148 204040
rect 450924 204036 450971 204038
rect 450905 204035 450971 204036
rect 452009 204035 452075 204038
rect 452142 204036 452148 204038
rect 452212 204036 452218 204100
rect 454534 204036 454540 204100
rect 454604 204098 454610 204100
rect 454677 204098 454743 204101
rect 454604 204096 454743 204098
rect 454604 204040 454682 204096
rect 454738 204040 454743 204096
rect 454604 204038 454743 204040
rect 454604 204036 454610 204038
rect 454677 204035 454743 204038
rect 456057 204098 456123 204101
rect 456558 204098 456564 204100
rect 456057 204096 456564 204098
rect 456057 204040 456062 204096
rect 456118 204040 456564 204096
rect 456057 204038 456564 204040
rect 456057 204035 456123 204038
rect 456558 204036 456564 204038
rect 456628 204036 456634 204100
rect 464470 204036 464476 204100
rect 464540 204098 464546 204100
rect 464981 204098 465047 204101
rect 464540 204096 465047 204098
rect 464540 204040 464986 204096
rect 465042 204040 465047 204096
rect 464540 204038 465047 204040
rect 464540 204036 464546 204038
rect 464981 204035 465047 204038
rect 465758 204036 465764 204100
rect 465828 204098 465834 204100
rect 466269 204098 466335 204101
rect 465828 204096 466335 204098
rect 465828 204040 466274 204096
rect 466330 204040 466335 204096
rect 465828 204038 466335 204040
rect 465828 204036 465834 204038
rect 466269 204035 466335 204038
rect 469254 204036 469260 204100
rect 469324 204098 469330 204100
rect 470409 204098 470475 204101
rect 469324 204096 470475 204098
rect 469324 204040 470414 204096
rect 470470 204040 470475 204096
rect 469324 204038 470475 204040
rect 469324 204036 469330 204038
rect 470409 204035 470475 204038
rect 475653 204098 475719 204101
rect 477493 204100 477559 204101
rect 476062 204098 476068 204100
rect 475653 204096 476068 204098
rect 475653 204040 475658 204096
rect 475714 204040 476068 204096
rect 475653 204038 476068 204040
rect 475653 204035 475719 204038
rect 476062 204036 476068 204038
rect 476132 204036 476138 204100
rect 477493 204098 477540 204100
rect 477448 204096 477540 204098
rect 477448 204040 477498 204096
rect 477448 204038 477540 204040
rect 477493 204036 477540 204038
rect 477604 204036 477610 204100
rect 483013 204098 483079 204101
rect 483422 204098 483428 204100
rect 483013 204096 483428 204098
rect 483013 204040 483018 204096
rect 483074 204040 483428 204096
rect 483013 204038 483428 204040
rect 477493 204035 477559 204036
rect 483013 204035 483079 204038
rect 483422 204036 483428 204038
rect 483492 204036 483498 204100
rect 485773 204098 485839 204101
rect 486366 204098 486372 204100
rect 485773 204096 486372 204098
rect 485773 204040 485778 204096
rect 485834 204040 486372 204096
rect 485773 204038 486372 204040
rect 485773 204035 485839 204038
rect 486366 204036 486372 204038
rect 486436 204036 486442 204100
rect 360510 203962 360516 203964
rect 357452 203960 357544 203962
rect 357494 203904 357544 203960
rect 357452 203902 357544 203904
rect 357758 203902 360516 203962
rect 357452 203900 357499 203902
rect 360510 203900 360516 203902
rect 360580 203900 360586 203964
rect 437473 203962 437539 203965
rect 451089 203962 451155 203965
rect 437473 203960 451155 203962
rect 437473 203904 437478 203960
rect 437534 203904 451094 203960
rect 451150 203904 451155 203960
rect 437473 203902 451155 203904
rect 357433 203899 357499 203900
rect 437473 203899 437539 203902
rect 451089 203899 451155 203902
rect 457478 203900 457484 203964
rect 457548 203962 457554 203964
rect 457989 203962 458055 203965
rect 457548 203960 458055 203962
rect 457548 203904 457994 203960
rect 458050 203904 458055 203960
rect 457548 203902 458055 203904
rect 457548 203900 457554 203902
rect 457989 203899 458055 203902
rect 460054 203900 460060 203964
rect 460124 203962 460130 203964
rect 460841 203962 460907 203965
rect 460124 203960 460907 203962
rect 460124 203904 460846 203960
rect 460902 203904 460907 203960
rect 460124 203902 460907 203904
rect 460124 203900 460130 203902
rect 460841 203899 460907 203902
rect 461577 203962 461643 203965
rect 466361 203962 466427 203965
rect 461577 203960 466427 203962
rect 461577 203904 461582 203960
rect 461638 203904 466366 203960
rect 466422 203904 466427 203960
rect 461577 203902 466427 203904
rect 461577 203899 461643 203902
rect 466361 203899 466427 203902
rect 471237 203962 471303 203965
rect 480161 203962 480227 203965
rect 490189 203964 490255 203965
rect 490189 203962 490236 203964
rect 471237 203960 480227 203962
rect 471237 203904 471242 203960
rect 471298 203904 480166 203960
rect 480222 203904 480227 203960
rect 471237 203902 480227 203904
rect 490144 203960 490236 203962
rect 490144 203904 490194 203960
rect 490144 203902 490236 203904
rect 471237 203899 471303 203902
rect 480161 203899 480227 203902
rect 490189 203900 490236 203902
rect 490300 203900 490306 203964
rect 490189 203899 490255 203900
rect 289721 203826 289787 203829
rect 361614 203826 361620 203828
rect 289721 203824 361620 203826
rect 289721 203768 289726 203824
rect 289782 203768 361620 203824
rect 289721 203766 361620 203768
rect 289721 203763 289787 203766
rect 361614 203764 361620 203766
rect 361684 203764 361690 203828
rect 376569 203826 376635 203829
rect 442257 203826 442323 203829
rect 376569 203824 442323 203826
rect 376569 203768 376574 203824
rect 376630 203768 442262 203824
rect 442318 203768 442323 203824
rect 376569 203766 442323 203768
rect 376569 203763 376635 203766
rect 442257 203763 442323 203766
rect 451089 203826 451155 203829
rect 485814 203826 485820 203828
rect 451089 203824 485820 203826
rect 451089 203768 451094 203824
rect 451150 203768 485820 203824
rect 451089 203766 485820 203768
rect 451089 203763 451155 203766
rect 485814 203764 485820 203766
rect 485884 203764 485890 203828
rect 330937 203692 331003 203693
rect 330886 203628 330892 203692
rect 330956 203690 331003 203692
rect 340965 203692 341031 203693
rect 340965 203690 341012 203692
rect 330956 203688 331048 203690
rect 330998 203632 331048 203688
rect 330956 203630 331048 203632
rect 340920 203688 341012 203690
rect 340920 203632 340970 203688
rect 340920 203630 341012 203632
rect 330956 203628 331003 203630
rect 330937 203627 331003 203628
rect 340965 203628 341012 203630
rect 341076 203628 341082 203692
rect 342253 203690 342319 203693
rect 347773 203692 347839 203693
rect 349153 203692 349219 203693
rect 342846 203690 342852 203692
rect 342253 203688 342852 203690
rect 342253 203632 342258 203688
rect 342314 203632 342852 203688
rect 342253 203630 342852 203632
rect 340965 203627 341031 203628
rect 342253 203627 342319 203630
rect 342846 203628 342852 203630
rect 342916 203628 342922 203692
rect 347773 203690 347820 203692
rect 347728 203688 347820 203690
rect 347728 203632 347778 203688
rect 347728 203630 347820 203632
rect 347773 203628 347820 203630
rect 347884 203628 347890 203692
rect 349102 203628 349108 203692
rect 349172 203690 349219 203692
rect 351913 203690 351979 203693
rect 352782 203690 352788 203692
rect 349172 203688 349264 203690
rect 349214 203632 349264 203688
rect 349172 203630 349264 203632
rect 351913 203688 352788 203690
rect 351913 203632 351918 203688
rect 351974 203632 352788 203688
rect 351913 203630 352788 203632
rect 349172 203628 349219 203630
rect 347773 203627 347839 203628
rect 349153 203627 349219 203628
rect 351913 203627 351979 203630
rect 352782 203628 352788 203630
rect 352852 203628 352858 203692
rect 358721 203690 358787 203693
rect 376385 203690 376451 203693
rect 358721 203688 376451 203690
rect 358721 203632 358726 203688
rect 358782 203632 376390 203688
rect 376446 203632 376451 203688
rect 358721 203630 376451 203632
rect 358721 203627 358787 203630
rect 376385 203627 376451 203630
rect 376569 203690 376635 203693
rect 437473 203690 437539 203693
rect 376569 203688 437539 203690
rect 376569 203632 376574 203688
rect 376630 203632 437478 203688
rect 437534 203632 437539 203688
rect 376569 203630 437539 203632
rect 376569 203627 376635 203630
rect 437473 203627 437539 203630
rect 451181 203690 451247 203693
rect 487470 203690 487476 203692
rect 451181 203688 487476 203690
rect 451181 203632 451186 203688
rect 451242 203632 487476 203688
rect 451181 203630 487476 203632
rect 451181 203627 451247 203630
rect 487470 203628 487476 203630
rect 487540 203628 487546 203692
rect 340045 203556 340111 203557
rect 342253 203556 342319 203557
rect 343633 203556 343699 203557
rect 340045 203552 340092 203556
rect 340156 203554 340162 203556
rect 342253 203554 342300 203556
rect 340045 203496 340050 203552
rect 340045 203492 340092 203496
rect 340156 203494 340202 203554
rect 342208 203552 342300 203554
rect 342208 203496 342258 203552
rect 342208 203494 342300 203496
rect 340156 203492 340162 203494
rect 342253 203492 342300 203494
rect 342364 203492 342370 203556
rect 343582 203554 343588 203556
rect 343542 203494 343588 203554
rect 343652 203552 343699 203556
rect 343694 203496 343699 203552
rect 343582 203492 343588 203494
rect 343652 203492 343699 203496
rect 340045 203491 340111 203492
rect 342253 203491 342319 203492
rect 343633 203491 343699 203492
rect 354673 203554 354739 203557
rect 354806 203554 354812 203556
rect 354673 203552 354812 203554
rect 354673 203496 354678 203552
rect 354734 203496 354812 203552
rect 354673 203494 354812 203496
rect 354673 203491 354739 203494
rect 354806 203492 354812 203494
rect 354876 203492 354882 203556
rect 355961 203554 356027 203557
rect 360193 203554 360259 203557
rect 466361 203554 466427 203557
rect 471237 203554 471303 203557
rect 355961 203552 360259 203554
rect 355961 203496 355966 203552
rect 356022 203496 360198 203552
rect 360254 203496 360259 203552
rect 355961 203494 360259 203496
rect 355961 203491 356027 203494
rect 360193 203491 360259 203494
rect 399526 203494 427922 203554
rect 329598 203356 329604 203420
rect 329668 203418 329674 203420
rect 329741 203418 329807 203421
rect 329668 203416 329807 203418
rect 329668 203360 329746 203416
rect 329802 203360 329807 203416
rect 329668 203358 329807 203360
rect 329668 203356 329674 203358
rect 329741 203355 329807 203358
rect 330702 203356 330708 203420
rect 330772 203418 330778 203420
rect 331121 203418 331187 203421
rect 330772 203416 331187 203418
rect 330772 203360 331126 203416
rect 331182 203360 331187 203416
rect 330772 203358 331187 203360
rect 330772 203356 330778 203358
rect 331121 203355 331187 203358
rect 334198 203356 334204 203420
rect 334268 203418 334274 203420
rect 335169 203418 335235 203421
rect 334268 203416 335235 203418
rect 334268 203360 335174 203416
rect 335230 203360 335235 203416
rect 334268 203358 335235 203360
rect 334268 203356 334274 203358
rect 335169 203355 335235 203358
rect 336733 203418 336799 203421
rect 336958 203418 336964 203420
rect 336733 203416 336964 203418
rect 336733 203360 336738 203416
rect 336794 203360 336964 203416
rect 336733 203358 336964 203360
rect 336733 203355 336799 203358
rect 336958 203356 336964 203358
rect 337028 203356 337034 203420
rect 341701 203418 341767 203421
rect 342478 203418 342484 203420
rect 341701 203416 342484 203418
rect 341701 203360 341706 203416
rect 341762 203360 342484 203416
rect 341701 203358 342484 203360
rect 341701 203355 341767 203358
rect 342478 203356 342484 203358
rect 342548 203418 342554 203420
rect 345565 203418 345631 203421
rect 342548 203416 345631 203418
rect 342548 203360 345570 203416
rect 345626 203360 345631 203416
rect 342548 203358 345631 203360
rect 342548 203356 342554 203358
rect 345565 203355 345631 203358
rect 355317 203418 355383 203421
rect 364333 203420 364399 203421
rect 362902 203418 362908 203420
rect 355317 203416 362908 203418
rect 355317 203360 355322 203416
rect 355378 203360 362908 203416
rect 355317 203358 362908 203360
rect 355317 203355 355383 203358
rect 362902 203356 362908 203358
rect 362972 203356 362978 203420
rect 364333 203418 364380 203420
rect 364288 203416 364380 203418
rect 364288 203360 364338 203416
rect 364288 203358 364380 203360
rect 364333 203356 364380 203358
rect 364444 203356 364450 203420
rect 366817 203418 366883 203421
rect 367502 203418 367508 203420
rect 366817 203416 367508 203418
rect 366817 203360 366822 203416
rect 366878 203360 367508 203416
rect 366817 203358 367508 203360
rect 364333 203355 364399 203356
rect 366817 203355 366883 203358
rect 367502 203356 367508 203358
rect 367572 203356 367578 203420
rect 399526 203418 399586 203494
rect 385174 203358 399586 203418
rect 427862 203418 427922 203494
rect 466361 203552 471303 203554
rect 466361 203496 466366 203552
rect 466422 203496 471242 203552
rect 471298 203496 471303 203552
rect 466361 203494 471303 203496
rect 466361 203491 466427 203494
rect 471237 203491 471303 203494
rect 473905 203554 473971 203557
rect 474222 203554 474228 203556
rect 473905 203552 474228 203554
rect 473905 203496 473910 203552
rect 473966 203496 474228 203552
rect 473905 203494 474228 203496
rect 473905 203491 473971 203494
rect 474222 203492 474228 203494
rect 474292 203554 474298 203556
rect 474457 203554 474523 203557
rect 474292 203552 474523 203554
rect 474292 203496 474462 203552
rect 474518 203496 474523 203552
rect 474292 203494 474523 203496
rect 474292 203492 474298 203494
rect 474457 203491 474523 203494
rect 480161 203554 480227 203557
rect 480621 203556 480687 203557
rect 480621 203554 480668 203556
rect 480161 203552 480362 203554
rect 480161 203496 480166 203552
rect 480222 203496 480362 203552
rect 480161 203494 480362 203496
rect 480576 203552 480668 203554
rect 480576 203496 480626 203552
rect 480576 203494 480668 203496
rect 480161 203491 480227 203494
rect 427862 203358 455890 203418
rect 328126 203220 328132 203284
rect 328196 203282 328202 203284
rect 328361 203282 328427 203285
rect 328196 203280 328427 203282
rect 328196 203224 328366 203280
rect 328422 203224 328427 203280
rect 328196 203222 328427 203224
rect 328196 203220 328202 203222
rect 328361 203219 328427 203222
rect 331622 203220 331628 203284
rect 331692 203282 331698 203284
rect 332501 203282 332567 203285
rect 331692 203280 332567 203282
rect 331692 203224 332506 203280
rect 332562 203224 332567 203280
rect 331692 203222 332567 203224
rect 331692 203220 331698 203222
rect 332501 203219 332567 203222
rect 332910 203220 332916 203284
rect 332980 203282 332986 203284
rect 333881 203282 333947 203285
rect 332980 203280 333947 203282
rect 332980 203224 333886 203280
rect 333942 203224 333947 203280
rect 332980 203222 333947 203224
rect 332980 203220 332986 203222
rect 333881 203219 333947 203222
rect 335118 203220 335124 203284
rect 335188 203282 335194 203284
rect 335261 203282 335327 203285
rect 335188 203280 335327 203282
rect 335188 203224 335266 203280
rect 335322 203224 335327 203280
rect 335188 203222 335327 203224
rect 335188 203220 335194 203222
rect 335261 203219 335327 203222
rect 338205 203282 338271 203285
rect 338430 203282 338436 203284
rect 338205 203280 338436 203282
rect 338205 203224 338210 203280
rect 338266 203224 338436 203280
rect 338205 203222 338436 203224
rect 338205 203219 338271 203222
rect 338430 203220 338436 203222
rect 338500 203220 338506 203284
rect 339585 203282 339651 203285
rect 339718 203282 339724 203284
rect 339585 203280 339724 203282
rect 339585 203224 339590 203280
rect 339646 203224 339724 203280
rect 339585 203222 339724 203224
rect 339585 203219 339651 203222
rect 339718 203220 339724 203222
rect 339788 203220 339794 203284
rect 346393 203282 346459 203285
rect 346526 203282 346532 203284
rect 346393 203280 346532 203282
rect 346393 203224 346398 203280
rect 346454 203224 346532 203280
rect 346393 203222 346532 203224
rect 346393 203219 346459 203222
rect 346526 203220 346532 203222
rect 346596 203220 346602 203284
rect 349153 203282 349219 203285
rect 356053 203284 356119 203285
rect 366909 203284 366975 203285
rect 349838 203282 349844 203284
rect 349153 203280 349844 203282
rect 349153 203224 349158 203280
rect 349214 203224 349844 203280
rect 349153 203222 349844 203224
rect 349153 203219 349219 203222
rect 349838 203220 349844 203222
rect 349908 203220 349914 203284
rect 356053 203282 356100 203284
rect 356008 203280 356100 203282
rect 356008 203224 356058 203280
rect 356008 203222 356100 203224
rect 356053 203220 356100 203222
rect 356164 203220 356170 203284
rect 366909 203282 366956 203284
rect 366864 203280 366956 203282
rect 366864 203224 366914 203280
rect 366864 203222 366956 203224
rect 366909 203220 366956 203222
rect 367020 203220 367026 203284
rect 368473 203282 368539 203285
rect 368606 203282 368612 203284
rect 368473 203280 368612 203282
rect 368473 203224 368478 203280
rect 368534 203224 368612 203280
rect 368473 203222 368612 203224
rect 356053 203219 356119 203220
rect 366909 203219 366975 203220
rect 368473 203219 368539 203222
rect 368606 203220 368612 203222
rect 368676 203220 368682 203284
rect 370998 203220 371004 203284
rect 371068 203282 371074 203284
rect 371141 203282 371207 203285
rect 371068 203280 371207 203282
rect 371068 203224 371146 203280
rect 371202 203224 371207 203280
rect 371068 203222 371207 203224
rect 371068 203220 371074 203222
rect 371141 203219 371207 203222
rect 375649 203282 375715 203285
rect 385174 203282 385234 203358
rect 375649 203280 385234 203282
rect 375649 203224 375654 203280
rect 375710 203224 385234 203280
rect 375649 203222 385234 203224
rect 442257 203282 442323 203285
rect 451089 203282 451155 203285
rect 442257 203280 451155 203282
rect 442257 203224 442262 203280
rect 442318 203224 451094 203280
rect 451150 203224 451155 203280
rect 442257 203222 451155 203224
rect 455830 203282 455890 203358
rect 456006 203356 456012 203420
rect 456076 203418 456082 203420
rect 456241 203418 456307 203421
rect 456701 203418 456767 203421
rect 461577 203418 461643 203421
rect 456076 203416 456767 203418
rect 456076 203360 456246 203416
rect 456302 203360 456706 203416
rect 456762 203360 456767 203416
rect 456076 203358 456767 203360
rect 456076 203356 456082 203358
rect 456241 203355 456307 203358
rect 456701 203355 456767 203358
rect 458590 203416 461643 203418
rect 458590 203360 461582 203416
rect 461638 203360 461643 203416
rect 458590 203358 461643 203360
rect 458590 203282 458650 203358
rect 461577 203355 461643 203358
rect 462262 203356 462268 203420
rect 462332 203418 462338 203420
rect 463601 203418 463667 203421
rect 464705 203420 464771 203421
rect 464654 203418 464660 203420
rect 462332 203416 463667 203418
rect 462332 203360 463606 203416
rect 463662 203360 463667 203416
rect 462332 203358 463667 203360
rect 464614 203358 464660 203418
rect 464724 203416 464771 203420
rect 464766 203360 464771 203416
rect 462332 203356 462338 203358
rect 463601 203355 463667 203358
rect 464654 203356 464660 203358
rect 464724 203356 464771 203360
rect 464705 203355 464771 203356
rect 467557 203418 467623 203421
rect 469489 203420 469555 203421
rect 469438 203418 469444 203420
rect 467557 203416 469444 203418
rect 469508 203418 469555 203420
rect 477493 203418 477559 203421
rect 478086 203418 478092 203420
rect 469508 203416 469636 203418
rect 467557 203360 467562 203416
rect 467618 203360 469444 203416
rect 469550 203360 469636 203416
rect 467557 203358 469444 203360
rect 467557 203355 467623 203358
rect 469438 203356 469444 203358
rect 469508 203358 469636 203360
rect 477493 203416 478092 203418
rect 477493 203360 477498 203416
rect 477554 203360 478092 203416
rect 477493 203358 478092 203360
rect 469508 203356 469555 203358
rect 469489 203355 469555 203356
rect 477493 203355 477559 203358
rect 478086 203356 478092 203358
rect 478156 203356 478162 203420
rect 478873 203418 478939 203421
rect 479190 203418 479196 203420
rect 478873 203416 479196 203418
rect 478873 203360 478878 203416
rect 478934 203360 479196 203416
rect 478873 203358 479196 203360
rect 478873 203355 478939 203358
rect 479190 203356 479196 203358
rect 479260 203356 479266 203420
rect 480302 203418 480362 203494
rect 480621 203492 480668 203494
rect 480732 203492 480738 203556
rect 484393 203554 484459 203557
rect 484526 203554 484532 203556
rect 484393 203552 484532 203554
rect 484393 203496 484398 203552
rect 484454 203496 484532 203552
rect 484393 203494 484532 203496
rect 480621 203491 480687 203492
rect 484393 203491 484459 203494
rect 484526 203492 484532 203494
rect 484596 203492 484602 203556
rect 488574 203418 488580 203420
rect 480302 203358 488580 203418
rect 488574 203356 488580 203358
rect 488644 203356 488650 203420
rect 455830 203222 458650 203282
rect 375649 203219 375715 203222
rect 442257 203219 442323 203222
rect 451089 203219 451155 203222
rect 458766 203220 458772 203284
rect 458836 203282 458842 203284
rect 459461 203282 459527 203285
rect 458836 203280 459527 203282
rect 458836 203224 459466 203280
rect 459522 203224 459527 203280
rect 458836 203222 459527 203224
rect 458836 203220 458842 203222
rect 459461 203219 459527 203222
rect 460974 203220 460980 203284
rect 461044 203282 461050 203284
rect 462221 203282 462287 203285
rect 461044 203280 462287 203282
rect 461044 203224 462226 203280
rect 462282 203224 462287 203280
rect 461044 203222 462287 203224
rect 461044 203220 461050 203222
rect 462221 203219 462287 203222
rect 463182 203220 463188 203284
rect 463252 203282 463258 203284
rect 463509 203282 463575 203285
rect 463252 203280 463575 203282
rect 463252 203224 463514 203280
rect 463570 203224 463575 203280
rect 463252 203222 463575 203224
rect 463252 203220 463258 203222
rect 463509 203219 463575 203222
rect 467046 203220 467052 203284
rect 467116 203282 467122 203284
rect 467741 203282 467807 203285
rect 467116 203280 467807 203282
rect 467116 203224 467746 203280
rect 467802 203224 467807 203280
rect 467116 203222 467807 203224
rect 467116 203220 467122 203222
rect 467741 203219 467807 203222
rect 470593 203282 470659 203285
rect 471094 203282 471100 203284
rect 470593 203280 471100 203282
rect 470593 203224 470598 203280
rect 470654 203224 471100 203280
rect 470593 203222 471100 203224
rect 470593 203219 470659 203222
rect 471094 203220 471100 203222
rect 471164 203282 471170 203284
rect 471329 203282 471395 203285
rect 471164 203280 471395 203282
rect 471164 203224 471334 203280
rect 471390 203224 471395 203280
rect 471164 203222 471395 203224
rect 471164 203220 471170 203222
rect 471329 203219 471395 203222
rect 471646 203220 471652 203284
rect 471716 203282 471722 203284
rect 471881 203282 471947 203285
rect 471716 203280 471947 203282
rect 471716 203224 471886 203280
rect 471942 203224 471947 203280
rect 471716 203222 471947 203224
rect 471716 203220 471722 203222
rect 471881 203219 471947 203222
rect 472617 203282 472683 203285
rect 472893 203284 472959 203285
rect 472750 203282 472756 203284
rect 472617 203280 472756 203282
rect 472617 203224 472622 203280
rect 472678 203224 472756 203280
rect 472617 203222 472756 203224
rect 472617 203219 472683 203222
rect 472750 203220 472756 203222
rect 472820 203220 472826 203284
rect 472893 203280 472940 203284
rect 473004 203282 473010 203284
rect 473353 203282 473419 203285
rect 473670 203282 473676 203284
rect 472893 203224 472898 203280
rect 472893 203220 472940 203224
rect 473004 203222 473050 203282
rect 473353 203280 473676 203282
rect 473353 203224 473358 203280
rect 473414 203224 473676 203280
rect 473353 203222 473676 203224
rect 473004 203220 473010 203222
rect 472893 203219 472959 203220
rect 473353 203219 473419 203222
rect 473670 203220 473676 203222
rect 473740 203220 473746 203284
rect 474825 203282 474891 203285
rect 474958 203282 474964 203284
rect 474825 203280 474964 203282
rect 474825 203224 474830 203280
rect 474886 203224 474964 203280
rect 474825 203222 474964 203224
rect 474825 203219 474891 203222
rect 474958 203220 474964 203222
rect 475028 203220 475034 203284
rect 477493 203282 477559 203285
rect 477718 203282 477724 203284
rect 477493 203280 477724 203282
rect 477493 203224 477498 203280
rect 477554 203224 477724 203280
rect 477493 203222 477724 203224
rect 477493 203219 477559 203222
rect 477718 203220 477724 203222
rect 477788 203220 477794 203284
rect 478965 203282 479031 203285
rect 479926 203282 479932 203284
rect 478965 203280 479932 203282
rect 478965 203224 478970 203280
rect 479026 203224 479932 203280
rect 478965 203222 479932 203224
rect 478965 203219 479031 203222
rect 479926 203220 479932 203222
rect 479996 203220 480002 203284
rect 481633 203282 481699 203285
rect 482134 203282 482140 203284
rect 481633 203280 482140 203282
rect 481633 203224 481638 203280
rect 481694 203224 482140 203280
rect 481633 203222 482140 203224
rect 481633 203219 481699 203222
rect 482134 203220 482140 203222
rect 482204 203220 482210 203284
rect 328269 203148 328335 203149
rect 332409 203148 332475 203149
rect 328269 203146 328316 203148
rect 328224 203144 328316 203146
rect 328224 203088 328274 203144
rect 328224 203086 328316 203088
rect 328269 203084 328316 203086
rect 328380 203084 328386 203148
rect 332358 203084 332364 203148
rect 332428 203146 332475 203148
rect 332428 203144 332520 203146
rect 332470 203088 332520 203144
rect 332428 203086 332520 203088
rect 332428 203084 332475 203086
rect 333646 203084 333652 203148
rect 333716 203146 333722 203148
rect 333789 203146 333855 203149
rect 336549 203148 336615 203149
rect 336549 203146 336596 203148
rect 333716 203144 333855 203146
rect 333716 203088 333794 203144
rect 333850 203088 333855 203144
rect 333716 203086 333855 203088
rect 336504 203144 336596 203146
rect 336504 203088 336554 203144
rect 336504 203086 336596 203088
rect 333716 203084 333722 203086
rect 328269 203083 328335 203084
rect 332409 203083 332475 203084
rect 333789 203083 333855 203086
rect 336549 203084 336596 203086
rect 336660 203084 336666 203148
rect 343633 203146 343699 203149
rect 343950 203146 343956 203148
rect 343633 203144 343956 203146
rect 343633 203088 343638 203144
rect 343694 203088 343956 203144
rect 343633 203086 343956 203088
rect 336549 203083 336615 203084
rect 343633 203083 343699 203086
rect 343950 203084 343956 203086
rect 344020 203084 344026 203148
rect 345013 203146 345079 203149
rect 351085 203148 351151 203149
rect 345238 203146 345244 203148
rect 345013 203144 345244 203146
rect 345013 203088 345018 203144
rect 345074 203088 345244 203144
rect 345013 203086 345244 203088
rect 345013 203083 345079 203086
rect 345238 203084 345244 203086
rect 345308 203084 345314 203148
rect 351085 203146 351132 203148
rect 351040 203144 351132 203146
rect 351040 203088 351090 203144
rect 351040 203086 351132 203088
rect 351085 203084 351132 203086
rect 351196 203084 351202 203148
rect 357750 203084 357756 203148
rect 357820 203146 357826 203148
rect 357985 203146 358051 203149
rect 357820 203144 358051 203146
rect 357820 203088 357990 203144
rect 358046 203088 358051 203144
rect 357820 203086 358051 203088
rect 357820 203084 357826 203086
rect 351085 203083 351151 203084
rect 357985 203083 358051 203086
rect 360193 203146 360259 203149
rect 360193 203144 365362 203146
rect 360193 203088 360198 203144
rect 360254 203088 365362 203144
rect 360193 203086 365362 203088
rect 360193 203083 360259 203086
rect 334750 202948 334756 203012
rect 334820 203010 334826 203012
rect 335261 203010 335327 203013
rect 334820 203008 335327 203010
rect 334820 202952 335266 203008
rect 335322 202952 335327 203008
rect 334820 202950 335327 202952
rect 334820 202948 334826 202950
rect 335261 202947 335327 202950
rect 336038 202948 336044 203012
rect 336108 203010 336114 203012
rect 336641 203010 336707 203013
rect 337929 203012 337995 203013
rect 339217 203012 339283 203013
rect 337878 203010 337884 203012
rect 336108 203008 336707 203010
rect 336108 202952 336646 203008
rect 336702 202952 336707 203008
rect 336108 202950 336707 202952
rect 337838 202950 337884 203010
rect 337948 203008 337995 203012
rect 339166 203010 339172 203012
rect 337990 202952 337995 203008
rect 336108 202948 336114 202950
rect 336641 202947 336707 202950
rect 337878 202948 337884 202950
rect 337948 202948 337995 202952
rect 339126 202950 339172 203010
rect 339236 203008 339283 203012
rect 339278 202952 339283 203008
rect 339166 202948 339172 202950
rect 339236 202948 339283 202952
rect 337929 202947 337995 202948
rect 339217 202947 339283 202948
rect 341333 203012 341399 203013
rect 344921 203012 344987 203013
rect 341333 203008 341380 203012
rect 341444 203010 341450 203012
rect 344870 203010 344876 203012
rect 341333 202952 341338 203008
rect 341333 202948 341380 202952
rect 341444 202950 341490 203010
rect 344830 202950 344876 203010
rect 344940 203008 344987 203012
rect 344982 202952 344987 203008
rect 341444 202948 341450 202950
rect 344870 202948 344876 202950
rect 344940 202948 344987 202952
rect 341333 202947 341399 202948
rect 344921 202947 344987 202948
rect 345933 203012 345999 203013
rect 347037 203012 347103 203013
rect 348417 203012 348483 203013
rect 345933 203008 345980 203012
rect 346044 203010 346050 203012
rect 345933 202952 345938 203008
rect 345933 202948 345980 202952
rect 346044 202950 346090 203010
rect 347037 203008 347084 203012
rect 347148 203010 347154 203012
rect 348366 203010 348372 203012
rect 347037 202952 347042 203008
rect 346044 202948 346050 202950
rect 347037 202948 347084 202952
rect 347148 202950 347194 203010
rect 348326 202950 348372 203010
rect 348436 203008 348483 203012
rect 348478 202952 348483 203008
rect 347148 202948 347154 202950
rect 348366 202948 348372 202950
rect 348436 202948 348483 202952
rect 345933 202947 345999 202948
rect 347037 202947 347103 202948
rect 348417 202947 348483 202948
rect 349429 203012 349495 203013
rect 349429 203008 349476 203012
rect 349540 203010 349546 203012
rect 349429 202952 349434 203008
rect 349429 202948 349476 202952
rect 349540 202950 349586 203010
rect 349540 202948 349546 202950
rect 350942 202948 350948 203012
rect 351012 203010 351018 203012
rect 351177 203010 351243 203013
rect 351012 203008 351243 203010
rect 351012 202952 351182 203008
rect 351238 202952 351243 203008
rect 351012 202950 351243 202952
rect 351012 202948 351018 202950
rect 349429 202947 349495 202948
rect 351177 202947 351243 202950
rect 351637 203012 351703 203013
rect 353017 203012 353083 203013
rect 351637 203008 351684 203012
rect 351748 203010 351754 203012
rect 352966 203010 352972 203012
rect 351637 202952 351642 203008
rect 351637 202948 351684 202952
rect 351748 202950 351794 203010
rect 352926 202950 352972 203010
rect 353036 203008 353083 203012
rect 353293 203012 353359 203013
rect 353293 203010 353340 203012
rect 353078 202952 353083 203008
rect 351748 202948 351754 202950
rect 352966 202948 352972 202950
rect 353036 202948 353083 202952
rect 353248 203008 353340 203010
rect 353248 202952 353298 203008
rect 353248 202950 353340 202952
rect 351637 202947 351703 202948
rect 353017 202947 353083 202948
rect 353293 202948 353340 202950
rect 353404 202948 353410 203012
rect 354438 202948 354444 203012
rect 354508 203010 354514 203012
rect 354581 203010 354647 203013
rect 355593 203012 355659 203013
rect 355542 203010 355548 203012
rect 354508 203008 354647 203010
rect 354508 202952 354586 203008
rect 354642 202952 354647 203008
rect 354508 202950 354647 202952
rect 355502 202950 355548 203010
rect 355612 203008 355659 203012
rect 355654 202952 355659 203008
rect 354508 202948 354514 202950
rect 353293 202947 353359 202948
rect 354581 202947 354647 202950
rect 355542 202948 355548 202950
rect 355612 202948 355659 202952
rect 355593 202947 355659 202948
rect 356421 203012 356487 203013
rect 356421 203008 356468 203012
rect 356532 203010 356538 203012
rect 357433 203010 357499 203013
rect 358629 203012 358695 203013
rect 357934 203010 357940 203012
rect 356421 202952 356426 203008
rect 356421 202948 356468 202952
rect 356532 202950 356578 203010
rect 357433 203008 357940 203010
rect 357433 202952 357438 203008
rect 357494 202952 357940 203008
rect 357433 202950 357940 202952
rect 356532 202948 356538 202950
rect 356421 202947 356487 202948
rect 357433 202947 357499 202950
rect 357934 202948 357940 202950
rect 358004 202948 358010 203012
rect 358629 203010 358676 203012
rect 358584 203008 358676 203010
rect 358584 202952 358634 203008
rect 358584 202950 358676 202952
rect 358629 202948 358676 202950
rect 358740 202948 358746 203012
rect 358813 203010 358879 203013
rect 360009 203012 360075 203013
rect 361297 203012 361363 203013
rect 359222 203010 359228 203012
rect 358813 203008 359228 203010
rect 358813 202952 358818 203008
rect 358874 202952 359228 203008
rect 358813 202950 359228 202952
rect 358629 202947 358695 202948
rect 358813 202947 358879 202950
rect 359222 202948 359228 202950
rect 359292 202948 359298 203012
rect 359958 203010 359964 203012
rect 359918 202950 359964 203010
rect 360028 203008 360075 203012
rect 361246 203010 361252 203012
rect 360070 202952 360075 203008
rect 359958 202948 359964 202950
rect 360028 202948 360075 202952
rect 361206 202950 361252 203010
rect 361316 203008 361363 203012
rect 361358 202952 361363 203008
rect 361246 202948 361252 202950
rect 361316 202948 361363 202952
rect 362718 202948 362724 203012
rect 362788 203010 362794 203012
rect 362861 203010 362927 203013
rect 362788 203008 362927 203010
rect 362788 202952 362866 203008
rect 362922 202952 362927 203008
rect 362788 202950 362927 202952
rect 362788 202948 362794 202950
rect 360009 202947 360075 202948
rect 361297 202947 361363 202948
rect 362861 202947 362927 202950
rect 363413 203012 363479 203013
rect 363413 203008 363460 203012
rect 363524 203010 363530 203012
rect 363413 202952 363418 203008
rect 363413 202948 363460 202952
rect 363524 202950 363570 203010
rect 363524 202948 363530 202950
rect 364926 202948 364932 203012
rect 364996 203010 365002 203012
rect 365069 203010 365135 203013
rect 364996 203008 365135 203010
rect 364996 202952 365074 203008
rect 365130 202952 365135 203008
rect 364996 202950 365135 202952
rect 365302 203010 365362 203086
rect 366398 203084 366404 203148
rect 366468 203146 366474 203148
rect 367001 203146 367067 203149
rect 366468 203144 367067 203146
rect 366468 203088 367006 203144
rect 367062 203088 367067 203144
rect 366468 203086 367067 203088
rect 366468 203084 366474 203086
rect 367001 203083 367067 203086
rect 373257 203146 373323 203149
rect 373390 203146 373396 203148
rect 373257 203144 373396 203146
rect 373257 203088 373262 203144
rect 373318 203088 373396 203144
rect 373257 203086 373396 203088
rect 373257 203083 373323 203086
rect 373390 203084 373396 203086
rect 373460 203146 373466 203148
rect 492806 203146 492812 203148
rect 373460 203086 492812 203146
rect 373460 203084 373466 203086
rect 492806 203084 492812 203086
rect 492876 203084 492882 203148
rect 375649 203010 375715 203013
rect 365302 203008 375715 203010
rect 365302 202952 375654 203008
rect 375710 202952 375715 203008
rect 365302 202950 375715 202952
rect 364996 202948 365002 202950
rect 363413 202947 363479 202948
rect 365069 202947 365135 202950
rect 375649 202947 375715 202950
rect 450670 202948 450676 203012
rect 450740 203010 450746 203012
rect 450997 203010 451063 203013
rect 450740 203008 451063 203010
rect 450740 202952 451002 203008
rect 451058 202952 451063 203008
rect 450740 202950 451063 202952
rect 450740 202948 450746 202950
rect 450997 202947 451063 202950
rect 452878 202948 452884 203012
rect 452948 203010 452954 203012
rect 453941 203010 454007 203013
rect 455321 203012 455387 203013
rect 457897 203012 457963 203013
rect 452948 203008 454007 203010
rect 452948 202952 453946 203008
rect 454002 202952 454007 203008
rect 452948 202950 454007 202952
rect 452948 202948 452954 202950
rect 453941 202947 454007 202950
rect 455270 202948 455276 203012
rect 455340 203010 455387 203012
rect 457846 203010 457852 203012
rect 455340 203008 455432 203010
rect 455382 202952 455432 203008
rect 455340 202950 455432 202952
rect 457806 202950 457852 203010
rect 457916 203008 457963 203012
rect 457958 202952 457963 203008
rect 455340 202948 455387 202950
rect 457846 202948 457852 202950
rect 457916 202948 457963 202952
rect 458950 202948 458956 203012
rect 459020 203010 459026 203012
rect 459093 203010 459159 203013
rect 460657 203012 460723 203013
rect 460606 203010 460612 203012
rect 459020 203008 459159 203010
rect 459020 202952 459098 203008
rect 459154 202952 459159 203008
rect 459020 202950 459159 202952
rect 460566 202950 460612 203010
rect 460676 203008 460723 203012
rect 460718 202952 460723 203008
rect 459020 202948 459026 202950
rect 455321 202947 455387 202948
rect 457897 202947 457963 202948
rect 459093 202947 459159 202950
rect 460606 202948 460612 202950
rect 460676 202948 460723 202952
rect 460657 202947 460723 202948
rect 461485 203012 461551 203013
rect 462405 203012 462471 203013
rect 461485 203008 461532 203012
rect 461596 203010 461602 203012
rect 461485 202952 461490 203008
rect 461485 202948 461532 202952
rect 461596 202950 461642 203010
rect 462405 203008 462452 203012
rect 462516 203010 462522 203012
rect 463049 203010 463115 203013
rect 465901 203012 465967 203013
rect 467189 203012 467255 203013
rect 468477 203012 468543 203013
rect 463550 203010 463556 203012
rect 462405 202952 462410 203008
rect 461596 202948 461602 202950
rect 462405 202948 462452 202952
rect 462516 202950 462562 203010
rect 463049 203008 463556 203010
rect 463049 202952 463054 203008
rect 463110 202952 463556 203008
rect 463049 202950 463556 202952
rect 462516 202948 462522 202950
rect 461485 202947 461551 202948
rect 462405 202947 462471 202948
rect 463049 202947 463115 202950
rect 463550 202948 463556 202950
rect 463620 202948 463626 203012
rect 465901 203008 465948 203012
rect 466012 203010 466018 203012
rect 465901 202952 465906 203008
rect 465901 202948 465948 202952
rect 466012 202950 466058 203010
rect 467189 203008 467236 203012
rect 467300 203010 467306 203012
rect 467189 202952 467194 203008
rect 466012 202948 466018 202950
rect 467189 202948 467236 202952
rect 467300 202950 467346 203010
rect 468477 203008 468524 203012
rect 468588 203010 468594 203012
rect 471053 203010 471119 203013
rect 471789 203012 471855 203013
rect 471789 203010 471836 203012
rect 468477 202952 468482 203008
rect 467300 202948 467306 202950
rect 468477 202948 468524 202952
rect 468588 202950 468634 203010
rect 471053 203008 471836 203010
rect 471053 202952 471058 203008
rect 471114 202952 471794 203008
rect 471053 202950 471836 202952
rect 468588 202948 468594 202950
rect 465901 202947 465967 202948
rect 467189 202947 467255 202948
rect 468477 202947 468543 202948
rect 471053 202947 471119 202950
rect 471789 202948 471836 202950
rect 471900 202948 471906 203012
rect 475510 202948 475516 203012
rect 475580 203010 475586 203012
rect 475745 203010 475811 203013
rect 475580 203008 475811 203010
rect 475580 202952 475750 203008
rect 475806 202952 475811 203008
rect 475580 202950 475811 202952
rect 475580 202948 475586 202950
rect 471789 202947 471855 202948
rect 475745 202947 475811 202950
rect 476113 203010 476179 203013
rect 476430 203010 476436 203012
rect 476113 203008 476436 203010
rect 476113 202952 476118 203008
rect 476174 202952 476436 203008
rect 476113 202950 476436 202952
rect 476113 202947 476179 202950
rect 476430 202948 476436 202950
rect 476500 202948 476506 203012
rect 477493 203010 477559 203013
rect 478638 203010 478644 203012
rect 477493 203008 478644 203010
rect 477493 202952 477498 203008
rect 477554 202952 478644 203008
rect 477493 202950 478644 202952
rect 477493 202947 477559 202950
rect 478638 202948 478644 202950
rect 478708 202948 478714 203012
rect 480529 203010 480595 203013
rect 481030 203010 481036 203012
rect 480529 203008 481036 203010
rect 480529 202952 480534 203008
rect 480590 202952 481036 203008
rect 480529 202950 481036 202952
rect 480529 202947 480595 202950
rect 481030 202948 481036 202950
rect 481100 202948 481106 203012
rect 481633 203010 481699 203013
rect 483013 203012 483079 203013
rect 481766 203010 481772 203012
rect 481633 203008 481772 203010
rect 481633 202952 481638 203008
rect 481694 202952 481772 203008
rect 481633 202950 481772 202952
rect 481633 202947 481699 202950
rect 481766 202948 481772 202950
rect 481836 202948 481842 203012
rect 483013 203010 483060 203012
rect 482968 203008 483060 203010
rect 482968 202952 483018 203008
rect 482968 202950 483060 202952
rect 483013 202948 483060 202950
rect 483124 202948 483130 203012
rect 483013 202947 483079 202948
rect 342294 201724 342300 201788
rect 342364 201724 342370 201788
rect 342302 201516 342362 201724
rect 342270 201452 342276 201516
rect 342340 201454 342362 201516
rect 342340 201452 342346 201454
rect 448421 201380 448487 201381
rect 448378 201378 448384 201380
rect 448330 201318 448384 201378
rect 448448 201376 448487 201380
rect 448482 201320 448487 201376
rect 448378 201316 448384 201318
rect 448448 201316 448487 201320
rect 448421 201315 448487 201316
rect 3693 200834 3759 200837
rect 522614 200834 522620 200836
rect 3693 200832 522620 200834
rect 3693 200776 3698 200832
rect 3754 200776 522620 200832
rect 3693 200774 522620 200776
rect 3693 200771 3759 200774
rect 522614 200772 522620 200774
rect 522684 200772 522690 200836
rect 3509 200698 3575 200701
rect 522430 200698 522436 200700
rect 3509 200696 522436 200698
rect 3509 200640 3514 200696
rect 3570 200640 522436 200696
rect 3509 200638 522436 200640
rect 3509 200635 3575 200638
rect 522430 200636 522436 200638
rect 522500 200636 522506 200700
rect -960 193898 480 193988
rect 2957 193898 3023 193901
rect -960 193896 3023 193898
rect -960 193840 2962 193896
rect 3018 193840 3023 193896
rect -960 193838 3023 193840
rect -960 193748 480 193838
rect 2957 193835 3023 193838
rect 583520 193476 584960 193716
rect 500309 183154 500375 183157
rect 497230 183152 500375 183154
rect 497230 183096 500314 183152
rect 500370 183096 500375 183152
rect 497230 183094 500375 183096
rect 379789 182746 379855 182749
rect 377814 182744 379855 182746
rect 377814 182722 379794 182744
rect 377292 182688 379794 182722
rect 379850 182688 379855 182744
rect 497230 182692 497290 183094
rect 500309 183091 500375 183094
rect 377292 182686 379855 182688
rect 377292 182662 377874 182686
rect 379789 182683 379855 182686
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect 496445 181386 496511 181389
rect 496445 181384 496554 181386
rect 496445 181328 496450 181384
rect 496506 181328 496554 181384
rect 496445 181323 496554 181328
rect 377292 180978 377874 181022
rect 496494 180992 496554 181323
rect 380525 180978 380591 180981
rect 377292 180976 380591 180978
rect 377292 180962 380530 180976
rect 377814 180920 380530 180962
rect 380586 180920 380591 180976
rect 377814 180918 380591 180920
rect 380525 180915 380591 180918
rect 417417 180570 417483 180573
rect 417417 180568 420378 180570
rect 417417 180512 417422 180568
rect 417478 180512 420378 180568
rect 417417 180510 420378 180512
rect 417417 180507 417483 180510
rect 297909 180298 297975 180301
rect 300166 180298 300226 180319
rect 297909 180296 300226 180298
rect 297909 180240 297914 180296
rect 297970 180240 300226 180296
rect 297909 180238 300226 180240
rect 297909 180235 297975 180238
rect -960 179482 480 179572
rect 3877 179482 3943 179485
rect -960 179480 3943 179482
rect -960 179424 3882 179480
rect 3938 179424 3943 179480
rect -960 179422 3943 179424
rect -960 179332 480 179422
rect 3877 179419 3943 179422
rect 297909 171866 297975 171869
rect 297909 171865 299674 171866
rect 300166 171865 300226 180238
rect 420318 171865 420378 180510
rect 297909 171864 300226 171865
rect 297909 171808 297914 171864
rect 297970 171835 300226 171864
rect 420164 171835 420378 171865
rect 297970 171808 300196 171835
rect 297909 171806 300196 171808
rect 297909 171803 297975 171806
rect 299614 171805 300196 171806
rect 420134 171805 420348 171835
rect 418061 171730 418127 171733
rect 420134 171730 420194 171805
rect 418061 171728 420194 171730
rect 418061 171672 418066 171728
rect 418122 171672 420194 171728
rect 418061 171670 420194 171672
rect 418061 171667 418127 171670
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3785 165066 3851 165069
rect -960 165064 3851 165066
rect -960 165008 3790 165064
rect 3846 165008 3851 165064
rect -960 165006 3851 165008
rect -960 164916 480 165006
rect 3785 165003 3851 165006
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect -960 150786 480 150876
rect 3601 150786 3667 150789
rect -960 150784 3667 150786
rect -960 150728 3606 150784
rect 3662 150728 3667 150784
rect -960 150726 3667 150728
rect -960 150636 480 150726
rect 3601 150723 3667 150726
rect 583520 146556 584960 146796
rect -960 136370 480 136460
rect 3693 136370 3759 136373
rect -960 136368 3759 136370
rect -960 136312 3698 136368
rect 3754 136312 3759 136368
rect -960 136310 3759 136312
rect -960 136220 480 136310
rect 3693 136307 3759 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 500125 123722 500191 123725
rect 497230 123720 500191 123722
rect 497230 123664 500130 123720
rect 500186 123664 500191 123720
rect 497230 123662 500191 123664
rect 379973 123178 380039 123181
rect 377814 123176 380039 123178
rect 377814 123174 379978 123176
rect 377292 123120 379978 123174
rect 380034 123120 380039 123176
rect 497230 123144 497290 123662
rect 500125 123659 500191 123662
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 377292 123118 380039 123120
rect 377292 123114 377874 123118
rect 379973 123115 380039 123118
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3509 122090 3575 122093
rect 380433 122090 380499 122093
rect 500033 122090 500099 122093
rect -960 122088 3575 122090
rect -960 122032 3514 122088
rect 3570 122032 3575 122088
rect -960 122030 3575 122032
rect -960 121940 480 122030
rect 3509 122027 3575 122030
rect 377078 122088 380499 122090
rect 377078 122032 380438 122088
rect 380494 122032 380499 122088
rect 377078 122030 380499 122032
rect 377078 121444 377138 122030
rect 380433 122027 380499 122030
rect 497230 122088 500099 122090
rect 497230 122032 500038 122088
rect 500094 122032 500099 122088
rect 497230 122030 500099 122032
rect 497230 121444 497290 122030
rect 500033 122027 500099 122030
rect 499941 120866 500007 120869
rect 497230 120864 500007 120866
rect 497230 120808 499946 120864
rect 500002 120808 500007 120864
rect 497230 120806 500007 120808
rect 377292 120322 377874 120346
rect 380341 120322 380407 120325
rect 377292 120320 380407 120322
rect 377292 120286 380346 120320
rect 377814 120264 380346 120286
rect 380402 120264 380407 120320
rect 497230 120316 497290 120806
rect 499941 120803 500007 120806
rect 377814 120262 380407 120264
rect 380341 120259 380407 120262
rect 380249 118690 380315 118693
rect 499757 118690 499823 118693
rect 377814 118688 380315 118690
rect 377814 118646 380254 118688
rect 377292 118632 380254 118646
rect 380310 118632 380315 118688
rect 377292 118630 380315 118632
rect 377292 118586 377874 118630
rect 380249 118627 380315 118630
rect 497230 118688 499823 118690
rect 497230 118632 499762 118688
rect 499818 118632 499823 118688
rect 497230 118630 499823 118632
rect 497230 118616 497290 118630
rect 499757 118627 499823 118630
rect 380065 118146 380131 118149
rect 499849 118146 499915 118149
rect 377078 118144 380131 118146
rect 377078 118088 380070 118144
rect 380126 118088 380131 118144
rect 377078 118086 380131 118088
rect 377078 117488 377138 118086
rect 380065 118083 380131 118086
rect 497230 118144 499915 118146
rect 497230 118088 499854 118144
rect 499910 118088 499915 118144
rect 497230 118086 499915 118088
rect 497230 117488 497290 118086
rect 499849 118083 499915 118086
rect 380157 115834 380223 115837
rect 500217 115834 500283 115837
rect 377814 115832 380223 115834
rect 377814 115818 380162 115832
rect 377292 115776 380162 115818
rect 380218 115776 380223 115832
rect 377292 115774 380223 115776
rect 497230 115832 500283 115834
rect 497230 115776 500222 115832
rect 500278 115776 500283 115832
rect 497230 115774 500283 115776
rect 377292 115758 377874 115774
rect 380157 115771 380223 115774
rect 500217 115771 500283 115774
rect 499665 115290 499731 115293
rect 497230 115288 499731 115290
rect 497230 115232 499670 115288
rect 499726 115232 499731 115288
rect 497230 115230 499731 115232
rect 379973 114746 380039 114749
rect 377814 114744 380039 114746
rect 377814 114690 379978 114744
rect 377292 114688 379978 114690
rect 380034 114688 380039 114744
rect 377292 114686 380039 114688
rect 377292 114630 377874 114686
rect 379973 114683 380039 114686
rect 497230 114660 497290 115230
rect 499665 115227 499731 115230
rect 297817 111754 297883 111757
rect 297817 111752 300778 111754
rect 297817 111696 297822 111752
rect 297878 111696 300778 111752
rect 297817 111694 300778 111696
rect 297817 111691 297883 111694
rect 300718 111349 300778 111694
rect 300718 111344 300827 111349
rect 300718 111288 300766 111344
rect 300822 111288 300827 111344
rect 300718 111286 300827 111288
rect 300761 111283 300827 111286
rect 416773 111346 416839 111349
rect 420134 111346 420194 111564
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 416773 111344 420194 111346
rect 416773 111288 416778 111344
rect 416834 111288 420194 111344
rect 583520 111332 584960 111422
rect 416773 111286 420194 111288
rect 416773 111283 416839 111286
rect 303613 109036 303679 109037
rect 303613 109032 303660 109036
rect 303724 109034 303730 109036
rect 307753 109034 307819 109037
rect 424225 109036 424291 109037
rect 308070 109034 308076 109036
rect 303613 108976 303618 109032
rect 303613 108972 303660 108976
rect 303724 108974 303770 109034
rect 307753 109032 308076 109034
rect 307753 108976 307758 109032
rect 307814 108976 308076 109032
rect 307753 108974 308076 108976
rect 303724 108972 303730 108974
rect 303613 108971 303679 108972
rect 307753 108971 307819 108974
rect 308070 108972 308076 108974
rect 308140 108972 308146 109036
rect 424174 109034 424180 109036
rect 424134 108974 424180 109034
rect 424244 109032 424291 109036
rect 424286 108976 424291 109032
rect 424174 108972 424180 108974
rect 424244 108972 424291 108976
rect 424225 108971 424291 108972
rect 427813 109034 427879 109037
rect 428038 109034 428044 109036
rect 427813 109032 428044 109034
rect 427813 108976 427818 109032
rect 427874 108976 428044 109032
rect 427813 108974 428044 108976
rect 427813 108971 427879 108974
rect 428038 108972 428044 108974
rect 428108 108972 428114 109036
rect 3509 108898 3575 108901
rect 520406 108898 520412 108900
rect 3509 108896 520412 108898
rect 3509 108840 3514 108896
rect 3570 108840 520412 108896
rect 3509 108838 520412 108840
rect 3509 108835 3575 108838
rect 520406 108836 520412 108838
rect 520476 108836 520482 108900
rect -960 107674 480 107764
rect 3509 107674 3575 107677
rect -960 107672 3575 107674
rect -960 107616 3514 107672
rect 3570 107616 3575 107672
rect -960 107614 3575 107616
rect -960 107524 480 107614
rect 3509 107611 3575 107614
rect 583520 99636 584960 99876
rect 522246 93802 522252 93804
rect 614 93742 522252 93802
rect -960 93258 480 93348
rect 614 93258 674 93742
rect 522246 93740 522252 93742
rect 522316 93740 522322 93804
rect -960 93198 674 93258
rect -960 93108 480 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 3509 80066 3575 80069
rect 522062 80066 522068 80068
rect 3509 80064 522068 80066
rect 3509 80008 3514 80064
rect 3570 80008 522068 80064
rect 3509 80006 522068 80008
rect 3509 80003 3575 80006
rect 522062 80004 522068 80006
rect 522132 80004 522138 80068
rect -960 78978 480 79068
rect 3509 78978 3575 78981
rect -960 78976 3575 78978
rect -960 78920 3514 78976
rect 3570 78920 3575 78976
rect -960 78918 3575 78920
rect -960 78828 480 78918
rect 3509 78915 3575 78918
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 520222 64834 520228 64836
rect 614 64774 520228 64834
rect -960 64562 480 64652
rect 614 64562 674 64774
rect 520222 64772 520228 64774
rect 520292 64772 520298 64836
rect -960 64502 674 64562
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect -960 64412 480 64502
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect 3325 50962 3391 50965
rect 521878 50962 521884 50964
rect 3325 50960 521884 50962
rect 3325 50904 3330 50960
rect 3386 50904 521884 50960
rect 3325 50902 521884 50904
rect 3325 50899 3391 50902
rect 521878 50900 521884 50902
rect 521948 50900 521954 50964
rect -960 50146 480 50236
rect 3325 50146 3391 50149
rect -960 50144 3391 50146
rect -960 50088 3330 50144
rect 3386 50088 3391 50144
rect -960 50086 3391 50088
rect -960 49996 480 50086
rect 3325 50083 3391 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 521694 35866 521700 35868
rect -960 35806 521700 35866
rect -960 35716 480 35806
rect 521694 35804 521700 35806
rect 521764 35804 521770 35868
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 3417 21450 3483 21453
rect -960 21448 3483 21450
rect -960 21392 3422 21448
rect 3478 21392 3483 21448
rect -960 21390 3483 21392
rect -960 21300 480 21390
rect 3417 21387 3483 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
<< via3 >>
rect 520596 700708 520660 700772
rect 518940 700572 519004 700636
rect 520780 700436 520844 700500
rect 519492 695540 519556 695604
rect 519492 695268 519556 695332
rect 519676 686080 519740 686084
rect 519676 686024 519690 686080
rect 519690 686024 519740 686080
rect 519676 686020 519740 686024
rect 519860 684388 519924 684452
rect 542492 684448 542556 684452
rect 542492 684392 542506 684448
rect 542506 684392 542556 684448
rect 542492 684388 542556 684392
rect 519308 681804 519372 681868
rect 542492 678872 542556 678876
rect 542492 678816 542542 678872
rect 542542 678816 542556 678872
rect 542492 678812 542556 678816
rect 520964 667932 521028 667996
rect 520044 666572 520108 666636
rect 519492 659636 519556 659700
rect 520044 659636 520108 659700
rect 519492 652836 519556 652900
rect 519124 644540 519188 644604
rect 519860 644540 519924 644604
rect 519124 644404 519188 644468
rect 519676 644404 519740 644468
rect 519124 634884 519188 634948
rect 519676 634884 519740 634948
rect 519124 625092 519188 625156
rect 519860 625092 519924 625156
rect 519676 623732 519740 623796
rect 519124 615572 519188 615636
rect 519860 615572 519924 615636
rect 373580 612776 373644 612780
rect 373580 612720 373630 612776
rect 373630 612720 373644 612776
rect 373580 612716 373644 612720
rect 488580 612776 488644 612780
rect 488580 612720 488594 612776
rect 488594 612720 488644 612776
rect 488580 612716 488644 612720
rect 493916 612776 493980 612780
rect 493916 612720 493966 612776
rect 493966 612720 493980 612776
rect 493916 612716 493980 612720
rect 369164 610948 369228 611012
rect 373028 610948 373092 611012
rect 519124 605780 519188 605844
rect 519860 605780 519924 605844
rect 519124 596260 519188 596324
rect 519860 596260 519924 596324
rect 519124 586332 519188 586396
rect 519860 586332 519924 586396
rect 519124 576812 519188 576876
rect 519860 576812 519924 576876
rect 519124 567020 519188 567084
rect 519860 567020 519924 567084
rect 519124 557500 519188 557564
rect 519860 557500 519924 557564
rect 519124 547708 519188 547772
rect 519860 547708 519924 547772
rect 519124 538188 519188 538252
rect 519860 538188 519924 538252
rect 519124 528396 519188 528460
rect 519860 528396 519924 528460
rect 427968 519692 428032 519756
rect 519124 518876 519188 518940
rect 519860 518876 519924 518940
rect 313780 518740 313844 518804
rect 316172 518740 316236 518804
rect 318564 518740 318628 518804
rect 321692 518800 321756 518804
rect 321692 518744 321742 518800
rect 321742 518744 321756 518800
rect 321692 518740 321756 518744
rect 323164 518800 323228 518804
rect 323164 518744 323178 518800
rect 323178 518744 323228 518800
rect 323164 518740 323228 518744
rect 324452 518740 324516 518804
rect 325188 518740 325252 518804
rect 326476 518800 326540 518804
rect 326476 518744 326490 518800
rect 326490 518744 326540 518800
rect 326476 518740 326540 518744
rect 327212 518800 327276 518804
rect 327212 518744 327226 518800
rect 327226 518744 327276 518800
rect 327212 518740 327276 518744
rect 328868 518800 328932 518804
rect 328868 518744 328918 518800
rect 328918 518744 328932 518800
rect 328868 518740 328932 518744
rect 330156 518800 330220 518804
rect 330156 518744 330170 518800
rect 330170 518744 330220 518800
rect 330156 518740 330220 518744
rect 332364 518800 332428 518804
rect 332364 518744 332378 518800
rect 332378 518744 332428 518800
rect 332364 518740 332428 518744
rect 335492 518800 335556 518804
rect 335492 518744 335542 518800
rect 335542 518744 335556 518800
rect 335492 518740 335556 518744
rect 337148 518800 337212 518804
rect 337148 518744 337198 518800
rect 337198 518744 337212 518800
rect 337148 518740 337212 518744
rect 339356 518740 339420 518804
rect 340460 518800 340524 518804
rect 340460 518744 340510 518800
rect 340510 518744 340524 518800
rect 340460 518740 340524 518744
rect 341564 518800 341628 518804
rect 341564 518744 341614 518800
rect 341614 518744 341628 518800
rect 341564 518740 341628 518744
rect 343036 518800 343100 518804
rect 343036 518744 343050 518800
rect 343050 518744 343100 518800
rect 343036 518740 343100 518744
rect 344140 518800 344204 518804
rect 344140 518744 344190 518800
rect 344190 518744 344204 518800
rect 344140 518740 344204 518744
rect 345428 518800 345492 518804
rect 345428 518744 345478 518800
rect 345478 518744 345492 518800
rect 345428 518740 345492 518744
rect 346532 518800 346596 518804
rect 346532 518744 346546 518800
rect 346546 518744 346596 518800
rect 346532 518740 346596 518744
rect 347636 518800 347700 518804
rect 347636 518744 347686 518800
rect 347686 518744 347700 518800
rect 347636 518740 347700 518744
rect 348556 518800 348620 518804
rect 348556 518744 348606 518800
rect 348606 518744 348620 518800
rect 348556 518740 348620 518744
rect 443132 518800 443196 518804
rect 443132 518744 443182 518800
rect 443182 518744 443196 518800
rect 443132 518740 443196 518744
rect 451228 518800 451292 518804
rect 451228 518744 451278 518800
rect 451278 518744 451292 518800
rect 451228 518740 451292 518744
rect 452516 518800 452580 518804
rect 452516 518744 452566 518800
rect 452566 518744 452580 518800
rect 452516 518740 452580 518744
rect 453620 518800 453684 518804
rect 453620 518744 453670 518800
rect 453670 518744 453684 518800
rect 453620 518740 453684 518744
rect 460428 518740 460492 518804
rect 461164 518740 461228 518804
rect 462452 518740 462516 518804
rect 314700 518604 314764 518668
rect 317276 518664 317340 518668
rect 317276 518608 317326 518664
rect 317326 518608 317340 518664
rect 317276 518604 317340 518608
rect 319668 518604 319732 518668
rect 324268 518604 324332 518668
rect 331260 518664 331324 518668
rect 331260 518608 331274 518664
rect 331274 518608 331324 518664
rect 331260 518604 331324 518608
rect 338068 518664 338132 518668
rect 338068 518608 338118 518664
rect 338118 518608 338132 518664
rect 338068 518604 338132 518608
rect 429700 518604 429764 518668
rect 454724 518604 454788 518668
rect 456012 518664 456076 518668
rect 456012 518608 456062 518664
rect 456062 518608 456076 518664
rect 456012 518604 456076 518608
rect 457116 518604 457180 518668
rect 458404 518604 458468 518668
rect 459508 518664 459572 518668
rect 459508 518608 459558 518664
rect 459558 518608 459572 518664
rect 459508 518604 459572 518608
rect 465212 518604 465276 518668
rect 467420 518604 467484 518668
rect 316540 518468 316604 518532
rect 318564 518468 318628 518532
rect 327948 518468 328012 518532
rect 333468 518528 333532 518532
rect 333468 518472 333482 518528
rect 333482 518472 333532 518528
rect 333468 518468 333532 518472
rect 334204 518528 334268 518532
rect 334204 518472 334218 518528
rect 334218 518472 334268 518528
rect 334204 518468 334268 518472
rect 426572 518468 426636 518532
rect 445340 518528 445404 518532
rect 445340 518472 445390 518528
rect 445390 518472 445404 518528
rect 445340 518468 445404 518472
rect 446628 518528 446692 518532
rect 446628 518472 446642 518528
rect 446642 518472 446692 518528
rect 446628 518468 446692 518472
rect 447732 518468 447796 518532
rect 466500 518528 466564 518532
rect 466500 518472 466514 518528
rect 466514 518472 466564 518528
rect 466500 518468 466564 518472
rect 312492 518332 312556 518396
rect 317460 518392 317524 518396
rect 317460 518336 317474 518392
rect 317474 518336 317524 518392
rect 317460 518332 317524 518336
rect 320772 518332 320836 518396
rect 430804 518332 430868 518396
rect 442028 518392 442092 518396
rect 442028 518336 442078 518392
rect 442078 518336 442092 518392
rect 442028 518332 442092 518336
rect 444052 518332 444116 518396
rect 448836 518392 448900 518396
rect 448836 518336 448850 518392
rect 448850 518336 448900 518392
rect 448836 518332 448900 518336
rect 449940 518392 450004 518396
rect 449940 518336 449954 518392
rect 449954 518336 450004 518392
rect 449940 518332 450004 518336
rect 463924 518332 463988 518396
rect 468524 518332 468588 518396
rect 303660 518256 303724 518260
rect 303660 518200 303674 518256
rect 303674 518200 303724 518256
rect 303660 518196 303724 518200
rect 315068 518196 315132 518260
rect 323532 518196 323596 518260
rect 423812 518196 423876 518260
rect 429148 518256 429212 518260
rect 429148 518200 429198 518256
rect 429198 518200 429212 518256
rect 429148 518196 429212 518200
rect 320036 518060 320100 518124
rect 322060 518060 322124 518124
rect 435036 518060 435100 518124
rect 312676 517924 312740 517988
rect 331444 517924 331508 517988
rect 332732 517924 332796 517988
rect 437244 517984 437308 517988
rect 437244 517928 437294 517984
rect 437294 517928 437308 517984
rect 437244 517924 437308 517928
rect 320956 517788 321020 517852
rect 334940 517788 335004 517852
rect 432644 517848 432708 517852
rect 432644 517792 432658 517848
rect 432658 517792 432708 517848
rect 432644 517788 432708 517792
rect 433748 517788 433812 517852
rect 440740 517788 440804 517852
rect 309732 517652 309796 517716
rect 313964 517652 314028 517716
rect 325556 517652 325620 517716
rect 330340 517652 330404 517716
rect 333836 517652 333900 517716
rect 336044 517652 336108 517716
rect 338436 517652 338500 517716
rect 339540 517712 339604 517716
rect 339540 517656 339554 517712
rect 339554 517656 339604 517712
rect 339540 517652 339604 517656
rect 343404 517652 343468 517716
rect 344324 517712 344388 517716
rect 344324 517656 344338 517712
rect 344338 517656 344388 517712
rect 344324 517652 344388 517656
rect 345796 517652 345860 517716
rect 347268 517652 347332 517716
rect 348924 517712 348988 517716
rect 348924 517656 348974 517712
rect 348974 517656 348988 517712
rect 348924 517652 348988 517656
rect 433012 517652 433076 517716
rect 433932 517652 433996 517716
rect 435772 517652 435836 517716
rect 436140 517652 436204 517716
rect 436876 517652 436940 517716
rect 437980 517652 438044 517716
rect 439636 517652 439700 517716
rect 444972 517652 445036 517716
rect 453252 517652 453316 517716
rect 460244 517652 460308 517716
rect 468340 517652 468404 517716
rect 307340 517516 307404 517580
rect 308628 517516 308692 517580
rect 310284 517576 310348 517580
rect 310284 517520 310298 517576
rect 310298 517520 310348 517576
rect 310284 517516 310348 517520
rect 311572 517516 311636 517580
rect 326660 517516 326724 517580
rect 329052 517516 329116 517580
rect 337332 517516 337396 517580
rect 340644 517516 340708 517580
rect 341932 517516 341996 517580
rect 348372 517516 348436 517580
rect 438348 517516 438412 517580
rect 438716 517576 438780 517580
rect 438716 517520 438766 517576
rect 438766 517520 438780 517576
rect 438716 517516 438780 517520
rect 440004 517516 440068 517580
rect 441476 517576 441540 517580
rect 441476 517520 441526 517576
rect 441526 517520 441540 517576
rect 441476 517516 441540 517520
rect 442764 517516 442828 517580
rect 443868 517516 443932 517580
rect 445524 517576 445588 517580
rect 445524 517520 445574 517576
rect 445574 517520 445588 517576
rect 445524 517516 445588 517520
rect 446996 517576 447060 517580
rect 446996 517520 447046 517576
rect 447046 517520 447060 517576
rect 446996 517516 447060 517520
rect 448284 517516 448348 517580
rect 449756 517576 449820 517580
rect 449756 517520 449806 517576
rect 449806 517520 449820 517576
rect 449756 517516 449820 517520
rect 450860 517516 450924 517580
rect 451964 517516 452028 517580
rect 453804 517576 453868 517580
rect 453804 517520 453854 517576
rect 453854 517520 453868 517576
rect 453804 517516 453868 517520
rect 455276 517576 455340 517580
rect 455276 517520 455326 517576
rect 455326 517520 455340 517576
rect 455276 517516 455340 517520
rect 456380 517516 456444 517580
rect 457852 517516 457916 517580
rect 459140 517516 459204 517580
rect 460796 517576 460860 517580
rect 460796 517520 460810 517576
rect 460810 517520 460860 517576
rect 460796 517516 460860 517520
rect 462084 517516 462148 517580
rect 463556 517576 463620 517580
rect 463556 517520 463606 517576
rect 463606 517520 463620 517576
rect 463556 517516 463620 517520
rect 464844 517516 464908 517580
rect 466132 517516 466196 517580
rect 467236 517516 467300 517580
rect 469076 517576 469140 517580
rect 469076 517520 469090 517576
rect 469090 517520 469140 517576
rect 469076 517516 469140 517520
rect 519124 509084 519188 509148
rect 519860 509084 519924 509148
rect 519124 499564 519188 499628
rect 519860 499564 519924 499628
rect 519124 489772 519188 489836
rect 519860 489772 519924 489836
rect 357388 479980 357452 480044
rect 376708 479980 376772 480044
rect 67588 479844 67652 479908
rect 434668 479708 434732 479772
rect 67588 479572 67652 479636
rect 106228 479572 106292 479636
rect 77524 479436 77588 479500
rect 86908 479436 86972 479500
rect 96476 479436 96540 479500
rect 77340 479300 77404 479364
rect 86908 479164 86972 479228
rect 96476 479164 96540 479228
rect 106228 479164 106292 479228
rect 269068 479300 269132 479364
rect 318748 479572 318812 479636
rect 318748 479300 318812 479364
rect 376708 479572 376772 479636
rect 357388 479300 357452 479364
rect 434668 479436 434732 479500
rect 511948 479572 512012 479636
rect 519124 479572 519188 479636
rect 519860 479572 519924 479636
rect 511948 479300 512012 479364
rect 519860 479300 519924 479364
rect 269068 479028 269132 479092
rect 522804 476852 522868 476916
rect 520412 476172 520476 476236
rect 520412 476036 520476 476100
rect 519308 475764 519372 475828
rect 519492 475764 519556 475828
rect 519676 475764 519740 475828
rect 519860 475764 519924 475828
rect 519308 475492 519372 475556
rect 519492 475492 519556 475556
rect 519676 475492 519740 475556
rect 519860 475492 519924 475556
rect 521700 474676 521764 474740
rect 520228 472636 520292 472700
rect 521884 470460 521948 470524
rect 519308 468692 519372 468756
rect 521332 468692 521396 468756
rect 519492 468556 519556 468620
rect 521148 468556 521212 468620
rect 522068 468420 522132 468484
rect 519860 466516 519924 466580
rect 519676 466380 519740 466444
rect 520412 466244 520476 466308
rect 519676 465972 519740 466036
rect 519860 465836 519924 465900
rect 519492 465564 519556 465628
rect 521148 465564 521212 465628
rect 519308 465428 519372 465492
rect 521332 465428 521396 465492
rect 522252 464204 522316 464268
rect 522436 462028 522500 462092
rect 522620 457812 522684 457876
rect 519492 452644 519556 452708
rect 519676 452644 519740 452708
rect 519860 452644 519924 452708
rect 519492 452372 519556 452436
rect 519676 452372 519740 452436
rect 519860 452372 519924 452436
rect 520044 437684 520108 437748
rect 521148 437684 521212 437748
rect 520044 437548 520108 437612
rect 520044 435236 520108 435300
rect 520044 435100 520108 435164
rect 521148 435100 521212 435164
rect 520044 429796 520108 429860
rect 521148 429796 521212 429860
rect 519676 429660 519740 429724
rect 520044 429660 520108 429724
rect 520044 428028 520108 428092
rect 519676 427892 519740 427956
rect 520044 425036 520108 425100
rect 521148 425036 521212 425100
rect 519308 415516 519372 415580
rect 519492 415244 519556 415308
rect 519308 414972 519372 415036
rect 519860 415244 519924 415308
rect 519860 414972 519924 415036
rect 519308 409124 519372 409188
rect 519676 408716 519740 408780
rect 519676 408308 519740 408372
rect 519308 406948 519372 407012
rect 520044 406948 520108 407012
rect 519492 406268 519556 406332
rect 519308 406132 519372 406196
rect 519492 406132 519556 406196
rect 519308 405996 519372 406060
rect 519676 399468 519740 399532
rect 520964 396748 521028 396812
rect 519308 396340 519372 396404
rect 519308 395524 519372 395588
rect 519492 395252 519556 395316
rect 519308 393348 519372 393412
rect 519676 393348 519740 393412
rect 519308 390628 519372 390692
rect 520780 390492 520844 390556
rect 519676 388860 519740 388924
rect 519860 386004 519924 386068
rect 520596 384100 520660 384164
rect 519308 382196 519372 382260
rect 522804 237084 522868 237148
rect 336412 220764 336476 220828
rect 329420 212528 329484 212532
rect 329420 212472 329434 212528
rect 329434 212472 329484 212528
rect 329420 212468 329484 212472
rect 357388 203960 357452 203964
rect 448284 204172 448348 204236
rect 449388 204172 449452 204236
rect 451780 204172 451844 204236
rect 453252 204232 453316 204236
rect 453252 204176 453302 204232
rect 453302 204176 453316 204232
rect 453252 204172 453316 204176
rect 454172 204172 454236 204236
rect 456380 204172 456444 204236
rect 468156 204172 468220 204236
rect 470364 204172 470428 204236
rect 484348 204232 484412 204236
rect 484348 204176 484398 204232
rect 484398 204176 484412 204232
rect 484348 204172 484412 204176
rect 449572 204036 449636 204100
rect 450860 204096 450924 204100
rect 450860 204040 450910 204096
rect 450910 204040 450924 204096
rect 450860 204036 450924 204040
rect 452148 204036 452212 204100
rect 454540 204036 454604 204100
rect 456564 204036 456628 204100
rect 464476 204036 464540 204100
rect 465764 204036 465828 204100
rect 469260 204036 469324 204100
rect 476068 204036 476132 204100
rect 477540 204096 477604 204100
rect 477540 204040 477554 204096
rect 477554 204040 477604 204096
rect 477540 204036 477604 204040
rect 483428 204036 483492 204100
rect 486372 204036 486436 204100
rect 357388 203904 357438 203960
rect 357438 203904 357452 203960
rect 357388 203900 357452 203904
rect 360516 203900 360580 203964
rect 457484 203900 457548 203964
rect 460060 203900 460124 203964
rect 490236 203960 490300 203964
rect 490236 203904 490250 203960
rect 490250 203904 490300 203960
rect 490236 203900 490300 203904
rect 361620 203764 361684 203828
rect 485820 203764 485884 203828
rect 330892 203688 330956 203692
rect 330892 203632 330942 203688
rect 330942 203632 330956 203688
rect 330892 203628 330956 203632
rect 341012 203688 341076 203692
rect 341012 203632 341026 203688
rect 341026 203632 341076 203688
rect 341012 203628 341076 203632
rect 342852 203628 342916 203692
rect 347820 203688 347884 203692
rect 347820 203632 347834 203688
rect 347834 203632 347884 203688
rect 347820 203628 347884 203632
rect 349108 203688 349172 203692
rect 349108 203632 349158 203688
rect 349158 203632 349172 203688
rect 349108 203628 349172 203632
rect 352788 203628 352852 203692
rect 487476 203628 487540 203692
rect 340092 203552 340156 203556
rect 340092 203496 340106 203552
rect 340106 203496 340156 203552
rect 340092 203492 340156 203496
rect 342300 203552 342364 203556
rect 342300 203496 342314 203552
rect 342314 203496 342364 203552
rect 342300 203492 342364 203496
rect 343588 203552 343652 203556
rect 343588 203496 343638 203552
rect 343638 203496 343652 203552
rect 343588 203492 343652 203496
rect 354812 203492 354876 203556
rect 329604 203356 329668 203420
rect 330708 203356 330772 203420
rect 334204 203356 334268 203420
rect 336964 203356 337028 203420
rect 342484 203356 342548 203420
rect 362908 203356 362972 203420
rect 364380 203416 364444 203420
rect 364380 203360 364394 203416
rect 364394 203360 364444 203416
rect 364380 203356 364444 203360
rect 367508 203356 367572 203420
rect 474228 203492 474292 203556
rect 480668 203552 480732 203556
rect 480668 203496 480682 203552
rect 480682 203496 480732 203552
rect 328132 203220 328196 203284
rect 331628 203220 331692 203284
rect 332916 203220 332980 203284
rect 335124 203220 335188 203284
rect 338436 203220 338500 203284
rect 339724 203220 339788 203284
rect 346532 203220 346596 203284
rect 349844 203220 349908 203284
rect 356100 203280 356164 203284
rect 356100 203224 356114 203280
rect 356114 203224 356164 203280
rect 356100 203220 356164 203224
rect 366956 203280 367020 203284
rect 366956 203224 366970 203280
rect 366970 203224 367020 203280
rect 366956 203220 367020 203224
rect 368612 203220 368676 203284
rect 371004 203220 371068 203284
rect 456012 203356 456076 203420
rect 462268 203356 462332 203420
rect 464660 203416 464724 203420
rect 464660 203360 464710 203416
rect 464710 203360 464724 203416
rect 464660 203356 464724 203360
rect 469444 203416 469508 203420
rect 469444 203360 469494 203416
rect 469494 203360 469508 203416
rect 469444 203356 469508 203360
rect 478092 203356 478156 203420
rect 479196 203356 479260 203420
rect 480668 203492 480732 203496
rect 484532 203492 484596 203556
rect 488580 203356 488644 203420
rect 458772 203220 458836 203284
rect 460980 203220 461044 203284
rect 463188 203220 463252 203284
rect 467052 203220 467116 203284
rect 471100 203220 471164 203284
rect 471652 203220 471716 203284
rect 472756 203220 472820 203284
rect 472940 203280 473004 203284
rect 472940 203224 472954 203280
rect 472954 203224 473004 203280
rect 472940 203220 473004 203224
rect 473676 203220 473740 203284
rect 474964 203220 475028 203284
rect 477724 203220 477788 203284
rect 479932 203220 479996 203284
rect 482140 203220 482204 203284
rect 328316 203144 328380 203148
rect 328316 203088 328330 203144
rect 328330 203088 328380 203144
rect 328316 203084 328380 203088
rect 332364 203144 332428 203148
rect 332364 203088 332414 203144
rect 332414 203088 332428 203144
rect 332364 203084 332428 203088
rect 333652 203084 333716 203148
rect 336596 203144 336660 203148
rect 336596 203088 336610 203144
rect 336610 203088 336660 203144
rect 336596 203084 336660 203088
rect 343956 203084 344020 203148
rect 345244 203084 345308 203148
rect 351132 203144 351196 203148
rect 351132 203088 351146 203144
rect 351146 203088 351196 203144
rect 351132 203084 351196 203088
rect 357756 203084 357820 203148
rect 334756 202948 334820 203012
rect 336044 202948 336108 203012
rect 337884 203008 337948 203012
rect 337884 202952 337934 203008
rect 337934 202952 337948 203008
rect 337884 202948 337948 202952
rect 339172 203008 339236 203012
rect 339172 202952 339222 203008
rect 339222 202952 339236 203008
rect 339172 202948 339236 202952
rect 341380 203008 341444 203012
rect 341380 202952 341394 203008
rect 341394 202952 341444 203008
rect 341380 202948 341444 202952
rect 344876 203008 344940 203012
rect 344876 202952 344926 203008
rect 344926 202952 344940 203008
rect 344876 202948 344940 202952
rect 345980 203008 346044 203012
rect 345980 202952 345994 203008
rect 345994 202952 346044 203008
rect 345980 202948 346044 202952
rect 347084 203008 347148 203012
rect 347084 202952 347098 203008
rect 347098 202952 347148 203008
rect 347084 202948 347148 202952
rect 348372 203008 348436 203012
rect 348372 202952 348422 203008
rect 348422 202952 348436 203008
rect 348372 202948 348436 202952
rect 349476 203008 349540 203012
rect 349476 202952 349490 203008
rect 349490 202952 349540 203008
rect 349476 202948 349540 202952
rect 350948 202948 351012 203012
rect 351684 203008 351748 203012
rect 351684 202952 351698 203008
rect 351698 202952 351748 203008
rect 351684 202948 351748 202952
rect 352972 203008 353036 203012
rect 352972 202952 353022 203008
rect 353022 202952 353036 203008
rect 352972 202948 353036 202952
rect 353340 203008 353404 203012
rect 353340 202952 353354 203008
rect 353354 202952 353404 203008
rect 353340 202948 353404 202952
rect 354444 202948 354508 203012
rect 355548 203008 355612 203012
rect 355548 202952 355598 203008
rect 355598 202952 355612 203008
rect 355548 202948 355612 202952
rect 356468 203008 356532 203012
rect 356468 202952 356482 203008
rect 356482 202952 356532 203008
rect 356468 202948 356532 202952
rect 357940 202948 358004 203012
rect 358676 203008 358740 203012
rect 358676 202952 358690 203008
rect 358690 202952 358740 203008
rect 358676 202948 358740 202952
rect 359228 202948 359292 203012
rect 359964 203008 360028 203012
rect 359964 202952 360014 203008
rect 360014 202952 360028 203008
rect 359964 202948 360028 202952
rect 361252 203008 361316 203012
rect 361252 202952 361302 203008
rect 361302 202952 361316 203008
rect 361252 202948 361316 202952
rect 362724 202948 362788 203012
rect 363460 203008 363524 203012
rect 363460 202952 363474 203008
rect 363474 202952 363524 203008
rect 363460 202948 363524 202952
rect 364932 202948 364996 203012
rect 366404 203084 366468 203148
rect 373396 203084 373460 203148
rect 492812 203084 492876 203148
rect 450676 202948 450740 203012
rect 452884 202948 452948 203012
rect 455276 203008 455340 203012
rect 455276 202952 455326 203008
rect 455326 202952 455340 203008
rect 455276 202948 455340 202952
rect 457852 203008 457916 203012
rect 457852 202952 457902 203008
rect 457902 202952 457916 203008
rect 457852 202948 457916 202952
rect 458956 202948 459020 203012
rect 460612 203008 460676 203012
rect 460612 202952 460662 203008
rect 460662 202952 460676 203008
rect 460612 202948 460676 202952
rect 461532 203008 461596 203012
rect 461532 202952 461546 203008
rect 461546 202952 461596 203008
rect 461532 202948 461596 202952
rect 462452 203008 462516 203012
rect 462452 202952 462466 203008
rect 462466 202952 462516 203008
rect 462452 202948 462516 202952
rect 463556 202948 463620 203012
rect 465948 203008 466012 203012
rect 465948 202952 465962 203008
rect 465962 202952 466012 203008
rect 465948 202948 466012 202952
rect 467236 203008 467300 203012
rect 467236 202952 467250 203008
rect 467250 202952 467300 203008
rect 467236 202948 467300 202952
rect 468524 203008 468588 203012
rect 468524 202952 468538 203008
rect 468538 202952 468588 203008
rect 468524 202948 468588 202952
rect 471836 203008 471900 203012
rect 471836 202952 471850 203008
rect 471850 202952 471900 203008
rect 471836 202948 471900 202952
rect 475516 202948 475580 203012
rect 476436 202948 476500 203012
rect 478644 202948 478708 203012
rect 481036 202948 481100 203012
rect 481772 202948 481836 203012
rect 483060 203008 483124 203012
rect 483060 202952 483074 203008
rect 483074 202952 483124 203008
rect 483060 202948 483124 202952
rect 342300 201724 342364 201788
rect 342276 201452 342340 201516
rect 448384 201376 448448 201380
rect 448384 201320 448426 201376
rect 448426 201320 448448 201376
rect 448384 201316 448448 201320
rect 522620 200772 522684 200836
rect 522436 200636 522500 200700
rect 303660 109032 303724 109036
rect 303660 108976 303674 109032
rect 303674 108976 303724 109032
rect 303660 108972 303724 108976
rect 308076 108972 308140 109036
rect 424180 109032 424244 109036
rect 424180 108976 424230 109032
rect 424230 108976 424244 109032
rect 424180 108972 424244 108976
rect 428044 108972 428108 109036
rect 520412 108836 520476 108900
rect 522252 93740 522316 93804
rect 522068 80004 522132 80068
rect 520228 64772 520292 64836
rect 521884 50900 521948 50964
rect 521700 35804 521764 35868
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 67587 479908 67653 479909
rect 67587 479844 67588 479908
rect 67652 479844 67653 479908
rect 67587 479843 67653 479844
rect 67590 479637 67650 479843
rect 67587 479636 67653 479637
rect 67587 479572 67588 479636
rect 67652 479572 67653 479636
rect 67587 479571 67653 479572
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 77523 479500 77589 479501
rect 77523 479436 77524 479500
rect 77588 479436 77589 479500
rect 77523 479435 77589 479436
rect 77339 479364 77405 479365
rect 77339 479300 77340 479364
rect 77404 479300 77405 479364
rect 77339 479299 77405 479300
rect 77342 479090 77402 479299
rect 77526 479090 77586 479435
rect 77342 479030 77586 479090
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 86907 479500 86973 479501
rect 86907 479436 86908 479500
rect 86972 479436 86973 479500
rect 86907 479435 86973 479436
rect 86910 479229 86970 479435
rect 86907 479228 86973 479229
rect 86907 479164 86908 479228
rect 86972 479164 86973 479228
rect 86907 479163 86973 479164
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 96475 479500 96541 479501
rect 96475 479436 96476 479500
rect 96540 479436 96541 479500
rect 96475 479435 96541 479436
rect 96478 479229 96538 479435
rect 96475 479228 96541 479229
rect 96475 479164 96476 479228
rect 96540 479164 96541 479228
rect 96475 479163 96541 479164
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 106227 479636 106293 479637
rect 106227 479572 106228 479636
rect 106292 479572 106293 479636
rect 106227 479571 106293 479572
rect 106230 479229 106290 479571
rect 106227 479228 106293 479229
rect 106227 479164 106228 479228
rect 106292 479164 106293 479228
rect 106227 479163 106293 479164
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 269067 479364 269133 479365
rect 269067 479300 269068 479364
rect 269132 479300 269133 479364
rect 269067 479299 269133 479300
rect 269070 479093 269130 479299
rect 269067 479092 269133 479093
rect 269067 479028 269068 479092
rect 269132 479028 269133 479092
rect 269067 479027 269133 479028
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 483000 278604 495098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 483000 282204 498698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 483000 289404 505898
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 483000 293004 509498
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 614247 300204 624698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 614247 307404 631898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 614247 311004 635498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 614247 314604 639098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 614247 318204 642698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614247 325404 649898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 614247 329004 617498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 614247 332604 621098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 614247 336204 624698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 614247 343404 631898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 614247 347004 635498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 614247 350604 639098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 614247 354204 642698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614247 361404 649898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 614247 365004 617498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 614247 368604 621098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 614247 372204 624698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 614247 379404 631898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 373579 612780 373645 612781
rect 373579 612716 373580 612780
rect 373644 612716 373645 612780
rect 373579 612715 373645 612716
rect 369163 611012 369229 611013
rect 369163 611010 369164 611012
rect 368608 610950 369164 611010
rect 369163 610948 369164 610950
rect 369228 610948 369229 611012
rect 369163 610947 369229 610948
rect 373027 611012 373093 611013
rect 373027 610948 373028 611012
rect 373092 611010 373093 611012
rect 373582 611010 373642 612715
rect 373092 610950 373642 611010
rect 373092 610948 373093 610950
rect 373027 610947 373093 610948
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 376938 596454 377262 596476
rect 376938 596218 376982 596454
rect 377218 596218 377262 596454
rect 376938 596134 377262 596218
rect 376938 595898 376982 596134
rect 377218 595898 377262 596134
rect 376938 595876 377262 595898
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 376494 578454 376814 578476
rect 376494 578218 376536 578454
rect 376772 578218 376814 578454
rect 376494 578134 376814 578218
rect 376494 577898 376536 578134
rect 376772 577898 376814 578134
rect 376494 577876 376814 577898
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 376938 560454 377262 560476
rect 376938 560218 376982 560454
rect 377218 560218 377262 560454
rect 376938 560134 377262 560218
rect 376938 559898 376982 560134
rect 377218 559898 377262 560134
rect 376938 559876 377262 559898
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 376494 542454 376814 542476
rect 376494 542218 376536 542454
rect 376772 542218 376814 542454
rect 376494 542134 376814 542218
rect 376494 541898 376536 542134
rect 376772 541898 376814 542134
rect 376494 541876 376814 541898
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 376938 524454 377262 524476
rect 376938 524218 376982 524454
rect 377218 524218 377262 524454
rect 376938 524134 377262 524218
rect 376938 523898 376982 524134
rect 377218 523898 377262 524134
rect 376938 523876 377262 523898
rect 314702 520510 315008 520570
rect 316300 520510 316602 520570
rect 319804 520510 320098 520570
rect 303662 520170 303833 520230
rect 306832 520170 307402 520230
rect 308000 520170 308690 520230
rect 309168 520170 309794 520230
rect 303662 518261 303722 520170
rect 303659 518260 303725 518261
rect 303659 518196 303660 518260
rect 303724 518196 303725 518260
rect 303659 518195 303725 518196
rect 307342 517581 307402 520170
rect 308630 517581 308690 520170
rect 309734 517717 309794 520170
rect 309731 517716 309797 517717
rect 309731 517652 309732 517716
rect 309796 517652 309797 517716
rect 309731 517651 309797 517652
rect 310286 517581 310346 520230
rect 311474 519890 311534 520200
rect 312494 520170 312672 520230
rect 311474 519830 311634 519890
rect 311574 517581 311634 519830
rect 312494 518397 312554 520170
rect 312766 519890 312826 520200
rect 312678 519830 312826 519890
rect 312491 518396 312557 518397
rect 312491 518332 312492 518396
rect 312556 518332 312557 518396
rect 312491 518331 312557 518332
rect 312678 517989 312738 519830
rect 313782 518805 313842 520230
rect 313964 520170 314026 520230
rect 313779 518804 313845 518805
rect 313779 518740 313780 518804
rect 313844 518740 313845 518804
rect 313779 518739 313845 518740
rect 312675 517988 312741 517989
rect 312675 517924 312676 517988
rect 312740 517924 312741 517988
rect 312675 517923 312741 517924
rect 313966 517717 314026 520170
rect 314702 518669 314762 520510
rect 315102 519890 315162 520200
rect 315070 519830 315162 519890
rect 316146 519890 316206 520200
rect 316146 519830 316234 519890
rect 314699 518668 314765 518669
rect 314699 518604 314700 518668
rect 314764 518604 314765 518668
rect 314699 518603 314765 518604
rect 315070 518261 315130 519830
rect 316174 518805 316234 519830
rect 316171 518804 316237 518805
rect 316171 518740 316172 518804
rect 316236 518740 316237 518804
rect 316171 518739 316237 518740
rect 316542 518533 316602 520510
rect 317278 520170 317344 520230
rect 317278 518669 317338 520170
rect 317275 518668 317341 518669
rect 317275 518604 317276 518668
rect 317340 518604 317341 518668
rect 317275 518603 317341 518604
rect 316539 518532 316605 518533
rect 316539 518468 316540 518532
rect 316604 518468 316605 518532
rect 316539 518467 316605 518468
rect 317462 518397 317522 520230
rect 318482 519890 318542 520200
rect 318636 520170 318810 520230
rect 318482 519830 318626 519890
rect 318566 518805 318626 519830
rect 318563 518804 318629 518805
rect 318563 518740 318564 518804
rect 318628 518740 318629 518804
rect 318563 518739 318629 518740
rect 318563 518532 318629 518533
rect 318563 518468 318564 518532
rect 318628 518530 318629 518532
rect 318750 518530 318810 520170
rect 319650 519890 319710 520200
rect 319650 519830 319730 519890
rect 319670 518669 319730 519830
rect 319667 518668 319733 518669
rect 319667 518604 319668 518668
rect 319732 518604 319733 518668
rect 319667 518603 319733 518604
rect 318628 518470 318810 518530
rect 318628 518468 318629 518470
rect 318563 518467 318629 518468
rect 317459 518396 317525 518397
rect 317459 518332 317460 518396
rect 317524 518332 317525 518396
rect 317459 518331 317525 518332
rect 315067 518260 315133 518261
rect 315067 518196 315068 518260
rect 315132 518196 315133 518260
rect 315067 518195 315133 518196
rect 320038 518125 320098 520510
rect 321694 520510 322016 520570
rect 323308 520510 323594 520570
rect 320774 520170 320848 520230
rect 320774 518397 320834 520170
rect 320771 518396 320837 518397
rect 320771 518332 320772 518396
rect 320836 518332 320837 518396
rect 320771 518331 320837 518332
rect 320035 518124 320101 518125
rect 320035 518060 320036 518124
rect 320100 518060 320101 518124
rect 320035 518059 320101 518060
rect 320958 517853 321018 520230
rect 321694 518805 321754 520510
rect 322110 519890 322170 520200
rect 322062 519830 322170 519890
rect 323154 519890 323214 520200
rect 323154 519830 323226 519890
rect 321691 518804 321757 518805
rect 321691 518740 321692 518804
rect 321756 518740 321757 518804
rect 321691 518739 321757 518740
rect 322062 518125 322122 519830
rect 323166 518805 323226 519830
rect 323163 518804 323229 518805
rect 323163 518740 323164 518804
rect 323228 518740 323229 518804
rect 323163 518739 323229 518740
rect 323534 518261 323594 520510
rect 325190 520510 325520 520570
rect 338070 520510 338368 520570
rect 341566 520510 341872 520570
rect 343164 520510 343466 520570
rect 324270 520170 324352 520230
rect 324270 518669 324330 520170
rect 324454 518805 324514 520230
rect 325190 518805 325250 520510
rect 325614 519890 325674 520200
rect 325558 519830 325674 519890
rect 326478 520170 326688 520230
rect 324451 518804 324517 518805
rect 324451 518740 324452 518804
rect 324516 518740 324517 518804
rect 324451 518739 324517 518740
rect 325187 518804 325253 518805
rect 325187 518740 325188 518804
rect 325252 518740 325253 518804
rect 325187 518739 325253 518740
rect 324267 518668 324333 518669
rect 324267 518604 324268 518668
rect 324332 518604 324333 518668
rect 324267 518603 324333 518604
rect 323531 518260 323597 518261
rect 323531 518196 323532 518260
rect 323596 518196 323597 518260
rect 323531 518195 323597 518196
rect 322059 518124 322125 518125
rect 322059 518060 322060 518124
rect 322124 518060 322125 518124
rect 322059 518059 322125 518060
rect 320955 517852 321021 517853
rect 320955 517788 320956 517852
rect 321020 517788 321021 517852
rect 320955 517787 321021 517788
rect 325558 517717 325618 519830
rect 326478 518805 326538 520170
rect 326782 519890 326842 520200
rect 326662 519830 326842 519890
rect 327214 520170 327856 520230
rect 326475 518804 326541 518805
rect 326475 518740 326476 518804
rect 326540 518740 326541 518804
rect 326475 518739 326541 518740
rect 313963 517716 314029 517717
rect 313963 517652 313964 517716
rect 314028 517652 314029 517716
rect 313963 517651 314029 517652
rect 325555 517716 325621 517717
rect 325555 517652 325556 517716
rect 325620 517652 325621 517716
rect 325555 517651 325621 517652
rect 326662 517581 326722 519830
rect 327214 518805 327274 520170
rect 327211 518804 327277 518805
rect 327211 518740 327212 518804
rect 327276 518740 327277 518804
rect 327211 518739 327277 518740
rect 327950 518533 328010 520200
rect 328870 520170 329024 520230
rect 328870 518805 328930 520170
rect 329118 519890 329178 520200
rect 329054 519830 329178 519890
rect 328867 518804 328933 518805
rect 328867 518740 328868 518804
rect 328932 518740 328933 518804
rect 328867 518739 328933 518740
rect 327947 518532 328013 518533
rect 327947 518468 327948 518532
rect 328012 518468 328013 518532
rect 327947 518467 328013 518468
rect 329054 517581 329114 519830
rect 330158 518805 330218 520230
rect 330316 520170 330402 520230
rect 330155 518804 330221 518805
rect 330155 518740 330156 518804
rect 330220 518740 330221 518804
rect 330155 518739 330221 518740
rect 330342 517717 330402 520170
rect 331308 519890 331368 520230
rect 331454 519890 331514 520200
rect 331262 519830 331368 519890
rect 331446 519830 331514 519890
rect 332366 520170 332528 520230
rect 331262 518669 331322 519830
rect 331259 518668 331325 518669
rect 331259 518604 331260 518668
rect 331324 518604 331325 518668
rect 331259 518603 331325 518604
rect 331446 517989 331506 519830
rect 332366 518805 332426 520170
rect 332622 519890 332682 520200
rect 333470 520170 333696 520230
rect 333820 520170 333898 520230
rect 332622 519830 332794 519890
rect 332363 518804 332429 518805
rect 332363 518740 332364 518804
rect 332428 518740 332429 518804
rect 332363 518739 332429 518740
rect 332734 517989 332794 519830
rect 333470 518533 333530 520170
rect 333467 518532 333533 518533
rect 333467 518468 333468 518532
rect 333532 518468 333533 518532
rect 333467 518467 333533 518468
rect 331443 517988 331509 517989
rect 331443 517924 331444 517988
rect 331508 517924 331509 517988
rect 331443 517923 331509 517924
rect 332731 517988 332797 517989
rect 332731 517924 332732 517988
rect 332796 517924 332797 517988
rect 332731 517923 332797 517924
rect 333838 517717 333898 520170
rect 334206 520170 334864 520230
rect 334206 518533 334266 520170
rect 334958 519890 335018 520200
rect 334942 519830 335018 519890
rect 335494 520170 336032 520230
rect 334203 518532 334269 518533
rect 334203 518468 334204 518532
rect 334268 518468 334269 518532
rect 334203 518467 334269 518468
rect 334942 517853 335002 519830
rect 335494 518805 335554 520170
rect 336126 519890 336186 520200
rect 336046 519830 336186 519890
rect 335491 518804 335557 518805
rect 335491 518740 335492 518804
rect 335556 518740 335557 518804
rect 335491 518739 335557 518740
rect 334939 517852 335005 517853
rect 334939 517788 334940 517852
rect 335004 517788 335005 517852
rect 334939 517787 335005 517788
rect 336046 517717 336106 519830
rect 337150 518805 337210 520230
rect 337324 520170 337394 520230
rect 337147 518804 337213 518805
rect 337147 518740 337148 518804
rect 337212 518740 337213 518804
rect 337147 518739 337213 518740
rect 330339 517716 330405 517717
rect 330339 517652 330340 517716
rect 330404 517652 330405 517716
rect 330339 517651 330405 517652
rect 333835 517716 333901 517717
rect 333835 517652 333836 517716
rect 333900 517652 333901 517716
rect 333835 517651 333901 517652
rect 336043 517716 336109 517717
rect 336043 517652 336044 517716
rect 336108 517652 336109 517716
rect 336043 517651 336109 517652
rect 337334 517581 337394 520170
rect 338070 518669 338130 520510
rect 338462 519890 338522 520200
rect 338438 519830 338522 519890
rect 339358 520170 339536 520230
rect 338067 518668 338133 518669
rect 338067 518604 338068 518668
rect 338132 518604 338133 518668
rect 338067 518603 338133 518604
rect 338438 517717 338498 519830
rect 339358 518805 339418 520170
rect 339630 519890 339690 520200
rect 339542 519830 339690 519890
rect 340462 520170 340704 520230
rect 339355 518804 339421 518805
rect 339355 518740 339356 518804
rect 339420 518740 339421 518804
rect 339355 518739 339421 518740
rect 339542 517717 339602 519830
rect 340462 518805 340522 520170
rect 340798 519890 340858 520200
rect 340646 519830 340858 519890
rect 340459 518804 340525 518805
rect 340459 518740 340460 518804
rect 340524 518740 340525 518804
rect 340459 518739 340525 518740
rect 338435 517716 338501 517717
rect 338435 517652 338436 517716
rect 338500 517652 338501 517716
rect 338435 517651 338501 517652
rect 339539 517716 339605 517717
rect 339539 517652 339540 517716
rect 339604 517652 339605 517716
rect 339539 517651 339605 517652
rect 340646 517581 340706 519830
rect 341566 518805 341626 520510
rect 341966 519890 342026 520200
rect 341934 519830 342026 519890
rect 343010 519890 343070 520200
rect 343010 519830 343098 519890
rect 341563 518804 341629 518805
rect 341563 518740 341564 518804
rect 341628 518740 341629 518804
rect 341563 518739 341629 518740
rect 341934 517581 341994 519830
rect 343038 518805 343098 519830
rect 343035 518804 343101 518805
rect 343035 518740 343036 518804
rect 343100 518740 343101 518804
rect 343035 518739 343101 518740
rect 343406 517717 343466 520510
rect 348558 520510 348880 520570
rect 344142 520170 344208 520230
rect 344142 518805 344202 520170
rect 344139 518804 344205 518805
rect 344139 518740 344140 518804
rect 344204 518740 344205 518804
rect 344139 518739 344205 518740
rect 344326 517717 344386 520230
rect 345346 519890 345406 520200
rect 345500 520170 345858 520230
rect 345346 519830 345490 519890
rect 345430 518805 345490 519830
rect 345427 518804 345493 518805
rect 345427 518740 345428 518804
rect 345492 518740 345493 518804
rect 345427 518739 345493 518740
rect 345798 517717 345858 520170
rect 346514 519890 346574 520200
rect 346668 520170 347330 520230
rect 346514 519830 346594 519890
rect 346534 518805 346594 519830
rect 346531 518804 346597 518805
rect 346531 518740 346532 518804
rect 346596 518740 346597 518804
rect 346531 518739 346597 518740
rect 347270 517717 347330 520170
rect 347638 520170 347712 520230
rect 347836 520170 348434 520230
rect 347638 518805 347698 520170
rect 347635 518804 347701 518805
rect 347635 518740 347636 518804
rect 347700 518740 347701 518804
rect 347635 518739 347701 518740
rect 343403 517716 343469 517717
rect 343403 517652 343404 517716
rect 343468 517652 343469 517716
rect 343403 517651 343469 517652
rect 344323 517716 344389 517717
rect 344323 517652 344324 517716
rect 344388 517652 344389 517716
rect 344323 517651 344389 517652
rect 345795 517716 345861 517717
rect 345795 517652 345796 517716
rect 345860 517652 345861 517716
rect 345795 517651 345861 517652
rect 347267 517716 347333 517717
rect 347267 517652 347268 517716
rect 347332 517652 347333 517716
rect 347267 517651 347333 517652
rect 348374 517581 348434 520170
rect 348558 518805 348618 520510
rect 348974 519890 349034 520200
rect 348926 519830 349034 519890
rect 348555 518804 348621 518805
rect 348555 518740 348556 518804
rect 348620 518740 348621 518804
rect 348555 518739 348621 518740
rect 348926 517717 348986 519830
rect 348923 517716 348989 517717
rect 348923 517652 348924 517716
rect 348988 517652 348989 517716
rect 348923 517651 348989 517652
rect 307339 517580 307405 517581
rect 307339 517516 307340 517580
rect 307404 517516 307405 517580
rect 307339 517515 307405 517516
rect 308627 517580 308693 517581
rect 308627 517516 308628 517580
rect 308692 517516 308693 517580
rect 308627 517515 308693 517516
rect 310283 517580 310349 517581
rect 310283 517516 310284 517580
rect 310348 517516 310349 517580
rect 310283 517515 310349 517516
rect 311571 517580 311637 517581
rect 311571 517516 311572 517580
rect 311636 517516 311637 517580
rect 311571 517515 311637 517516
rect 326659 517580 326725 517581
rect 326659 517516 326660 517580
rect 326724 517516 326725 517580
rect 326659 517515 326725 517516
rect 329051 517580 329117 517581
rect 329051 517516 329052 517580
rect 329116 517516 329117 517580
rect 329051 517515 329117 517516
rect 337331 517580 337397 517581
rect 337331 517516 337332 517580
rect 337396 517516 337397 517580
rect 337331 517515 337397 517516
rect 340643 517580 340709 517581
rect 340643 517516 340644 517580
rect 340708 517516 340709 517580
rect 340643 517515 340709 517516
rect 341931 517580 341997 517581
rect 341931 517516 341932 517580
rect 341996 517516 341997 517580
rect 341931 517515 341997 517516
rect 348371 517580 348437 517581
rect 348371 517516 348372 517580
rect 348436 517516 348437 517580
rect 348371 517515 348437 517516
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 483000 296604 513098
rect 299604 483000 300204 517000
rect 306804 488454 307404 517000
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 483000 307404 487898
rect 310404 492054 311004 517000
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 483000 311004 491498
rect 314004 495654 314604 517000
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 483000 314604 495098
rect 317604 499254 318204 517000
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 483000 318204 498698
rect 324804 506454 325404 517000
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 483000 325404 505898
rect 328404 510054 329004 517000
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 483000 329004 509498
rect 332004 513654 332604 517000
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 483000 332604 513098
rect 335604 483000 336204 517000
rect 342804 488454 343404 517000
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 483000 343404 487898
rect 346404 492054 347004 517000
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 483000 347004 491498
rect 350004 495654 350604 517000
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 483000 350604 495098
rect 353604 499254 354204 517000
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 483000 354204 498698
rect 360804 506454 361404 517000
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 483000 361404 505898
rect 364404 510054 365004 517000
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 483000 365004 509498
rect 368004 513654 368604 517000
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 483000 368604 513098
rect 371604 483000 372204 517000
rect 378804 488454 379404 517000
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 483000 379404 487898
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 483000 383004 491498
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 483000 386604 495098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 483000 390204 498698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 483000 397404 505898
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 483000 401004 509498
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 483000 404604 513098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 483000 408204 516698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 614247 419004 635498
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 614247 422604 639098
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 614247 426204 642698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614247 433404 649898
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 614247 437004 617498
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 614247 440604 621098
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 614247 444204 624698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 614247 451404 631898
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 614247 455004 635498
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 614247 458604 639098
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 614247 462204 642698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614247 469404 649898
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 614247 473004 617498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 614247 476604 621098
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 614247 480204 624698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 614247 487404 631898
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 614247 491004 635498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 614247 494604 639098
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 614247 498204 642698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 488579 612780 488645 612781
rect 488579 612716 488580 612780
rect 488644 612716 488645 612780
rect 488579 612715 488645 612716
rect 493915 612780 493981 612781
rect 493915 612716 493916 612780
rect 493980 612716 493981 612780
rect 493915 612715 493981 612716
rect 488582 610950 488642 612715
rect 493918 611010 493978 612715
rect 493603 610950 493978 611010
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 496938 596454 497262 596476
rect 496938 596218 496982 596454
rect 497218 596218 497262 596454
rect 496938 596134 497262 596218
rect 496938 595898 496982 596134
rect 497218 595898 497262 596134
rect 496938 595876 497262 595898
rect 496494 578454 496814 578476
rect 496494 578218 496536 578454
rect 496772 578218 496814 578454
rect 496494 578134 496814 578218
rect 496494 577898 496536 578134
rect 496772 577898 496814 578134
rect 496494 577876 496814 577898
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 496938 560454 497262 560476
rect 496938 560218 496982 560454
rect 497218 560218 497262 560454
rect 496938 560134 497262 560218
rect 496938 559898 496982 560134
rect 497218 559898 497262 560134
rect 496938 559876 497262 559898
rect 496494 542454 496814 542476
rect 496494 542218 496536 542454
rect 496772 542218 496814 542454
rect 496494 542134 496814 542218
rect 496494 541898 496536 542134
rect 496772 541898 496814 542134
rect 496494 541876 496814 541898
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 496938 524454 497262 524476
rect 496938 524218 496982 524454
rect 497218 524218 497262 524454
rect 496938 524134 497262 524218
rect 496938 523898 496982 524134
rect 497218 523898 497262 524134
rect 496938 523876 497262 523898
rect 423814 518261 423874 520230
rect 426574 520170 426832 520230
rect 426574 518533 426634 520170
rect 427970 519757 428030 520200
rect 427967 519756 428033 519757
rect 427967 519692 427968 519756
rect 428032 519692 428033 519756
rect 427967 519691 428033 519692
rect 426571 518532 426637 518533
rect 426571 518468 426572 518532
rect 426636 518468 426637 518532
rect 426571 518467 426637 518468
rect 429150 518261 429210 520230
rect 429702 520170 430336 520230
rect 430806 520170 431504 520230
rect 429702 518669 429762 520170
rect 429699 518668 429765 518669
rect 429699 518604 429700 518668
rect 429764 518604 429765 518668
rect 429699 518603 429765 518604
rect 430806 518397 430866 520170
rect 432642 519890 432702 520200
rect 432796 520170 433074 520230
rect 432642 519830 432706 519890
rect 430803 518396 430869 518397
rect 430803 518332 430804 518396
rect 430868 518332 430869 518396
rect 430803 518331 430869 518332
rect 423811 518260 423877 518261
rect 423811 518196 423812 518260
rect 423876 518196 423877 518260
rect 423811 518195 423877 518196
rect 429147 518260 429213 518261
rect 429147 518196 429148 518260
rect 429212 518196 429213 518260
rect 429147 518195 429213 518196
rect 432646 517853 432706 519830
rect 432643 517852 432709 517853
rect 432643 517788 432644 517852
rect 432708 517788 432709 517852
rect 432643 517787 432709 517788
rect 433014 517717 433074 520170
rect 433750 520170 433840 520230
rect 433750 517853 433810 520170
rect 433747 517852 433813 517853
rect 433747 517788 433748 517852
rect 433812 517788 433813 517852
rect 433747 517787 433813 517788
rect 433934 517717 433994 520200
rect 434978 519890 435038 520200
rect 435132 520170 435834 520230
rect 434978 519830 435098 519890
rect 435038 518125 435098 519830
rect 435035 518124 435101 518125
rect 435035 518060 435036 518124
rect 435100 518060 435101 518124
rect 435035 518059 435101 518060
rect 435774 517717 435834 520170
rect 436142 517717 436202 520230
rect 436300 520170 436938 520230
rect 436878 517717 436938 520170
rect 437314 519890 437374 520200
rect 437468 520170 438042 520230
rect 437246 519830 437374 519890
rect 437246 517989 437306 519830
rect 437243 517988 437309 517989
rect 437243 517924 437244 517988
rect 437308 517924 437309 517988
rect 437243 517923 437309 517924
rect 437982 517717 438042 520170
rect 438350 520170 438512 520230
rect 433011 517716 433077 517717
rect 433011 517652 433012 517716
rect 433076 517652 433077 517716
rect 433011 517651 433077 517652
rect 433931 517716 433997 517717
rect 433931 517652 433932 517716
rect 433996 517652 433997 517716
rect 433931 517651 433997 517652
rect 435771 517716 435837 517717
rect 435771 517652 435772 517716
rect 435836 517652 435837 517716
rect 435771 517651 435837 517652
rect 436139 517716 436205 517717
rect 436139 517652 436140 517716
rect 436204 517652 436205 517716
rect 436139 517651 436205 517652
rect 436875 517716 436941 517717
rect 436875 517652 436876 517716
rect 436940 517652 436941 517716
rect 436875 517651 436941 517652
rect 437979 517716 438045 517717
rect 437979 517652 437980 517716
rect 438044 517652 438045 517716
rect 437979 517651 438045 517652
rect 438350 517581 438410 520170
rect 438606 519890 438666 520200
rect 438606 519830 438778 519890
rect 438718 517581 438778 519830
rect 439638 517717 439698 520230
rect 439804 520170 440066 520230
rect 439635 517716 439701 517717
rect 439635 517652 439636 517716
rect 439700 517652 439701 517716
rect 439635 517651 439701 517652
rect 440006 517581 440066 520170
rect 440818 519890 440878 520200
rect 440972 520170 441538 520230
rect 440742 519830 440878 519890
rect 440742 517853 440802 519830
rect 440739 517852 440805 517853
rect 440739 517788 440740 517852
rect 440804 517788 440805 517852
rect 440739 517787 440805 517788
rect 441478 517581 441538 520170
rect 441986 519890 442046 520200
rect 442140 520170 442826 520230
rect 441986 519830 442090 519890
rect 442030 518397 442090 519830
rect 442027 518396 442093 518397
rect 442027 518332 442028 518396
rect 442092 518332 442093 518396
rect 442027 518331 442093 518332
rect 442766 517581 442826 520170
rect 443134 518805 443194 520230
rect 443308 520170 443930 520230
rect 443131 518804 443197 518805
rect 443131 518740 443132 518804
rect 443196 518740 443197 518804
rect 443131 518739 443197 518740
rect 443870 517581 443930 520170
rect 444054 520170 444352 520230
rect 444476 520170 445034 520230
rect 444054 518397 444114 520170
rect 444051 518396 444117 518397
rect 444051 518332 444052 518396
rect 444116 518332 444117 518396
rect 444051 518331 444117 518332
rect 444974 517717 445034 520170
rect 445342 520170 445520 520230
rect 445342 518533 445402 520170
rect 445614 519890 445674 520200
rect 445526 519830 445674 519890
rect 445339 518532 445405 518533
rect 445339 518468 445340 518532
rect 445404 518468 445405 518532
rect 445339 518467 445405 518468
rect 444971 517716 445037 517717
rect 444971 517652 444972 517716
rect 445036 517652 445037 517716
rect 444971 517651 445037 517652
rect 445526 517581 445586 519830
rect 446630 518533 446690 520230
rect 446812 520170 447058 520230
rect 446627 518532 446693 518533
rect 446627 518468 446628 518532
rect 446692 518468 446693 518532
rect 446627 518467 446693 518468
rect 446998 517581 447058 520170
rect 447826 519890 447886 520200
rect 447980 520170 448346 520230
rect 447734 519830 447886 519890
rect 447734 518533 447794 519830
rect 447731 518532 447797 518533
rect 447731 518468 447732 518532
rect 447796 518468 447797 518532
rect 447731 518467 447797 518468
rect 448286 517581 448346 520170
rect 448838 520170 449024 520230
rect 449148 520170 449818 520230
rect 448838 518397 448898 520170
rect 448835 518396 448901 518397
rect 448835 518332 448836 518396
rect 448900 518332 448901 518396
rect 448835 518331 448901 518332
rect 449758 517581 449818 520170
rect 449942 520170 450192 520230
rect 450316 520170 450922 520230
rect 449942 518397 450002 520170
rect 449939 518396 450005 518397
rect 449939 518332 449940 518396
rect 450004 518332 450005 518396
rect 449939 518331 450005 518332
rect 450862 517581 450922 520170
rect 451330 519890 451390 520200
rect 451484 520170 452026 520230
rect 451230 519830 451390 519890
rect 451230 518805 451290 519830
rect 451227 518804 451293 518805
rect 451227 518740 451228 518804
rect 451292 518740 451293 518804
rect 451227 518739 451293 518740
rect 451966 517581 452026 520170
rect 452498 519890 452558 520200
rect 452652 520170 453314 520230
rect 452498 519830 452578 519890
rect 452518 518805 452578 519830
rect 452515 518804 452581 518805
rect 452515 518740 452516 518804
rect 452580 518740 452581 518804
rect 452515 518739 452581 518740
rect 453254 517717 453314 520170
rect 453622 520170 453696 520230
rect 453622 518805 453682 520170
rect 453619 518804 453685 518805
rect 453619 518740 453620 518804
rect 453684 518740 453685 518804
rect 453619 518739 453685 518740
rect 453251 517716 453317 517717
rect 453251 517652 453252 517716
rect 453316 517652 453317 517716
rect 453251 517651 453317 517652
rect 453806 517581 453866 520230
rect 454834 519890 454894 520200
rect 454988 520170 455338 520230
rect 454726 519830 454894 519890
rect 454726 518669 454786 519830
rect 454723 518668 454789 518669
rect 454723 518604 454724 518668
rect 454788 518604 454789 518668
rect 454723 518603 454789 518604
rect 455278 517581 455338 520170
rect 456002 519890 456062 520200
rect 456156 520170 456442 520230
rect 456002 519830 456074 519890
rect 456014 518669 456074 519830
rect 456011 518668 456077 518669
rect 456011 518604 456012 518668
rect 456076 518604 456077 518668
rect 456011 518603 456077 518604
rect 456382 517581 456442 520170
rect 457118 520170 457200 520230
rect 457324 520170 457914 520230
rect 457118 518669 457178 520170
rect 457115 518668 457181 518669
rect 457115 518604 457116 518668
rect 457180 518604 457181 518668
rect 457115 518603 457181 518604
rect 457854 517581 457914 520170
rect 458338 519890 458398 520200
rect 458492 520170 459202 520230
rect 458338 519830 458466 519890
rect 458406 518669 458466 519830
rect 458403 518668 458469 518669
rect 458403 518604 458404 518668
rect 458468 518604 458469 518668
rect 458403 518603 458469 518604
rect 459142 517581 459202 520170
rect 459506 519890 459566 520200
rect 459660 520170 460306 520230
rect 459506 519830 459570 519890
rect 459510 518669 459570 519830
rect 459507 518668 459573 518669
rect 459507 518604 459508 518668
rect 459572 518604 459573 518668
rect 459507 518603 459573 518604
rect 460246 517717 460306 520170
rect 460430 520170 460704 520230
rect 460430 518805 460490 520170
rect 460427 518804 460493 518805
rect 460427 518740 460428 518804
rect 460492 518740 460493 518804
rect 460427 518739 460493 518740
rect 460243 517716 460309 517717
rect 460243 517652 460244 517716
rect 460308 517652 460309 517716
rect 460243 517651 460309 517652
rect 460798 517581 460858 520200
rect 461166 520170 461872 520230
rect 461996 520170 462146 520230
rect 461166 518805 461226 520170
rect 461163 518804 461229 518805
rect 461163 518740 461164 518804
rect 461228 518740 461229 518804
rect 461163 518739 461229 518740
rect 462086 517581 462146 520170
rect 462454 520170 463040 520230
rect 463164 520170 463618 520230
rect 462454 518805 462514 520170
rect 462451 518804 462517 518805
rect 462451 518740 462452 518804
rect 462516 518740 462517 518804
rect 462451 518739 462517 518740
rect 463558 517581 463618 520170
rect 463926 520170 464208 520230
rect 464332 520170 464906 520230
rect 463926 518397 463986 520170
rect 463923 518396 463989 518397
rect 463923 518332 463924 518396
rect 463988 518332 463989 518396
rect 463923 518331 463989 518332
rect 464846 517581 464906 520170
rect 465214 520170 465376 520230
rect 465500 520170 466194 520230
rect 465214 518669 465274 520170
rect 465211 518668 465277 518669
rect 465211 518604 465212 518668
rect 465276 518604 465277 518668
rect 465211 518603 465277 518604
rect 466134 517581 466194 520170
rect 466502 518533 466562 520230
rect 466668 520170 467298 520230
rect 466499 518532 466565 518533
rect 466499 518468 466500 518532
rect 466564 518468 466565 518532
rect 466499 518467 466565 518468
rect 467238 517581 467298 520170
rect 467422 520170 467712 520230
rect 467836 520170 468402 520230
rect 467422 518669 467482 520170
rect 467419 518668 467485 518669
rect 467419 518604 467420 518668
rect 467484 518604 467485 518668
rect 467419 518603 467485 518604
rect 468342 517717 468402 520170
rect 468526 520170 468880 520230
rect 468526 518397 468586 520170
rect 468974 519890 469034 520200
rect 468974 519830 469138 519890
rect 468523 518396 468589 518397
rect 468523 518332 468524 518396
rect 468588 518332 468589 518396
rect 468523 518331 468589 518332
rect 468339 517716 468405 517717
rect 468339 517652 468340 517716
rect 468404 517652 468405 517716
rect 468339 517651 468405 517652
rect 469078 517581 469138 519830
rect 438347 517580 438413 517581
rect 438347 517516 438348 517580
rect 438412 517516 438413 517580
rect 438347 517515 438413 517516
rect 438715 517580 438781 517581
rect 438715 517516 438716 517580
rect 438780 517516 438781 517580
rect 438715 517515 438781 517516
rect 440003 517580 440069 517581
rect 440003 517516 440004 517580
rect 440068 517516 440069 517580
rect 440003 517515 440069 517516
rect 441475 517580 441541 517581
rect 441475 517516 441476 517580
rect 441540 517516 441541 517580
rect 441475 517515 441541 517516
rect 442763 517580 442829 517581
rect 442763 517516 442764 517580
rect 442828 517516 442829 517580
rect 442763 517515 442829 517516
rect 443867 517580 443933 517581
rect 443867 517516 443868 517580
rect 443932 517516 443933 517580
rect 443867 517515 443933 517516
rect 445523 517580 445589 517581
rect 445523 517516 445524 517580
rect 445588 517516 445589 517580
rect 445523 517515 445589 517516
rect 446995 517580 447061 517581
rect 446995 517516 446996 517580
rect 447060 517516 447061 517580
rect 446995 517515 447061 517516
rect 448283 517580 448349 517581
rect 448283 517516 448284 517580
rect 448348 517516 448349 517580
rect 448283 517515 448349 517516
rect 449755 517580 449821 517581
rect 449755 517516 449756 517580
rect 449820 517516 449821 517580
rect 449755 517515 449821 517516
rect 450859 517580 450925 517581
rect 450859 517516 450860 517580
rect 450924 517516 450925 517580
rect 450859 517515 450925 517516
rect 451963 517580 452029 517581
rect 451963 517516 451964 517580
rect 452028 517516 452029 517580
rect 451963 517515 452029 517516
rect 453803 517580 453869 517581
rect 453803 517516 453804 517580
rect 453868 517516 453869 517580
rect 453803 517515 453869 517516
rect 455275 517580 455341 517581
rect 455275 517516 455276 517580
rect 455340 517516 455341 517580
rect 455275 517515 455341 517516
rect 456379 517580 456445 517581
rect 456379 517516 456380 517580
rect 456444 517516 456445 517580
rect 456379 517515 456445 517516
rect 457851 517580 457917 517581
rect 457851 517516 457852 517580
rect 457916 517516 457917 517580
rect 457851 517515 457917 517516
rect 459139 517580 459205 517581
rect 459139 517516 459140 517580
rect 459204 517516 459205 517580
rect 459139 517515 459205 517516
rect 460795 517580 460861 517581
rect 460795 517516 460796 517580
rect 460860 517516 460861 517580
rect 460795 517515 460861 517516
rect 462083 517580 462149 517581
rect 462083 517516 462084 517580
rect 462148 517516 462149 517580
rect 462083 517515 462149 517516
rect 463555 517580 463621 517581
rect 463555 517516 463556 517580
rect 463620 517516 463621 517580
rect 463555 517515 463621 517516
rect 464843 517580 464909 517581
rect 464843 517516 464844 517580
rect 464908 517516 464909 517580
rect 464843 517515 464909 517516
rect 466131 517580 466197 517581
rect 466131 517516 466132 517580
rect 466196 517516 466197 517580
rect 466131 517515 466197 517516
rect 467235 517580 467301 517581
rect 467235 517516 467236 517580
rect 467300 517516 467301 517580
rect 467235 517515 467301 517516
rect 469075 517580 469141 517581
rect 469075 517516 469076 517580
rect 469140 517516 469141 517580
rect 469075 517515 469141 517516
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 483000 415404 487898
rect 418404 492054 419004 517000
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 483000 419004 491498
rect 422004 495654 422604 517000
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 483000 422604 495098
rect 425604 499254 426204 517000
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 483000 426204 498698
rect 432804 506454 433404 517000
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 483000 433404 505898
rect 436404 510054 437004 517000
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 483000 437004 509498
rect 440004 513654 440604 517000
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 483000 440604 513098
rect 443604 483000 444204 517000
rect 450804 488454 451404 517000
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 483000 451404 487898
rect 454404 492054 455004 517000
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 483000 455004 491498
rect 458004 495654 458604 517000
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 483000 458604 495098
rect 461604 499254 462204 517000
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 483000 462204 498698
rect 468804 506454 469404 517000
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 483000 469404 505898
rect 472404 510054 473004 517000
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 483000 473004 509498
rect 476004 513654 476604 517000
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 483000 476604 513098
rect 479604 483000 480204 517000
rect 486804 488454 487404 517000
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 483000 487404 487898
rect 490404 492054 491004 517000
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 483000 491004 491498
rect 494004 495654 494604 517000
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 483000 494604 495098
rect 497604 499254 498204 517000
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 483000 498204 498698
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 483000 505404 505898
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 483000 509004 509498
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 483000 512604 513098
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 520595 700772 520661 700773
rect 520595 700708 520596 700772
rect 520660 700708 520661 700772
rect 520595 700707 520661 700708
rect 518939 700636 519005 700637
rect 518939 700572 518940 700636
rect 519004 700572 519005 700636
rect 518939 700571 519005 700572
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 483000 516204 516698
rect 357387 480044 357453 480045
rect 357387 479980 357388 480044
rect 357452 479980 357453 480044
rect 357387 479979 357453 479980
rect 376707 480044 376773 480045
rect 376707 479980 376708 480044
rect 376772 479980 376773 480044
rect 376707 479979 376773 479980
rect 318747 479636 318813 479637
rect 318747 479572 318748 479636
rect 318812 479572 318813 479636
rect 318747 479571 318813 479572
rect 318750 479365 318810 479571
rect 357390 479365 357450 479979
rect 376710 479637 376770 479979
rect 434667 479772 434733 479773
rect 434667 479708 434668 479772
rect 434732 479708 434733 479772
rect 434667 479707 434733 479708
rect 376707 479636 376773 479637
rect 376707 479572 376708 479636
rect 376772 479572 376773 479636
rect 376707 479571 376773 479572
rect 434670 479501 434730 479707
rect 511947 479636 512013 479637
rect 511947 479572 511948 479636
rect 512012 479572 512013 479636
rect 511947 479571 512013 479572
rect 434667 479500 434733 479501
rect 434667 479436 434668 479500
rect 434732 479436 434733 479500
rect 434667 479435 434733 479436
rect 511950 479365 512010 479571
rect 318747 479364 318813 479365
rect 318747 479300 318748 479364
rect 318812 479300 318813 479364
rect 318747 479299 318813 479300
rect 357387 479364 357453 479365
rect 357387 479300 357388 479364
rect 357452 479300 357453 479364
rect 357387 479299 357453 479300
rect 511947 479364 512013 479365
rect 511947 479300 511948 479364
rect 512012 479300 512013 479364
rect 511947 479299 512013 479300
rect 284208 470454 284528 470476
rect 284208 470218 284250 470454
rect 284486 470218 284528 470454
rect 284208 470134 284528 470218
rect 284208 469898 284250 470134
rect 284486 469898 284528 470134
rect 284208 469876 284528 469898
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 299568 452454 299888 452476
rect 299568 452218 299610 452454
rect 299846 452218 299888 452454
rect 299568 452134 299888 452218
rect 299568 451898 299610 452134
rect 299846 451898 299888 452134
rect 299568 451876 299888 451898
rect 284208 434454 284528 434476
rect 284208 434218 284250 434454
rect 284486 434218 284528 434454
rect 284208 434134 284528 434218
rect 284208 433898 284250 434134
rect 284486 433898 284528 434134
rect 284208 433876 284528 433898
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 299568 416454 299888 416476
rect 299568 416218 299610 416454
rect 299846 416218 299888 416454
rect 299568 416134 299888 416218
rect 299568 415898 299610 416134
rect 299846 415898 299888 416134
rect 299568 415876 299888 415898
rect 518942 409050 519002 700571
rect 519491 695604 519557 695605
rect 519491 695540 519492 695604
rect 519556 695540 519557 695604
rect 519491 695539 519557 695540
rect 519494 695333 519554 695539
rect 519491 695332 519557 695333
rect 519491 695268 519492 695332
rect 519556 695268 519557 695332
rect 519491 695267 519557 695268
rect 519675 686084 519741 686085
rect 519675 686020 519676 686084
rect 519740 686020 519741 686084
rect 519675 686019 519741 686020
rect 519678 685810 519738 686019
rect 519678 685750 519922 685810
rect 519862 684453 519922 685750
rect 519859 684452 519925 684453
rect 519859 684388 519860 684452
rect 519924 684388 519925 684452
rect 519859 684387 519925 684388
rect 519307 681868 519373 681869
rect 519307 681804 519308 681868
rect 519372 681804 519373 681868
rect 519307 681803 519373 681804
rect 519123 644604 519189 644605
rect 519123 644540 519124 644604
rect 519188 644540 519189 644604
rect 519123 644539 519189 644540
rect 519126 644469 519186 644539
rect 519123 644468 519189 644469
rect 519123 644404 519124 644468
rect 519188 644404 519189 644468
rect 519123 644403 519189 644404
rect 519123 634948 519189 634949
rect 519123 634884 519124 634948
rect 519188 634884 519189 634948
rect 519123 634883 519189 634884
rect 519126 625157 519186 634883
rect 519123 625156 519189 625157
rect 519123 625092 519124 625156
rect 519188 625092 519189 625156
rect 519123 625091 519189 625092
rect 519123 615636 519189 615637
rect 519123 615572 519124 615636
rect 519188 615572 519189 615636
rect 519123 615571 519189 615572
rect 519126 605845 519186 615571
rect 519123 605844 519189 605845
rect 519123 605780 519124 605844
rect 519188 605780 519189 605844
rect 519123 605779 519189 605780
rect 519123 596324 519189 596325
rect 519123 596260 519124 596324
rect 519188 596260 519189 596324
rect 519123 596259 519189 596260
rect 519126 586397 519186 596259
rect 519123 586396 519189 586397
rect 519123 586332 519124 586396
rect 519188 586332 519189 586396
rect 519123 586331 519189 586332
rect 519123 576876 519189 576877
rect 519123 576812 519124 576876
rect 519188 576812 519189 576876
rect 519123 576811 519189 576812
rect 519126 567085 519186 576811
rect 519123 567084 519189 567085
rect 519123 567020 519124 567084
rect 519188 567020 519189 567084
rect 519123 567019 519189 567020
rect 519123 557564 519189 557565
rect 519123 557500 519124 557564
rect 519188 557500 519189 557564
rect 519123 557499 519189 557500
rect 519126 547773 519186 557499
rect 519123 547772 519189 547773
rect 519123 547708 519124 547772
rect 519188 547708 519189 547772
rect 519123 547707 519189 547708
rect 519123 538252 519189 538253
rect 519123 538188 519124 538252
rect 519188 538188 519189 538252
rect 519123 538187 519189 538188
rect 519126 528461 519186 538187
rect 519123 528460 519189 528461
rect 519123 528396 519124 528460
rect 519188 528396 519189 528460
rect 519123 528395 519189 528396
rect 519123 518940 519189 518941
rect 519123 518876 519124 518940
rect 519188 518876 519189 518940
rect 519123 518875 519189 518876
rect 519126 509149 519186 518875
rect 519123 509148 519189 509149
rect 519123 509084 519124 509148
rect 519188 509084 519189 509148
rect 519123 509083 519189 509084
rect 519123 499628 519189 499629
rect 519123 499564 519124 499628
rect 519188 499564 519189 499628
rect 519123 499563 519189 499564
rect 519126 489837 519186 499563
rect 519123 489836 519189 489837
rect 519123 489772 519124 489836
rect 519188 489772 519189 489836
rect 519123 489771 519189 489772
rect 519123 479636 519189 479637
rect 519123 479572 519124 479636
rect 519188 479572 519189 479636
rect 519123 479571 519189 479572
rect 519126 466306 519186 479571
rect 519310 475829 519370 681803
rect 520043 666636 520109 666637
rect 520043 666572 520044 666636
rect 520108 666572 520109 666636
rect 520043 666571 520109 666572
rect 520046 659701 520106 666571
rect 519491 659700 519557 659701
rect 519491 659636 519492 659700
rect 519556 659636 519557 659700
rect 519491 659635 519557 659636
rect 520043 659700 520109 659701
rect 520043 659636 520044 659700
rect 520108 659636 520109 659700
rect 520043 659635 520109 659636
rect 519494 653170 519554 659635
rect 519494 653110 519922 653170
rect 519491 652900 519557 652901
rect 519491 652836 519492 652900
rect 519556 652836 519557 652900
rect 519491 652835 519557 652836
rect 519494 475829 519554 652835
rect 519862 644605 519922 653110
rect 519859 644604 519925 644605
rect 519859 644540 519860 644604
rect 519924 644540 519925 644604
rect 519859 644539 519925 644540
rect 519675 644468 519741 644469
rect 519675 644404 519676 644468
rect 519740 644404 519741 644468
rect 519675 644403 519741 644404
rect 519678 634949 519738 644403
rect 519675 634948 519741 634949
rect 519675 634884 519676 634948
rect 519740 634884 519741 634948
rect 519675 634883 519741 634884
rect 519859 625156 519925 625157
rect 519859 625092 519860 625156
rect 519924 625092 519925 625156
rect 519859 625091 519925 625092
rect 519675 623796 519741 623797
rect 519675 623732 519676 623796
rect 519740 623732 519741 623796
rect 519675 623731 519741 623732
rect 519678 475829 519738 623731
rect 519862 615637 519922 625091
rect 519859 615636 519925 615637
rect 519859 615572 519860 615636
rect 519924 615572 519925 615636
rect 519859 615571 519925 615572
rect 519859 605844 519925 605845
rect 519859 605780 519860 605844
rect 519924 605780 519925 605844
rect 519859 605779 519925 605780
rect 519862 596325 519922 605779
rect 519859 596324 519925 596325
rect 519859 596260 519860 596324
rect 519924 596260 519925 596324
rect 519859 596259 519925 596260
rect 519859 586396 519925 586397
rect 519859 586332 519860 586396
rect 519924 586332 519925 586396
rect 519859 586331 519925 586332
rect 519862 576877 519922 586331
rect 519859 576876 519925 576877
rect 519859 576812 519860 576876
rect 519924 576812 519925 576876
rect 519859 576811 519925 576812
rect 519859 567084 519925 567085
rect 519859 567020 519860 567084
rect 519924 567020 519925 567084
rect 519859 567019 519925 567020
rect 519862 557565 519922 567019
rect 519859 557564 519925 557565
rect 519859 557500 519860 557564
rect 519924 557500 519925 557564
rect 519859 557499 519925 557500
rect 519859 547772 519925 547773
rect 519859 547708 519860 547772
rect 519924 547708 519925 547772
rect 519859 547707 519925 547708
rect 519862 538253 519922 547707
rect 519859 538252 519925 538253
rect 519859 538188 519860 538252
rect 519924 538188 519925 538252
rect 519859 538187 519925 538188
rect 519859 528460 519925 528461
rect 519859 528396 519860 528460
rect 519924 528396 519925 528460
rect 519859 528395 519925 528396
rect 519862 518941 519922 528395
rect 519859 518940 519925 518941
rect 519859 518876 519860 518940
rect 519924 518876 519925 518940
rect 519859 518875 519925 518876
rect 519859 509148 519925 509149
rect 519859 509084 519860 509148
rect 519924 509084 519925 509148
rect 519859 509083 519925 509084
rect 519862 499629 519922 509083
rect 519859 499628 519925 499629
rect 519859 499564 519860 499628
rect 519924 499564 519925 499628
rect 519859 499563 519925 499564
rect 519859 489836 519925 489837
rect 519859 489772 519860 489836
rect 519924 489772 519925 489836
rect 519859 489771 519925 489772
rect 519862 479637 519922 489771
rect 519859 479636 519925 479637
rect 519859 479572 519860 479636
rect 519924 479572 519925 479636
rect 519859 479571 519925 479572
rect 519859 479364 519925 479365
rect 519859 479300 519860 479364
rect 519924 479300 519925 479364
rect 519859 479299 519925 479300
rect 519862 475829 519922 479299
rect 520411 476236 520477 476237
rect 520411 476172 520412 476236
rect 520476 476172 520477 476236
rect 520411 476171 520477 476172
rect 520414 476101 520474 476171
rect 520411 476100 520477 476101
rect 520411 476036 520412 476100
rect 520476 476036 520477 476100
rect 520411 476035 520477 476036
rect 519307 475828 519373 475829
rect 519307 475764 519308 475828
rect 519372 475764 519373 475828
rect 519307 475763 519373 475764
rect 519491 475828 519557 475829
rect 519491 475764 519492 475828
rect 519556 475764 519557 475828
rect 519491 475763 519557 475764
rect 519675 475828 519741 475829
rect 519675 475764 519676 475828
rect 519740 475764 519741 475828
rect 519675 475763 519741 475764
rect 519859 475828 519925 475829
rect 519859 475764 519860 475828
rect 519924 475764 519925 475828
rect 519859 475763 519925 475764
rect 519307 475556 519373 475557
rect 519307 475492 519308 475556
rect 519372 475492 519373 475556
rect 519307 475491 519373 475492
rect 519491 475556 519557 475557
rect 519491 475492 519492 475556
rect 519556 475492 519557 475556
rect 519491 475491 519557 475492
rect 519675 475556 519741 475557
rect 519675 475492 519676 475556
rect 519740 475492 519741 475556
rect 519675 475491 519741 475492
rect 519859 475556 519925 475557
rect 519859 475492 519860 475556
rect 519924 475492 519925 475556
rect 519859 475491 519925 475492
rect 519310 468757 519370 475491
rect 519307 468756 519373 468757
rect 519307 468692 519308 468756
rect 519372 468692 519373 468756
rect 519307 468691 519373 468692
rect 519494 468621 519554 475491
rect 519491 468620 519557 468621
rect 519491 468556 519492 468620
rect 519556 468556 519557 468620
rect 519491 468555 519557 468556
rect 519678 466445 519738 475491
rect 519862 466581 519922 475491
rect 520227 472700 520293 472701
rect 520227 472636 520228 472700
rect 520292 472636 520293 472700
rect 520227 472635 520293 472636
rect 519859 466580 519925 466581
rect 519859 466516 519860 466580
rect 519924 466516 519925 466580
rect 519859 466515 519925 466516
rect 519675 466444 519741 466445
rect 519675 466380 519676 466444
rect 519740 466380 519741 466444
rect 519675 466379 519741 466380
rect 519126 466246 520106 466306
rect 519675 466036 519741 466037
rect 519675 465972 519676 466036
rect 519740 465972 519741 466036
rect 519675 465971 519741 465972
rect 519491 465628 519557 465629
rect 519491 465564 519492 465628
rect 519556 465564 519557 465628
rect 519491 465563 519557 465564
rect 519307 465492 519373 465493
rect 519307 465428 519308 465492
rect 519372 465428 519373 465492
rect 519307 465427 519373 465428
rect 519310 453250 519370 465427
rect 519126 453190 519370 453250
rect 519126 446994 519186 453190
rect 519494 452709 519554 465563
rect 519678 452709 519738 465971
rect 519859 465900 519925 465901
rect 519859 465836 519860 465900
rect 519924 465836 519925 465900
rect 519859 465835 519925 465836
rect 519862 452709 519922 465835
rect 519491 452708 519557 452709
rect 519491 452644 519492 452708
rect 519556 452644 519557 452708
rect 519491 452643 519557 452644
rect 519675 452708 519741 452709
rect 519675 452644 519676 452708
rect 519740 452644 519741 452708
rect 519675 452643 519741 452644
rect 519859 452708 519925 452709
rect 519859 452644 519860 452708
rect 519924 452644 519925 452708
rect 519859 452643 519925 452644
rect 519491 452436 519557 452437
rect 519491 452372 519492 452436
rect 519556 452372 519557 452436
rect 519491 452371 519557 452372
rect 519675 452436 519741 452437
rect 519675 452372 519676 452436
rect 519740 452372 519741 452436
rect 519675 452371 519741 452372
rect 519859 452436 519925 452437
rect 519859 452372 519860 452436
rect 519924 452372 519925 452436
rect 519859 452371 519925 452372
rect 519126 446934 519370 446994
rect 519310 428770 519370 446934
rect 519126 428710 519370 428770
rect 519126 427410 519186 428710
rect 519126 427350 519370 427410
rect 519310 415581 519370 427350
rect 519307 415580 519373 415581
rect 519307 415516 519308 415580
rect 519372 415516 519373 415580
rect 519307 415515 519373 415516
rect 519494 415309 519554 452371
rect 519678 429725 519738 452371
rect 519675 429724 519741 429725
rect 519675 429660 519676 429724
rect 519740 429660 519741 429724
rect 519675 429659 519741 429660
rect 519675 427956 519741 427957
rect 519675 427892 519676 427956
rect 519740 427892 519741 427956
rect 519675 427891 519741 427892
rect 519491 415308 519557 415309
rect 519491 415244 519492 415308
rect 519556 415244 519557 415308
rect 519491 415243 519557 415244
rect 519307 415036 519373 415037
rect 519307 414972 519308 415036
rect 519372 414972 519373 415036
rect 519307 414971 519373 414972
rect 519310 409189 519370 414971
rect 519307 409188 519373 409189
rect 519307 409124 519308 409188
rect 519372 409124 519373 409188
rect 519307 409123 519373 409124
rect 518942 408990 519554 409050
rect 519307 407012 519373 407013
rect 519307 407010 519308 407012
rect 518758 406950 519308 407010
rect 518758 405650 518818 406950
rect 519307 406948 519308 406950
rect 519372 406948 519373 407012
rect 519307 406947 519373 406948
rect 519494 406333 519554 408990
rect 519678 408781 519738 427891
rect 519862 415309 519922 452371
rect 520046 437749 520106 466246
rect 520043 437748 520109 437749
rect 520043 437684 520044 437748
rect 520108 437684 520109 437748
rect 520043 437683 520109 437684
rect 520043 437612 520109 437613
rect 520043 437548 520044 437612
rect 520108 437548 520109 437612
rect 520043 437547 520109 437548
rect 520046 435301 520106 437547
rect 520043 435300 520109 435301
rect 520043 435236 520044 435300
rect 520108 435236 520109 435300
rect 520043 435235 520109 435236
rect 520043 435164 520109 435165
rect 520043 435100 520044 435164
rect 520108 435100 520109 435164
rect 520043 435099 520109 435100
rect 520046 429861 520106 435099
rect 520043 429860 520109 429861
rect 520043 429796 520044 429860
rect 520108 429796 520109 429860
rect 520043 429795 520109 429796
rect 520043 429724 520109 429725
rect 520043 429660 520044 429724
rect 520108 429660 520109 429724
rect 520043 429659 520109 429660
rect 520046 428093 520106 429659
rect 520043 428092 520109 428093
rect 520043 428028 520044 428092
rect 520108 428028 520109 428092
rect 520043 428027 520109 428028
rect 520043 425100 520109 425101
rect 520043 425036 520044 425100
rect 520108 425036 520109 425100
rect 520043 425035 520109 425036
rect 519859 415308 519925 415309
rect 519859 415244 519860 415308
rect 519924 415244 519925 415308
rect 519859 415243 519925 415244
rect 519859 415036 519925 415037
rect 519859 414972 519860 415036
rect 519924 414972 519925 415036
rect 519859 414971 519925 414972
rect 519675 408780 519741 408781
rect 519675 408716 519676 408780
rect 519740 408716 519741 408780
rect 519675 408715 519741 408716
rect 519675 408372 519741 408373
rect 519675 408308 519676 408372
rect 519740 408308 519741 408372
rect 519675 408307 519741 408308
rect 519491 406332 519557 406333
rect 519491 406268 519492 406332
rect 519556 406268 519557 406332
rect 519491 406267 519557 406268
rect 519307 406196 519373 406197
rect 519307 406194 519308 406196
rect 518574 405590 518818 405650
rect 518942 406134 519308 406194
rect 284208 398454 284528 398476
rect 284208 398218 284250 398454
rect 284486 398218 284528 398454
rect 284208 398134 284528 398218
rect 284208 397898 284250 398134
rect 284486 397898 284528 398134
rect 284208 397876 284528 397898
rect 518574 393410 518634 405590
rect 518942 396130 519002 406134
rect 519307 406132 519308 406134
rect 519372 406132 519373 406196
rect 519307 406131 519373 406132
rect 519491 406196 519557 406197
rect 519491 406132 519492 406196
rect 519556 406132 519557 406196
rect 519491 406131 519557 406132
rect 519307 406060 519373 406061
rect 519307 405996 519308 406060
rect 519372 405996 519373 406060
rect 519307 405995 519373 405996
rect 519310 396405 519370 405995
rect 519307 396404 519373 396405
rect 519307 396340 519308 396404
rect 519372 396340 519373 396404
rect 519307 396339 519373 396340
rect 518942 396070 519370 396130
rect 519310 395589 519370 396070
rect 519307 395588 519373 395589
rect 519307 395524 519308 395588
rect 519372 395524 519373 395588
rect 519307 395523 519373 395524
rect 519494 395317 519554 406131
rect 519678 399533 519738 408307
rect 519675 399532 519741 399533
rect 519675 399468 519676 399532
rect 519740 399468 519741 399532
rect 519675 399467 519741 399468
rect 519491 395316 519557 395317
rect 519491 395252 519492 395316
rect 519556 395252 519557 395316
rect 519491 395251 519557 395252
rect 519307 393412 519373 393413
rect 519307 393410 519308 393412
rect 518574 393350 519308 393410
rect 519307 393348 519308 393350
rect 519372 393348 519373 393412
rect 519307 393347 519373 393348
rect 519675 393412 519741 393413
rect 519675 393348 519676 393412
rect 519740 393348 519741 393412
rect 519675 393347 519741 393348
rect 519307 390692 519373 390693
rect 519307 390628 519308 390692
rect 519372 390628 519373 390692
rect 519307 390627 519373 390628
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 519310 382261 519370 390627
rect 519678 388925 519738 393347
rect 519675 388924 519741 388925
rect 519675 388860 519676 388924
rect 519740 388860 519741 388924
rect 519675 388859 519741 388860
rect 519862 386069 519922 414971
rect 520046 407013 520106 425035
rect 520043 407012 520109 407013
rect 520043 406948 520044 407012
rect 520108 406948 520109 407012
rect 520043 406947 520109 406948
rect 519859 386068 519925 386069
rect 519859 386004 519860 386068
rect 519924 386004 519925 386068
rect 519859 386003 519925 386004
rect 519307 382260 519373 382261
rect 519307 382196 519308 382260
rect 519372 382196 519373 382260
rect 519307 382195 519373 382196
rect 299568 380454 299888 380476
rect 299568 380218 299610 380454
rect 299846 380218 299888 380454
rect 299568 380134 299888 380218
rect 299568 379898 299610 380134
rect 299846 379898 299888 380134
rect 299568 379876 299888 379898
rect 284208 362454 284528 362476
rect 284208 362218 284250 362454
rect 284486 362218 284528 362454
rect 284208 362134 284528 362218
rect 284208 361898 284250 362134
rect 284486 361898 284528 362134
rect 284208 361876 284528 361898
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 299568 344454 299888 344476
rect 299568 344218 299610 344454
rect 299846 344218 299888 344454
rect 299568 344134 299888 344218
rect 299568 343898 299610 344134
rect 299846 343898 299888 344134
rect 299568 343876 299888 343898
rect 284208 326454 284528 326476
rect 284208 326218 284250 326454
rect 284486 326218 284528 326454
rect 284208 326134 284528 326218
rect 284208 325898 284250 326134
rect 284486 325898 284528 326134
rect 284208 325876 284528 325898
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 299568 308454 299888 308476
rect 299568 308218 299610 308454
rect 299846 308218 299888 308454
rect 299568 308134 299888 308218
rect 299568 307898 299610 308134
rect 299846 307898 299888 308134
rect 299568 307876 299888 307898
rect 284208 290454 284528 290476
rect 284208 290218 284250 290454
rect 284486 290218 284528 290454
rect 284208 290134 284528 290218
rect 284208 289898 284250 290134
rect 284486 289898 284528 290134
rect 284208 289876 284528 289898
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 299568 272454 299888 272476
rect 299568 272218 299610 272454
rect 299846 272218 299888 272454
rect 299568 272134 299888 272218
rect 299568 271898 299610 272134
rect 299846 271898 299888 272134
rect 299568 271876 299888 271898
rect 284208 254454 284528 254476
rect 284208 254218 284250 254454
rect 284486 254218 284528 254454
rect 284208 254134 284528 254218
rect 284208 253898 284250 254134
rect 284486 253898 284528 254134
rect 284208 253876 284528 253898
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 207654 278604 237000
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 211254 282204 237000
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 218454 289404 237000
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 222054 293004 237000
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 225654 296604 237000
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 299604 229254 300204 237000
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 204247 300204 228698
rect 306804 236454 307404 237000
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 204247 307404 235898
rect 310404 204247 311004 237000
rect 314004 207654 314604 237000
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 204247 314604 207098
rect 317604 211254 318204 237000
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 204247 318204 210698
rect 324804 218454 325404 237000
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 204247 325404 217898
rect 328404 222054 329004 237000
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 204247 329004 221498
rect 332004 225654 332604 237000
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 329419 212532 329485 212533
rect 329419 212468 329420 212532
rect 329484 212468 329485 212532
rect 329419 212467 329485 212468
rect 328131 203284 328197 203285
rect 328131 203220 328132 203284
rect 328196 203220 328197 203284
rect 328131 203219 328197 203220
rect 328134 200970 328194 203219
rect 328315 203148 328381 203149
rect 328315 203084 328316 203148
rect 328380 203084 328381 203148
rect 328315 203083 328381 203084
rect 328318 201650 328378 203083
rect 328318 201590 328446 201650
rect 328134 200910 328292 200970
rect 328386 200940 328446 201590
rect 329422 200910 329482 212467
rect 332004 204247 332604 225098
rect 335604 229254 336204 237000
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 204247 336204 228698
rect 342804 236454 343404 237000
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 336411 220828 336477 220829
rect 336411 220764 336412 220828
rect 336476 220764 336477 220828
rect 336411 220763 336477 220764
rect 330891 203692 330957 203693
rect 330891 203628 330892 203692
rect 330956 203628 330957 203692
rect 330891 203627 330957 203628
rect 329603 203420 329669 203421
rect 329603 203356 329604 203420
rect 329668 203356 329669 203420
rect 329603 203355 329669 203356
rect 330707 203420 330773 203421
rect 330707 203356 330708 203420
rect 330772 203356 330773 203420
rect 330707 203355 330773 203356
rect 329606 200970 329666 203355
rect 330710 201650 330770 203355
rect 329584 200910 329666 200970
rect 330598 201590 330770 201650
rect 330598 200940 330658 201590
rect 330894 200970 330954 203627
rect 334203 203420 334269 203421
rect 334203 203356 334204 203420
rect 334268 203356 334269 203420
rect 334203 203355 334269 203356
rect 331627 203284 331693 203285
rect 331627 203220 331628 203284
rect 331692 203220 331693 203284
rect 331627 203219 331693 203220
rect 332915 203284 332981 203285
rect 332915 203220 332916 203284
rect 332980 203220 332981 203284
rect 332915 203219 332981 203220
rect 330752 200910 330954 200970
rect 331630 200970 331690 203219
rect 332363 203148 332429 203149
rect 332363 203084 332364 203148
rect 332428 203084 332429 203148
rect 332363 203083 332429 203084
rect 332366 200970 332426 203083
rect 331630 200910 331796 200970
rect 331920 200910 332426 200970
rect 332918 200910 332978 203219
rect 333651 203148 333717 203149
rect 333651 203084 333652 203148
rect 333716 203084 333717 203148
rect 333651 203083 333717 203084
rect 333654 200970 333714 203083
rect 334206 201650 334266 203355
rect 335123 203284 335189 203285
rect 335123 203220 335124 203284
rect 335188 203220 335189 203284
rect 335123 203219 335189 203220
rect 334755 203012 334821 203013
rect 334755 202948 334756 203012
rect 334820 202948 334821 203012
rect 334755 202947 334821 202948
rect 333088 200910 333714 200970
rect 334102 201590 334266 201650
rect 334102 200940 334162 201590
rect 334758 200970 334818 202947
rect 334256 200910 334818 200970
rect 335126 200970 335186 203219
rect 336043 203012 336109 203013
rect 336043 202948 336044 203012
rect 336108 202948 336109 203012
rect 336043 202947 336109 202948
rect 336046 200970 336106 202947
rect 335126 200910 335300 200970
rect 335424 200910 336106 200970
rect 336414 200910 336474 220763
rect 342804 204247 343404 235898
rect 346404 204247 347004 237000
rect 350004 207654 350604 237000
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 204247 350604 207098
rect 353604 211254 354204 237000
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 204247 354204 210698
rect 360804 218454 361404 237000
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 204247 361404 217898
rect 364404 222054 365004 237000
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 204247 365004 221498
rect 368004 225654 368604 237000
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 204247 368604 225098
rect 371604 229254 372204 237000
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 204247 372204 228698
rect 378804 236454 379404 237000
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 204247 379404 235898
rect 382404 204054 383004 237000
rect 357387 203964 357453 203965
rect 357387 203900 357388 203964
rect 357452 203900 357453 203964
rect 357387 203899 357453 203900
rect 360515 203964 360581 203965
rect 360515 203900 360516 203964
rect 360580 203900 360581 203964
rect 360515 203899 360581 203900
rect 341011 203692 341077 203693
rect 341011 203628 341012 203692
rect 341076 203628 341077 203692
rect 341011 203627 341077 203628
rect 342851 203692 342917 203693
rect 342851 203628 342852 203692
rect 342916 203628 342917 203692
rect 342851 203627 342917 203628
rect 347819 203692 347885 203693
rect 347819 203628 347820 203692
rect 347884 203628 347885 203692
rect 347819 203627 347885 203628
rect 349107 203692 349173 203693
rect 349107 203628 349108 203692
rect 349172 203628 349173 203692
rect 349107 203627 349173 203628
rect 352787 203692 352853 203693
rect 352787 203628 352788 203692
rect 352852 203628 352853 203692
rect 352787 203627 352853 203628
rect 340091 203556 340157 203557
rect 340091 203492 340092 203556
rect 340156 203492 340157 203556
rect 340091 203491 340157 203492
rect 336963 203420 337029 203421
rect 336963 203356 336964 203420
rect 337028 203356 337029 203420
rect 336963 203355 337029 203356
rect 336595 203148 336661 203149
rect 336595 203084 336596 203148
rect 336660 203084 336661 203148
rect 336595 203083 336661 203084
rect 336598 200970 336658 203083
rect 336592 200910 336658 200970
rect 336966 200970 337026 203355
rect 338435 203284 338501 203285
rect 338435 203220 338436 203284
rect 338500 203220 338501 203284
rect 338435 203219 338501 203220
rect 339723 203284 339789 203285
rect 339723 203220 339724 203284
rect 339788 203220 339789 203284
rect 339723 203219 339789 203220
rect 337883 203012 337949 203013
rect 337883 202948 337884 203012
rect 337948 202948 337949 203012
rect 337883 202947 337949 202948
rect 337886 200970 337946 202947
rect 336966 200910 337636 200970
rect 337760 200910 337946 200970
rect 338438 200970 338498 203219
rect 339171 203012 339237 203013
rect 339171 202948 339172 203012
rect 339236 202948 339237 203012
rect 339171 202947 339237 202948
rect 338438 200910 338804 200970
rect 339174 200817 339234 202947
rect 339726 200970 339786 203219
rect 339726 200910 339972 200970
rect 340094 200910 340154 203491
rect 341014 201650 341074 203627
rect 342299 203556 342365 203557
rect 342299 203492 342300 203556
rect 342364 203492 342365 203556
rect 342299 203491 342365 203492
rect 341379 203012 341445 203013
rect 341379 202948 341380 203012
rect 341444 202948 341445 203012
rect 341379 202947 341445 202948
rect 341014 201590 341170 201650
rect 341110 200940 341170 201590
rect 341382 200970 341442 202947
rect 342302 201789 342362 203491
rect 342483 203420 342549 203421
rect 342483 203356 342484 203420
rect 342548 203356 342549 203420
rect 342483 203355 342549 203356
rect 342299 201788 342365 201789
rect 342299 201724 342300 201788
rect 342364 201724 342365 201788
rect 342299 201723 342365 201724
rect 342486 201650 342546 203355
rect 342402 201590 342546 201650
rect 342275 201516 342341 201517
rect 342275 201452 342276 201516
rect 342340 201452 342341 201516
rect 342275 201451 342341 201452
rect 341264 200910 341442 200970
rect 342278 200940 342338 201451
rect 342402 200940 342462 201590
rect 342854 200970 342914 203627
rect 343587 203556 343653 203557
rect 343587 203492 343588 203556
rect 343652 203492 343653 203556
rect 343587 203491 343653 203492
rect 342854 200910 343476 200970
rect 343590 200910 343650 203491
rect 346531 203284 346597 203285
rect 346531 203220 346532 203284
rect 346596 203220 346597 203284
rect 346531 203219 346597 203220
rect 343955 203148 344021 203149
rect 343955 203084 343956 203148
rect 344020 203084 344021 203148
rect 343955 203083 344021 203084
rect 345243 203148 345309 203149
rect 345243 203084 345244 203148
rect 345308 203084 345309 203148
rect 345243 203083 345309 203084
rect 343958 200970 344018 203083
rect 344875 203012 344941 203013
rect 344875 202948 344876 203012
rect 344940 202948 344941 203012
rect 344875 202947 344941 202948
rect 344878 200970 344938 202947
rect 343958 200910 344644 200970
rect 344768 200910 344938 200970
rect 345246 200970 345306 203083
rect 345979 203012 346045 203013
rect 345979 202948 345980 203012
rect 346044 202948 346045 203012
rect 345979 202947 346045 202948
rect 345982 201650 346042 202947
rect 345906 201590 346042 201650
rect 345246 200910 345812 200970
rect 345906 200940 345966 201590
rect 346534 200970 346594 203219
rect 347083 203012 347149 203013
rect 347083 202948 347084 203012
rect 347148 202948 347149 203012
rect 347083 202947 347149 202948
rect 346534 200910 346980 200970
rect 347086 200910 347146 202947
rect 347822 200970 347882 203627
rect 348371 203012 348437 203013
rect 348371 202948 348372 203012
rect 348436 202948 348437 203012
rect 348371 202947 348437 202948
rect 348374 200970 348434 202947
rect 347822 200910 348148 200970
rect 348272 200910 348434 200970
rect 349110 200970 349170 203627
rect 349843 203284 349909 203285
rect 349843 203220 349844 203284
rect 349908 203220 349909 203284
rect 349843 203219 349909 203220
rect 349475 203012 349541 203013
rect 349475 202948 349476 203012
rect 349540 202948 349541 203012
rect 349475 202947 349541 202948
rect 349478 201650 349538 202947
rect 349410 201590 349538 201650
rect 349110 200910 349316 200970
rect 349410 200940 349470 201590
rect 349846 200970 349906 203219
rect 351131 203148 351197 203149
rect 351131 203084 351132 203148
rect 351196 203084 351197 203148
rect 351131 203083 351197 203084
rect 350947 203012 351013 203013
rect 350947 202948 350948 203012
rect 351012 202948 351013 203012
rect 350947 202947 351013 202948
rect 350950 200970 351010 202947
rect 349846 200910 350484 200970
rect 350608 200910 351010 200970
rect 351134 200970 351194 203083
rect 351683 203012 351749 203013
rect 351683 202948 351684 203012
rect 351748 202948 351749 203012
rect 351683 202947 351749 202948
rect 351686 201650 351746 202947
rect 351686 201590 351806 201650
rect 351134 200910 351652 200970
rect 351746 200940 351806 201590
rect 352790 200940 352850 203627
rect 354811 203556 354877 203557
rect 354811 203492 354812 203556
rect 354876 203492 354877 203556
rect 354811 203491 354877 203492
rect 352971 203012 353037 203013
rect 352971 202948 352972 203012
rect 353036 202948 353037 203012
rect 352971 202947 353037 202948
rect 353339 203012 353405 203013
rect 353339 202948 353340 203012
rect 353404 202948 353405 203012
rect 353339 202947 353405 202948
rect 354443 203012 354509 203013
rect 354443 202948 354444 203012
rect 354508 202948 354509 203012
rect 354443 202947 354509 202948
rect 352974 200970 353034 202947
rect 352944 200910 353034 200970
rect 353342 200970 353402 202947
rect 354446 200970 354506 202947
rect 353342 200910 353988 200970
rect 354112 200910 354506 200970
rect 354814 200970 354874 203491
rect 356099 203284 356165 203285
rect 356099 203220 356100 203284
rect 356164 203220 356165 203284
rect 356099 203219 356165 203220
rect 355547 203012 355613 203013
rect 355547 202948 355548 203012
rect 355612 202948 355613 203012
rect 355547 202947 355613 202948
rect 354814 200910 355156 200970
rect 355550 200817 355610 202947
rect 356102 200970 356162 203219
rect 356467 203012 356533 203013
rect 356467 202948 356468 203012
rect 356532 202948 356533 203012
rect 356467 202947 356533 202948
rect 356470 200970 356530 202947
rect 357390 201650 357450 203899
rect 357755 203148 357821 203149
rect 357755 203084 357756 203148
rect 357820 203084 357821 203148
rect 357755 203083 357821 203084
rect 357390 201590 357522 201650
rect 356102 200910 356324 200970
rect 356448 200910 356530 200970
rect 357462 200940 357522 201590
rect 357758 200970 357818 203083
rect 357939 203012 358005 203013
rect 357939 202948 357940 203012
rect 358004 202948 358005 203012
rect 357939 202947 358005 202948
rect 358675 203012 358741 203013
rect 358675 202948 358676 203012
rect 358740 202948 358741 203012
rect 358675 202947 358741 202948
rect 359227 203012 359293 203013
rect 359227 202948 359228 203012
rect 359292 202948 359293 203012
rect 359227 202947 359293 202948
rect 359963 203012 360029 203013
rect 359963 202948 359964 203012
rect 360028 202948 360029 203012
rect 359963 202947 360029 202948
rect 357616 200910 357818 200970
rect 357942 200970 358002 202947
rect 358678 201650 358738 202947
rect 358678 201590 358814 201650
rect 357942 200910 358660 200970
rect 358754 200940 358814 201590
rect 359230 200970 359290 202947
rect 359966 200970 360026 202947
rect 359230 200910 359828 200970
rect 359952 200910 360026 200970
rect 360518 200970 360578 203899
rect 361619 203828 361685 203829
rect 361619 203764 361620 203828
rect 361684 203764 361685 203828
rect 361619 203763 361685 203764
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 361251 203012 361317 203013
rect 361251 202948 361252 203012
rect 361316 202948 361317 203012
rect 361251 202947 361317 202948
rect 361254 200970 361314 202947
rect 360518 200910 360996 200970
rect 361120 200910 361314 200970
rect 361622 200970 361682 203763
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 362907 203420 362973 203421
rect 362907 203356 362908 203420
rect 362972 203356 362973 203420
rect 362907 203355 362973 203356
rect 364379 203420 364445 203421
rect 364379 203356 364380 203420
rect 364444 203356 364445 203420
rect 364379 203355 364445 203356
rect 367507 203420 367573 203421
rect 367507 203356 367508 203420
rect 367572 203356 367573 203420
rect 367507 203355 367573 203356
rect 362723 203012 362789 203013
rect 362723 202948 362724 203012
rect 362788 202948 362789 203012
rect 362723 202947 362789 202948
rect 361622 200910 362164 200970
rect 362726 200817 362786 202947
rect 362910 200970 362970 203355
rect 363459 203012 363525 203013
rect 363459 202948 363460 203012
rect 363524 202948 363525 203012
rect 363459 202947 363525 202948
rect 363462 200970 363522 202947
rect 364382 201650 364442 203355
rect 366955 203284 367021 203285
rect 366955 203220 366956 203284
rect 367020 203220 367021 203284
rect 366955 203219 367021 203220
rect 366403 203148 366469 203149
rect 366403 203084 366404 203148
rect 366468 203084 366469 203148
rect 366403 203083 366469 203084
rect 364931 203012 364997 203013
rect 364931 202948 364932 203012
rect 364996 202948 364997 203012
rect 364931 202947 364997 202948
rect 364382 201590 364530 201650
rect 362910 200910 363332 200970
rect 363456 200910 363522 200970
rect 364470 200940 364530 201590
rect 364934 200970 364994 202947
rect 366406 200970 366466 203083
rect 364624 200910 364994 200970
rect 365792 200910 366466 200970
rect 366958 200910 367018 203219
rect 367510 200970 367570 203355
rect 368611 203284 368677 203285
rect 368611 203220 368612 203284
rect 368676 203220 368677 203284
rect 368611 203219 368677 203220
rect 371003 203284 371069 203285
rect 371003 203220 371004 203284
rect 371068 203220 371069 203284
rect 371003 203219 371069 203220
rect 368614 200970 368674 203219
rect 371006 200970 371066 203219
rect 373395 203148 373461 203149
rect 373395 203084 373396 203148
rect 373460 203084 373461 203148
rect 373395 203083 373461 203084
rect 367510 200910 368128 200970
rect 368614 200910 369296 200970
rect 370464 200910 371066 200970
rect 373398 200970 373458 203083
rect 373398 200910 373463 200970
rect 338928 200757 339234 200817
rect 355280 200757 355610 200817
rect 362288 200757 362786 200817
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 300482 182454 300802 182476
rect 300482 182218 300524 182454
rect 300760 182218 300802 182454
rect 300482 182134 300802 182218
rect 300482 181898 300524 182134
rect 300760 181898 300802 182134
rect 300482 181876 300802 181898
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 300034 164454 300358 164476
rect 300034 164218 300078 164454
rect 300314 164218 300358 164454
rect 300034 164134 300358 164218
rect 300034 163898 300078 164134
rect 300314 163898 300358 164134
rect 300034 163876 300358 163898
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 300482 146454 300802 146476
rect 300482 146218 300524 146454
rect 300760 146218 300802 146454
rect 300482 146134 300802 146218
rect 300482 145898 300524 146134
rect 300760 145898 300802 146134
rect 300482 145876 300802 145898
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 300034 128454 300358 128476
rect 300034 128218 300078 128454
rect 300314 128218 300358 128454
rect 300034 128134 300358 128218
rect 300034 127898 300078 128134
rect 300314 127898 300358 128134
rect 300034 127876 300358 127898
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 303662 109037 303722 110190
rect 308078 110130 308688 110190
rect 308078 109037 308138 110130
rect 303659 109036 303725 109037
rect 303659 108972 303660 109036
rect 303724 108972 303725 109036
rect 303659 108971 303725 108972
rect 308075 109036 308141 109037
rect 308075 108972 308076 109036
rect 308140 108972 308141 109036
rect 308075 108971 308141 108972
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 85254 300204 107000
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 92454 307404 107000
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 96054 311004 107000
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 99654 314604 107000
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 103254 318204 107000
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 74454 325404 107000
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 78054 329004 107000
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 81654 332604 107000
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 85254 336204 107000
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 92454 343404 107000
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 96054 347004 107000
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 99654 350604 107000
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 103254 354204 107000
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 74454 361404 107000
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 78054 365004 107000
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 81654 368604 107000
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 85254 372204 107000
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 92454 379404 107000
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 207654 386604 237000
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 211254 390204 237000
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 218454 397404 237000
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 222054 401004 237000
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 225654 404604 237000
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 229254 408204 237000
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 236454 415404 237000
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 418404 204247 419004 237000
rect 422004 207654 422604 237000
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 204247 422604 207098
rect 425604 211254 426204 237000
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 204247 426204 210698
rect 432804 218454 433404 237000
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 204247 433404 217898
rect 436404 222054 437004 237000
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 204247 437004 221498
rect 440004 225654 440604 237000
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 204247 440604 225098
rect 443604 229254 444204 237000
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 204247 444204 228698
rect 450804 236454 451404 237000
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 204247 451404 235898
rect 454404 204247 455004 237000
rect 458004 207654 458604 237000
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 204247 458604 207098
rect 461604 211254 462204 237000
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 204247 462204 210698
rect 468804 218454 469404 237000
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 204247 469404 217898
rect 472404 222054 473004 237000
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 204247 473004 221498
rect 476004 225654 476604 237000
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 204247 476604 225098
rect 479604 229254 480204 237000
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 204247 480204 228698
rect 486804 236454 487404 237000
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 204247 487404 235898
rect 490404 204247 491004 237000
rect 494004 207654 494604 237000
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 204247 494604 207098
rect 497604 211254 498204 237000
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 204247 498204 210698
rect 504804 218454 505404 237000
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 448283 204236 448349 204237
rect 448283 204172 448284 204236
rect 448348 204172 448349 204236
rect 448283 204171 448349 204172
rect 449387 204236 449453 204237
rect 449387 204172 449388 204236
rect 449452 204172 449453 204236
rect 449387 204171 449453 204172
rect 451779 204236 451845 204237
rect 451779 204172 451780 204236
rect 451844 204172 451845 204236
rect 451779 204171 451845 204172
rect 453251 204236 453317 204237
rect 453251 204172 453252 204236
rect 453316 204172 453317 204236
rect 453251 204171 453317 204172
rect 454171 204236 454237 204237
rect 454171 204172 454172 204236
rect 454236 204172 454237 204236
rect 454171 204171 454237 204172
rect 456379 204236 456445 204237
rect 456379 204172 456380 204236
rect 456444 204172 456445 204236
rect 456379 204171 456445 204172
rect 468155 204236 468221 204237
rect 468155 204172 468156 204236
rect 468220 204172 468221 204236
rect 468155 204171 468221 204172
rect 470363 204236 470429 204237
rect 470363 204172 470364 204236
rect 470428 204172 470429 204236
rect 470363 204171 470429 204172
rect 484347 204236 484413 204237
rect 484347 204172 484348 204236
rect 484412 204172 484413 204236
rect 484347 204171 484413 204172
rect 448286 201514 448346 204171
rect 448262 201454 448346 201514
rect 448262 200940 448322 201454
rect 448383 201380 448449 201381
rect 448383 201316 448384 201380
rect 448448 201316 448449 201380
rect 448383 201315 448449 201316
rect 448386 200940 448446 201315
rect 449390 200970 449450 204171
rect 449571 204100 449637 204101
rect 449571 204036 449572 204100
rect 449636 204036 449637 204100
rect 449571 204035 449637 204036
rect 450859 204100 450925 204101
rect 450859 204036 450860 204100
rect 450924 204036 450925 204100
rect 450859 204035 450925 204036
rect 449390 200910 449460 200970
rect 449574 200910 449634 204035
rect 450675 203012 450741 203013
rect 450675 202948 450676 203012
rect 450740 202948 450741 203012
rect 450675 202947 450741 202948
rect 450678 201514 450738 202947
rect 450598 201454 450738 201514
rect 450598 200940 450658 201454
rect 450862 200970 450922 204035
rect 451782 201514 451842 204171
rect 452147 204100 452213 204101
rect 452147 204036 452148 204100
rect 452212 204036 452213 204100
rect 452147 204035 452213 204036
rect 450752 200910 450922 200970
rect 451766 201454 451842 201514
rect 451766 200940 451826 201454
rect 452150 200817 452210 204035
rect 452883 203012 452949 203013
rect 452883 202948 452884 203012
rect 452948 202948 452949 203012
rect 452883 202947 452949 202948
rect 452886 200970 452946 202947
rect 453254 200970 453314 204171
rect 454174 201514 454234 204171
rect 454539 204100 454605 204101
rect 454539 204036 454540 204100
rect 454604 204036 454605 204100
rect 454539 204035 454605 204036
rect 452886 200910 452964 200970
rect 453088 200910 453314 200970
rect 454102 201454 454234 201514
rect 454102 200940 454162 201454
rect 454542 200970 454602 204035
rect 456011 203420 456077 203421
rect 456011 203356 456012 203420
rect 456076 203356 456077 203420
rect 456011 203355 456077 203356
rect 455275 203012 455341 203013
rect 455275 202948 455276 203012
rect 455340 202948 455341 203012
rect 455275 202947 455341 202948
rect 455278 201514 455338 202947
rect 454256 200910 454602 200970
rect 455270 201454 455338 201514
rect 455270 200940 455330 201454
rect 456014 200970 456074 203355
rect 455424 200910 456074 200970
rect 456382 200970 456442 204171
rect 456563 204100 456629 204101
rect 456563 204036 456564 204100
rect 456628 204036 456629 204100
rect 456563 204035 456629 204036
rect 464475 204100 464541 204101
rect 464475 204036 464476 204100
rect 464540 204036 464541 204100
rect 464475 204035 464541 204036
rect 465763 204100 465829 204101
rect 465763 204036 465764 204100
rect 465828 204036 465829 204100
rect 465763 204035 465829 204036
rect 456382 200910 456468 200970
rect 456566 200910 456626 204035
rect 457483 203964 457549 203965
rect 457483 203900 457484 203964
rect 457548 203900 457549 203964
rect 457483 203899 457549 203900
rect 460059 203964 460125 203965
rect 460059 203900 460060 203964
rect 460124 203900 460125 203964
rect 460059 203899 460125 203900
rect 457486 200970 457546 203899
rect 458771 203284 458837 203285
rect 458771 203220 458772 203284
rect 458836 203220 458837 203284
rect 458771 203219 458837 203220
rect 457851 203012 457917 203013
rect 457851 202948 457852 203012
rect 457916 202948 457917 203012
rect 457851 202947 457917 202948
rect 457854 200970 457914 202947
rect 457486 200910 457636 200970
rect 457760 200910 457914 200970
rect 458774 200940 458834 203219
rect 458955 203012 459021 203013
rect 458955 202948 458956 203012
rect 459020 202948 459021 203012
rect 458955 202947 459021 202948
rect 458958 200970 459018 202947
rect 460062 201650 460122 203899
rect 462267 203420 462333 203421
rect 462267 203356 462268 203420
rect 462332 203356 462333 203420
rect 462267 203355 462333 203356
rect 460979 203284 461045 203285
rect 460979 203220 460980 203284
rect 461044 203220 461045 203284
rect 460979 203219 461045 203220
rect 460611 203012 460677 203013
rect 460611 202948 460612 203012
rect 460676 202948 460677 203012
rect 460611 202947 460677 202948
rect 458928 200910 459018 200970
rect 459942 201590 460122 201650
rect 459942 200940 460002 201590
rect 460614 200970 460674 202947
rect 460096 200910 460674 200970
rect 460982 200970 461042 203219
rect 461531 203012 461597 203013
rect 461531 202948 461532 203012
rect 461596 202948 461597 203012
rect 461531 202947 461597 202948
rect 460982 200910 461140 200970
rect 461534 200817 461594 202947
rect 462270 200910 462330 203355
rect 463187 203284 463253 203285
rect 463187 203220 463188 203284
rect 463252 203220 463253 203284
rect 463187 203219 463253 203220
rect 462451 203012 462517 203013
rect 462451 202948 462452 203012
rect 462516 202948 462517 203012
rect 462451 202947 462517 202948
rect 462454 200970 462514 202947
rect 462432 200910 462514 200970
rect 451920 200757 452210 200817
rect 461264 200757 461594 200817
rect 463190 200817 463250 203219
rect 463555 203012 463621 203013
rect 463555 202948 463556 203012
rect 463620 202948 463621 203012
rect 463555 202947 463621 202948
rect 463558 201650 463618 202947
rect 463558 201590 463630 201650
rect 463570 200940 463630 201590
rect 464478 200970 464538 204035
rect 464659 203420 464725 203421
rect 464659 203356 464660 203420
rect 464724 203356 464725 203420
rect 464659 203355 464725 203356
rect 464662 201650 464722 203355
rect 464662 201590 464798 201650
rect 464478 200910 464644 200970
rect 464738 200940 464798 201590
rect 465766 200910 465826 204035
rect 467051 203284 467117 203285
rect 467051 203220 467052 203284
rect 467116 203220 467117 203284
rect 467051 203219 467117 203220
rect 465947 203012 466013 203013
rect 465947 202948 465948 203012
rect 466012 202948 466013 203012
rect 465947 202947 466013 202948
rect 465950 200970 466010 202947
rect 467054 201650 467114 203219
rect 467235 203012 467301 203013
rect 467235 202948 467236 203012
rect 467300 202948 467301 203012
rect 467235 202947 467301 202948
rect 465936 200910 466010 200970
rect 466950 201590 467114 201650
rect 466950 200940 467010 201590
rect 467238 200970 467298 202947
rect 468158 201650 468218 204171
rect 469259 204100 469325 204101
rect 469259 204036 469260 204100
rect 469324 204036 469325 204100
rect 469259 204035 469325 204036
rect 468523 203012 468589 203013
rect 468523 202948 468524 203012
rect 468588 202948 468589 203012
rect 468523 202947 468589 202948
rect 467104 200910 467298 200970
rect 468118 201590 468218 201650
rect 468118 200940 468178 201590
rect 468526 200817 468586 202947
rect 469262 200910 469322 204035
rect 469443 203420 469509 203421
rect 469443 203356 469444 203420
rect 469508 203356 469509 203420
rect 469443 203355 469509 203356
rect 469446 200970 469506 203355
rect 470366 201650 470426 204171
rect 476067 204100 476133 204101
rect 476067 204036 476068 204100
rect 476132 204036 476133 204100
rect 476067 204035 476133 204036
rect 477539 204100 477605 204101
rect 477539 204036 477540 204100
rect 477604 204036 477605 204100
rect 477539 204035 477605 204036
rect 483427 204100 483493 204101
rect 483427 204036 483428 204100
rect 483492 204036 483493 204100
rect 483427 204035 483493 204036
rect 474227 203556 474293 203557
rect 474227 203492 474228 203556
rect 474292 203492 474293 203556
rect 474227 203491 474293 203492
rect 471099 203284 471165 203285
rect 471099 203220 471100 203284
rect 471164 203220 471165 203284
rect 471099 203219 471165 203220
rect 471651 203284 471717 203285
rect 471651 203220 471652 203284
rect 471716 203220 471717 203284
rect 471651 203219 471717 203220
rect 472755 203284 472821 203285
rect 472755 203220 472756 203284
rect 472820 203220 472821 203284
rect 472755 203219 472821 203220
rect 472939 203284 473005 203285
rect 472939 203220 472940 203284
rect 473004 203220 473005 203284
rect 472939 203219 473005 203220
rect 473675 203284 473741 203285
rect 473675 203220 473676 203284
rect 473740 203220 473741 203284
rect 473675 203219 473741 203220
rect 470366 201590 470514 201650
rect 469440 200910 469506 200970
rect 470454 200940 470514 201590
rect 471102 200970 471162 203219
rect 471654 201650 471714 203219
rect 471835 203012 471901 203013
rect 471835 202948 471836 203012
rect 471900 202948 471901 203012
rect 471835 202947 471901 202948
rect 470608 200910 471162 200970
rect 471622 201590 471714 201650
rect 471838 201650 471898 202947
rect 471838 201590 472082 201650
rect 471622 200940 471682 201590
rect 472022 200817 472082 201590
rect 472758 200970 472818 203219
rect 472758 200910 472820 200970
rect 472942 200910 473002 203219
rect 473678 200970 473738 203219
rect 474230 200970 474290 203491
rect 474963 203284 475029 203285
rect 474963 203220 474964 203284
rect 475028 203220 475029 203284
rect 474963 203219 475029 203220
rect 473678 200910 473988 200970
rect 474112 200910 474290 200970
rect 474966 200970 475026 203219
rect 475515 203012 475581 203013
rect 475515 202948 475516 203012
rect 475580 202948 475581 203012
rect 475515 202947 475581 202948
rect 474966 200910 475156 200970
rect 475518 200817 475578 202947
rect 476070 200970 476130 204035
rect 476435 203012 476501 203013
rect 476435 202948 476436 203012
rect 476500 202948 476501 203012
rect 476435 202947 476501 202948
rect 476070 200910 476324 200970
rect 476438 200910 476498 202947
rect 477542 201514 477602 204035
rect 480667 203556 480733 203557
rect 480667 203492 480668 203556
rect 480732 203492 480733 203556
rect 480667 203491 480733 203492
rect 478091 203420 478157 203421
rect 478091 203356 478092 203420
rect 478156 203356 478157 203420
rect 478091 203355 478157 203356
rect 479195 203420 479261 203421
rect 479195 203356 479196 203420
rect 479260 203356 479261 203420
rect 479195 203355 479261 203356
rect 477723 203284 477789 203285
rect 477723 203220 477724 203284
rect 477788 203220 477789 203284
rect 477723 203219 477789 203220
rect 477462 201454 477602 201514
rect 477462 200940 477522 201454
rect 477726 200970 477786 203219
rect 477616 200910 477786 200970
rect 478094 200970 478154 203355
rect 478643 203012 478709 203013
rect 478643 202948 478644 203012
rect 478708 202948 478709 203012
rect 478643 202947 478709 202948
rect 478646 201514 478706 202947
rect 478646 201454 478814 201514
rect 478094 200910 478660 200970
rect 478754 200940 478814 201454
rect 479198 200970 479258 203355
rect 479931 203284 479997 203285
rect 479931 203220 479932 203284
rect 479996 203220 479997 203284
rect 479931 203219 479997 203220
rect 479198 200910 479828 200970
rect 479934 200910 479994 203219
rect 480670 200970 480730 203491
rect 482139 203284 482205 203285
rect 482139 203220 482140 203284
rect 482204 203220 482205 203284
rect 482139 203219 482205 203220
rect 481035 203012 481101 203013
rect 481035 202948 481036 203012
rect 481100 202948 481101 203012
rect 481035 202947 481101 202948
rect 481771 203012 481837 203013
rect 481771 202948 481772 203012
rect 481836 202948 481837 203012
rect 481771 202947 481837 202948
rect 481038 201514 481098 202947
rect 481038 201454 481150 201514
rect 480670 200910 480996 200970
rect 481090 200940 481150 201454
rect 481774 200970 481834 202947
rect 482142 201514 482202 203219
rect 483059 203012 483125 203013
rect 483059 202948 483060 203012
rect 483124 202948 483125 203012
rect 483059 202947 483125 202948
rect 482142 201454 482318 201514
rect 481774 200910 482164 200970
rect 482258 200940 482318 201454
rect 483062 200970 483122 202947
rect 483062 200910 483332 200970
rect 483430 200910 483490 204035
rect 484350 200970 484410 204171
rect 486371 204100 486437 204101
rect 486371 204036 486372 204100
rect 486436 204036 486437 204100
rect 486371 204035 486437 204036
rect 485819 203828 485885 203829
rect 485819 203764 485820 203828
rect 485884 203764 485885 203828
rect 485819 203763 485885 203764
rect 484531 203556 484597 203557
rect 484531 203492 484532 203556
rect 484596 203492 484597 203556
rect 484531 203491 484597 203492
rect 484534 201514 484594 203491
rect 484534 201454 484654 201514
rect 484350 200910 484500 200970
rect 484594 200940 484654 201454
rect 485822 200970 485882 203763
rect 485792 200910 485882 200970
rect 486374 200970 486434 204035
rect 490235 203964 490301 203965
rect 490235 203900 490236 203964
rect 490300 203900 490301 203964
rect 490235 203899 490301 203900
rect 487475 203692 487541 203693
rect 487475 203628 487476 203692
rect 487540 203628 487541 203692
rect 487475 203627 487541 203628
rect 487478 200970 487538 203627
rect 488579 203420 488645 203421
rect 488579 203356 488580 203420
rect 488644 203356 488645 203420
rect 488579 203355 488645 203356
rect 488582 200970 488642 203355
rect 490238 200970 490298 203899
rect 492811 203148 492877 203149
rect 492811 203084 492812 203148
rect 492876 203084 492877 203148
rect 492811 203083 492877 203084
rect 492814 200970 492874 203083
rect 486374 200910 486960 200970
rect 487478 200910 488128 200970
rect 488582 200910 489296 200970
rect 490238 200910 490464 200970
rect 492814 200910 493463 200970
rect 463190 200757 463476 200817
rect 468272 200757 468586 200817
rect 471776 200757 472082 200817
rect 475280 200757 475578 200817
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 420482 182454 420802 182476
rect 420482 182218 420524 182454
rect 420760 182218 420802 182454
rect 420482 182134 420802 182218
rect 420482 181898 420524 182134
rect 420760 181898 420802 182134
rect 420482 181876 420802 181898
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 420034 164454 420358 164476
rect 420034 164218 420078 164454
rect 420314 164218 420358 164454
rect 420034 164134 420358 164218
rect 420034 163898 420078 164134
rect 420314 163898 420358 164134
rect 420034 163876 420358 163898
rect 420482 146454 420802 146476
rect 420482 146218 420524 146454
rect 420760 146218 420802 146454
rect 420482 146134 420802 146218
rect 420482 145898 420524 146134
rect 420760 145898 420802 146134
rect 420482 145876 420802 145898
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 420034 128454 420358 128476
rect 420034 128218 420078 128454
rect 420314 128218 420358 128454
rect 420034 128134 420358 128218
rect 420034 127898 420078 128134
rect 420314 127898 420358 128134
rect 420034 127876 420358 127898
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 423693 110130 424242 110190
rect 424182 109037 424242 110130
rect 428046 110130 428688 110190
rect 504804 110134 505404 110218
rect 428046 109037 428106 110130
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 424179 109036 424245 109037
rect 424179 108972 424180 109036
rect 424244 108972 424245 109036
rect 424179 108971 424245 108972
rect 428043 109036 428109 109037
rect 428043 108972 428044 109036
rect 428108 108972 428109 109036
rect 428043 108971 428109 108972
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 96054 419004 107000
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 99654 422604 107000
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 103254 426204 107000
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 74454 433404 107000
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 78054 437004 107000
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 81654 440604 107000
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 85254 444204 107000
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 92454 451404 107000
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 96054 455004 107000
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 99654 458604 107000
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 103254 462204 107000
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 74454 469404 107000
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 78054 473004 107000
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 81654 476604 107000
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 85254 480204 107000
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 92454 487404 107000
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 96054 491004 107000
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 99654 494604 107000
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 103254 498204 107000
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 222054 509004 237000
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 225654 512604 237000
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 229254 516204 237000
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 520230 64837 520290 472635
rect 520411 466308 520477 466309
rect 520411 466244 520412 466308
rect 520476 466244 520477 466308
rect 520411 466243 520477 466244
rect 520414 108901 520474 466243
rect 520598 384165 520658 700707
rect 520779 700500 520845 700501
rect 520779 700436 520780 700500
rect 520844 700436 520845 700500
rect 520779 700435 520845 700436
rect 520782 390557 520842 700435
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 520963 667996 521029 667997
rect 520963 667932 520964 667996
rect 521028 667932 521029 667996
rect 520963 667931 521029 667932
rect 520966 396813 521026 667931
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 483000 523404 487898
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 522803 476916 522869 476917
rect 522803 476852 522804 476916
rect 522868 476852 522869 476916
rect 522803 476851 522869 476852
rect 521699 474740 521765 474741
rect 521699 474676 521700 474740
rect 521764 474676 521765 474740
rect 521699 474675 521765 474676
rect 521331 468756 521397 468757
rect 521331 468692 521332 468756
rect 521396 468692 521397 468756
rect 521331 468691 521397 468692
rect 521147 468620 521213 468621
rect 521147 468556 521148 468620
rect 521212 468556 521213 468620
rect 521147 468555 521213 468556
rect 521150 465629 521210 468555
rect 521147 465628 521213 465629
rect 521147 465564 521148 465628
rect 521212 465564 521213 465628
rect 521147 465563 521213 465564
rect 521334 465493 521394 468691
rect 521331 465492 521397 465493
rect 521331 465428 521332 465492
rect 521396 465428 521397 465492
rect 521331 465427 521397 465428
rect 521147 437748 521213 437749
rect 521147 437684 521148 437748
rect 521212 437684 521213 437748
rect 521147 437683 521213 437684
rect 521150 435165 521210 437683
rect 521147 435164 521213 435165
rect 521147 435100 521148 435164
rect 521212 435100 521213 435164
rect 521147 435099 521213 435100
rect 521147 429860 521213 429861
rect 521147 429796 521148 429860
rect 521212 429796 521213 429860
rect 521147 429795 521213 429796
rect 521150 425101 521210 429795
rect 521147 425100 521213 425101
rect 521147 425036 521148 425100
rect 521212 425036 521213 425100
rect 521147 425035 521213 425036
rect 520963 396812 521029 396813
rect 520963 396748 520964 396812
rect 521028 396748 521029 396812
rect 520963 396747 521029 396748
rect 520779 390556 520845 390557
rect 520779 390492 520780 390556
rect 520844 390492 520845 390556
rect 520779 390491 520845 390492
rect 520595 384164 520661 384165
rect 520595 384100 520596 384164
rect 520660 384100 520661 384164
rect 520595 384099 520661 384100
rect 520411 108900 520477 108901
rect 520411 108836 520412 108900
rect 520476 108836 520477 108900
rect 520411 108835 520477 108836
rect 520227 64836 520293 64837
rect 520227 64772 520228 64836
rect 520292 64772 520293 64836
rect 520227 64771 520293 64772
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 521702 35869 521762 474675
rect 521883 470524 521949 470525
rect 521883 470460 521884 470524
rect 521948 470460 521949 470524
rect 521883 470459 521949 470460
rect 521886 50965 521946 470459
rect 522067 468484 522133 468485
rect 522067 468420 522068 468484
rect 522132 468420 522133 468484
rect 522067 468419 522133 468420
rect 522070 80069 522130 468419
rect 522251 464268 522317 464269
rect 522251 464204 522252 464268
rect 522316 464204 522317 464268
rect 522251 464203 522317 464204
rect 522254 93805 522314 464203
rect 522435 462092 522501 462093
rect 522435 462028 522436 462092
rect 522500 462028 522501 462092
rect 522435 462027 522501 462028
rect 522438 200701 522498 462027
rect 522619 457876 522685 457877
rect 522619 457812 522620 457876
rect 522684 457812 522685 457876
rect 522619 457811 522685 457812
rect 522622 200837 522682 457811
rect 522806 237149 522866 476851
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 522803 237148 522869 237149
rect 522803 237084 522804 237148
rect 522868 237084 522869 237148
rect 522803 237083 522869 237084
rect 522804 236454 523404 237000
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522619 200836 522685 200837
rect 522619 200772 522620 200836
rect 522684 200772 522685 200836
rect 522619 200771 522685 200772
rect 522435 200700 522501 200701
rect 522435 200636 522436 200700
rect 522500 200636 522501 200700
rect 522435 200635 522501 200636
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522251 93804 522317 93805
rect 522251 93740 522252 93804
rect 522316 93740 522317 93804
rect 522251 93739 522317 93740
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522067 80068 522133 80069
rect 522067 80004 522068 80068
rect 522132 80004 522133 80068
rect 522067 80003 522133 80004
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 521883 50964 521949 50965
rect 521883 50900 521884 50964
rect 521948 50900 521949 50964
rect 521883 50899 521949 50900
rect 521699 35868 521765 35869
rect 521699 35804 521700 35868
rect 521764 35804 521765 35868
rect 521699 35803 521765 35804
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 542491 684452 542557 684453
rect 542491 684388 542492 684452
rect 542556 684388 542557 684452
rect 542491 684387 542557 684388
rect 542494 678877 542554 684387
rect 542491 678876 542557 678877
rect 542491 678812 542492 678876
rect 542556 678812 542557 678876
rect 542491 678811 542557 678812
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 376982 596218 377218 596454
rect 376982 595898 377218 596134
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 376536 578218 376772 578454
rect 376536 577898 376772 578134
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 376982 560218 377218 560454
rect 376982 559898 377218 560134
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 376536 542218 376772 542454
rect 376536 541898 376772 542134
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 376982 524218 377218 524454
rect 376982 523898 377218 524134
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 496982 596218 497218 596454
rect 496982 595898 497218 596134
rect 496536 578218 496772 578454
rect 496536 577898 496772 578134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 496982 560218 497218 560454
rect 496982 559898 497218 560134
rect 496536 542218 496772 542454
rect 496536 541898 496772 542134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 496982 524218 497218 524454
rect 496982 523898 497218 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 284250 470218 284486 470454
rect 284250 469898 284486 470134
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 299610 452218 299846 452454
rect 299610 451898 299846 452134
rect 284250 434218 284486 434454
rect 284250 433898 284486 434134
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 299610 416218 299846 416454
rect 299610 415898 299846 416134
rect 284250 398218 284486 398454
rect 284250 397898 284486 398134
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 299610 380218 299846 380454
rect 299610 379898 299846 380134
rect 284250 362218 284486 362454
rect 284250 361898 284486 362134
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 299610 344218 299846 344454
rect 299610 343898 299846 344134
rect 284250 326218 284486 326454
rect 284250 325898 284486 326134
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 299610 308218 299846 308454
rect 299610 307898 299846 308134
rect 284250 290218 284486 290454
rect 284250 289898 284486 290134
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 299610 272218 299846 272454
rect 299610 271898 299846 272134
rect 284250 254218 284486 254454
rect 284250 253898 284486 254134
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 300524 182218 300760 182454
rect 300524 181898 300760 182134
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 300078 164218 300314 164454
rect 300078 163898 300314 164134
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 300524 146218 300760 146454
rect 300524 145898 300760 146134
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 300078 128218 300314 128454
rect 300078 127898 300314 128134
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 420524 182218 420760 182454
rect 420524 181898 420760 182134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 420078 164218 420314 164454
rect 420078 163898 420314 164134
rect 420524 146218 420760 146454
rect 420524 145898 420760 146134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 420078 128218 420314 128454
rect 420078 127898 420314 128134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 396804 614476 397404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 396986 614454
rect 397222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 396986 614134
rect 397222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 396804 613874 397404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 389604 607276 390204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 389786 607254
rect 390022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 389786 606934
rect 390022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 389604 606674 390204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 386004 603676 386604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 386186 603654
rect 386422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 386186 603334
rect 386422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 386004 603074 386604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 382404 600076 383004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 382586 600054
rect 382822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 382586 599734
rect 382822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 382404 599474 383004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 376938 596476 377262 596478
rect 414804 596476 415404 596478
rect 496938 596476 497262 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 376982 596454
rect 377218 596218 414986 596454
rect 415222 596218 496982 596454
rect 497218 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 376982 596134
rect 377218 595898 414986 596134
rect 415222 595898 496982 596134
rect 497218 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 376938 595874 377262 595876
rect 414804 595874 415404 595876
rect 496938 595874 497262 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 407604 589276 408204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 407786 589254
rect 408022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 407786 588934
rect 408022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 407604 588674 408204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 404004 585676 404604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 404186 585654
rect 404422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 404186 585334
rect 404422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 404004 585074 404604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 400404 582076 401004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 400586 582054
rect 400822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 400586 581734
rect 400822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 400404 581474 401004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 376494 578476 376814 578478
rect 396804 578476 397404 578478
rect 496494 578476 496814 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 376536 578454
rect 376772 578218 396986 578454
rect 397222 578218 496536 578454
rect 496772 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 376536 578134
rect 376772 577898 396986 578134
rect 397222 577898 496536 578134
rect 496772 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 376494 577874 376814 577876
rect 396804 577874 397404 577876
rect 496494 577874 496814 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 389604 571276 390204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 389786 571254
rect 390022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 389786 570934
rect 390022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 389604 570674 390204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 386004 567676 386604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 386186 567654
rect 386422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 386186 567334
rect 386422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 386004 567074 386604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 382404 564076 383004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 382586 564054
rect 382822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 382586 563734
rect 382822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 382404 563474 383004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 376938 560476 377262 560478
rect 414804 560476 415404 560478
rect 496938 560476 497262 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 376982 560454
rect 377218 560218 414986 560454
rect 415222 560218 496982 560454
rect 497218 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 376982 560134
rect 377218 559898 414986 560134
rect 415222 559898 496982 560134
rect 497218 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 376938 559874 377262 559876
rect 414804 559874 415404 559876
rect 496938 559874 497262 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 407604 553276 408204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 407786 553254
rect 408022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 407786 552934
rect 408022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 407604 552674 408204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 404004 549676 404604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 404186 549654
rect 404422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 404186 549334
rect 404422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 404004 549074 404604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 400404 546076 401004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 400586 546054
rect 400822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 400586 545734
rect 400822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 400404 545474 401004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 376494 542476 376814 542478
rect 396804 542476 397404 542478
rect 496494 542476 496814 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 376536 542454
rect 376772 542218 396986 542454
rect 397222 542218 496536 542454
rect 496772 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 376536 542134
rect 376772 541898 396986 542134
rect 397222 541898 496536 542134
rect 496772 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 376494 541874 376814 541876
rect 396804 541874 397404 541876
rect 496494 541874 496814 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 389604 535276 390204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 389786 535254
rect 390022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 389786 534934
rect 390022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 389604 534674 390204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 386004 531676 386604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 386186 531654
rect 386422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 386186 531334
rect 386422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 386004 531074 386604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 382404 528076 383004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 382586 528054
rect 382822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 382586 527734
rect 382822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 382404 527474 383004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 376938 524476 377262 524478
rect 414804 524476 415404 524478
rect 496938 524476 497262 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 376982 524454
rect 377218 524218 414986 524454
rect 415222 524218 496982 524454
rect 497218 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 376982 524134
rect 377218 523898 414986 524134
rect 415222 523898 496982 524134
rect 497218 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 376938 523874 377262 523876
rect 414804 523874 415404 523876
rect 496938 523874 497262 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 407604 517276 408204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 407786 517254
rect 408022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 407786 516934
rect 408022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 407604 516674 408204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 284208 470476 284528 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 284250 470454
rect 284486 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 284250 470134
rect 284486 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 284208 469874 284528 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 299568 452476 299888 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 299610 452454
rect 299846 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 299610 452134
rect 299846 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 299568 451874 299888 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 284208 434476 284528 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 284250 434454
rect 284486 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 284250 434134
rect 284486 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 284208 433874 284528 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 299568 416476 299888 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 299610 416454
rect 299846 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 299610 416134
rect 299846 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 299568 415874 299888 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 284208 398476 284528 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 284250 398454
rect 284486 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 284250 398134
rect 284486 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 284208 397874 284528 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 299568 380476 299888 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 299610 380454
rect 299846 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 299610 380134
rect 299846 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 299568 379874 299888 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 284208 362476 284528 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 284250 362454
rect 284486 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 284250 362134
rect 284486 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 284208 361874 284528 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 299568 344476 299888 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 299610 344454
rect 299846 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 299610 344134
rect 299846 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 299568 343874 299888 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 284208 326476 284528 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 284250 326454
rect 284486 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 284250 326134
rect 284486 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 284208 325874 284528 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 299568 308476 299888 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 299610 308454
rect 299846 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 299610 308134
rect 299846 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 299568 307874 299888 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 284208 290476 284528 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 284250 290454
rect 284486 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 284250 290134
rect 284486 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 284208 289874 284528 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 299568 272476 299888 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 299610 272454
rect 299846 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 299610 272134
rect 299846 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 299568 271874 299888 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 284208 254476 284528 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 284250 254454
rect 284486 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 284250 254134
rect 284486 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 284208 253874 284528 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 382404 204076 383004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 382586 204054
rect 382822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 382586 203734
rect 382822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 382404 203474 383004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 414804 200476 415404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 414986 200454
rect 415222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 414986 200134
rect 415222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 414804 199874 415404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 407604 193276 408204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 407786 193254
rect 408022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 407786 192934
rect 408022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 407604 192674 408204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 404004 189676 404604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 404186 189654
rect 404422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 404186 189334
rect 404422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 404004 189074 404604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 400404 186076 401004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 400586 186054
rect 400822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 400586 185734
rect 400822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 400404 185474 401004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 300482 182476 300802 182478
rect 396804 182476 397404 182478
rect 420482 182476 420802 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 300524 182454
rect 300760 182218 396986 182454
rect 397222 182218 420524 182454
rect 420760 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 300524 182134
rect 300760 181898 396986 182134
rect 397222 181898 420524 182134
rect 420760 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 300482 181874 300802 181876
rect 396804 181874 397404 181876
rect 420482 181874 420802 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 389604 175276 390204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 389786 175254
rect 390022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 389786 174934
rect 390022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 389604 174674 390204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 386004 171676 386604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 386186 171654
rect 386422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 386186 171334
rect 386422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 386004 171074 386604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 382404 168076 383004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 382586 168054
rect 382822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 382586 167734
rect 382822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 382404 167474 383004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 300034 164476 300358 164478
rect 414804 164476 415404 164478
rect 420034 164476 420358 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 300078 164454
rect 300314 164218 414986 164454
rect 415222 164218 420078 164454
rect 420314 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 300078 164134
rect 300314 163898 414986 164134
rect 415222 163898 420078 164134
rect 420314 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 300034 163874 300358 163876
rect 414804 163874 415404 163876
rect 420034 163874 420358 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 407604 157276 408204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 407786 157254
rect 408022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 407786 156934
rect 408022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 407604 156674 408204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 404004 153676 404604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 404186 153654
rect 404422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 404186 153334
rect 404422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 404004 153074 404604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 400404 150076 401004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 400586 150054
rect 400822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 400586 149734
rect 400822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 400404 149474 401004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 300482 146476 300802 146478
rect 396804 146476 397404 146478
rect 420482 146476 420802 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 300524 146454
rect 300760 146218 396986 146454
rect 397222 146218 420524 146454
rect 420760 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 300524 146134
rect 300760 145898 396986 146134
rect 397222 145898 420524 146134
rect 420760 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 300482 145874 300802 145876
rect 396804 145874 397404 145876
rect 420482 145874 420802 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 389604 139276 390204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 389786 139254
rect 390022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 389786 138934
rect 390022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 389604 138674 390204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 386004 135676 386604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 386186 135654
rect 386422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 386186 135334
rect 386422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 386004 135074 386604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 382404 132076 383004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 382586 132054
rect 382822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 382586 131734
rect 382822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 382404 131474 383004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 300034 128476 300358 128478
rect 414804 128476 415404 128478
rect 420034 128476 420358 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 300078 128454
rect 300314 128218 414986 128454
rect 415222 128218 420078 128454
rect 420314 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 300078 128134
rect 300314 127898 414986 128134
rect 415222 127898 420078 128134
rect 420314 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 300034 127874 300358 127876
rect 414804 127874 415404 127876
rect 420034 127874 420358 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 407604 121276 408204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 407786 121254
rect 408022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 407786 120934
rect 408022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 407604 120674 408204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 404004 117676 404604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 404186 117654
rect 404422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 404186 117334
rect 404422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 404004 117074 404604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 400404 114076 401004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 400586 114054
rect 400822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 400586 113734
rect 400822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 400404 113474 401004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 396804 110476 397404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 396986 110454
rect 397222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 396986 110134
rect 397222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 396804 109874 397404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use sram_1rw1r_32_256_8_sky130  sram3
timestamp 1608929960
transform -1 0 497296 0 -1 201247
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram2
timestamp 1608929960
transform -1 0 377296 0 -1 201247
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram1
timestamp 1608929960
transform 1 0 420000 0 1 520000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram0
timestamp 1608929960
transform 1 0 300000 0 1 520000
box 0 0 77296 91247
use hs32_core1  core1
timestamp 1608929960
transform 1 0 280000 0 1 240000
box 0 0 240000 240000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 274 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 275 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 276 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 277 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 278 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 279 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 280 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 281 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 282 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 283 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 284 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 285 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 286 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 287 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 288 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 289 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 290 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 291 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 292 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 293 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 294 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 295 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 296 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 297 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 298 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 299 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 300 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 301 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 302 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 303 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 304 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 305 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 306 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 307 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 308 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 309 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 310 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 311 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 312 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 313 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 314 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 315 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 316 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 317 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 318 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 319 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 320 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 321 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 322 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 323 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 324 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 325 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 326 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 327 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 328 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 329 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 330 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 331 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 332 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 333 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 334 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 335 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 336 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 337 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 338 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 339 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 340 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 341 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 342 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 343 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 344 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 345 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 346 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 347 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 348 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 349 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 350 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 351 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 352 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 353 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 354 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 355 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 356 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 357 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 358 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 359 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 360 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 361 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 362 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 363 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 364 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 365 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 366 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 367 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 368 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 369 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 370 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 371 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 372 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 373 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 374 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 375 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 376 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 377 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 378 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 379 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 380 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 381 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 382 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 383 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 384 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 385 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 386 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 387 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 388 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 389 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 390 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 391 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 392 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 393 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 394 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 395 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 396 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 397 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 398 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 399 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 400 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 401 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 402 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 403 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 404 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 405 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 406 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 407 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 408 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 409 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 410 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 411 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 412 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 413 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 414 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 415 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 416 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 417 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 418 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 419 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 420 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 421 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 422 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 423 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 424 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 425 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 426 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 427 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 428 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 429 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 430 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 431 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 432 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 433 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 434 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 435 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 436 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 437 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 438 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 439 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 440 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 441 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 442 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 443 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 444 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 445 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 446 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 447 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 448 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 449 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 450 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 451 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 452 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 453 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 454 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 455 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 456 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 457 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 458 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 459 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 460 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 461 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 462 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 463 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 464 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 465 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 466 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 467 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 468 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 469 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 470 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 471 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 472 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 473 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 474 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 475 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 476 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 477 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 478 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 479 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 480 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 481 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 482 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 483 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 484 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 485 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 486 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 487 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 488 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 489 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 490 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 491 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 492 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 493 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 494 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 495 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 496 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 497 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 498 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 499 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 500 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 501 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 502 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 503 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 504 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 505 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 506 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 507 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 508 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 509 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 510 nsew default input
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 511 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 512 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 513 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 514 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 515 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 516 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 517 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 518 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 519 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 520 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 521 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 522 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 523 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 524 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 525 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 526 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 527 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 528 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 529 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 530 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 531 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 532 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 533 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 534 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 535 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 536 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 537 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 538 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 539 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 540 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 541 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 542 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 543 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 544 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 545 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 546 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 547 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 548 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 549 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 550 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 551 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 552 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 553 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 554 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 555 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 556 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 557 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 558 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 559 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 560 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 561 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 562 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 563 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 564 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 565 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 566 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 567 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 568 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 569 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 570 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 571 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 572 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 573 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 574 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 575 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 576 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 577 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 578 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 579 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 580 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 581 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 582 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 583 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 584 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 585 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 586 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 587 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 588 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 589 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 590 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 591 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 592 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 593 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 594 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 595 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 596 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 597 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 598 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 599 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 600 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 601 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 602 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 603 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 604 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 605 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 606 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 607 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 608 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 609 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 610 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 611 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 612 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 613 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 614 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 615 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 616 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 617 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 618 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 619 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 620 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 621 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 622 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 623 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 624 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 625 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 626 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 627 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 628 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 629 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 630 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 631 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 632 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 633 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 634 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 635 nsew default tristate
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
