magic
tech sky130A
magscale 1 2
timestamp 1608756459
<< metal1 >>
rect 57698 700952 57704 701004
rect 57756 700992 57762 701004
rect 170306 700992 170312 701004
rect 57756 700964 170312 700992
rect 57756 700952 57762 700964
rect 170306 700952 170312 700964
rect 170364 700952 170370 701004
rect 58802 700884 58808 700936
rect 58860 700924 58866 700936
rect 202782 700924 202788 700936
rect 58860 700896 202788 700924
rect 58860 700884 58866 700896
rect 202782 700884 202788 700896
rect 202840 700884 202846 700936
rect 57790 700816 57796 700868
rect 57848 700856 57854 700868
rect 218974 700856 218980 700868
rect 57848 700828 218980 700856
rect 57848 700816 57854 700828
rect 218974 700816 218980 700828
rect 219032 700816 219038 700868
rect 58894 700748 58900 700800
rect 58952 700788 58958 700800
rect 267642 700788 267648 700800
rect 58952 700760 267648 700788
rect 58952 700748 58958 700760
rect 267642 700748 267648 700760
rect 267700 700748 267706 700800
rect 59446 700680 59452 700732
rect 59504 700720 59510 700732
rect 283834 700720 283840 700732
rect 59504 700692 283840 700720
rect 59504 700680 59510 700692
rect 283834 700680 283840 700692
rect 283892 700680 283898 700732
rect 59538 700612 59544 700664
rect 59596 700652 59602 700664
rect 105446 700652 105452 700664
rect 59596 700624 105452 700652
rect 59596 700612 59602 700624
rect 105446 700612 105452 700624
rect 105504 700612 105510 700664
rect 136358 700612 136364 700664
rect 136416 700652 136422 700664
rect 364978 700652 364984 700664
rect 136416 700624 364984 700652
rect 136416 700612 136422 700624
rect 364978 700612 364984 700624
rect 365036 700612 365042 700664
rect 58986 700544 58992 700596
rect 59044 700584 59050 700596
rect 332502 700584 332508 700596
rect 59044 700556 332508 700584
rect 59044 700544 59050 700556
rect 332502 700544 332508 700556
rect 332560 700544 332566 700596
rect 57882 700476 57888 700528
rect 57940 700516 57946 700528
rect 348786 700516 348792 700528
rect 57940 700488 348792 700516
rect 57940 700476 57946 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 59170 700408 59176 700460
rect 59228 700448 59234 700460
rect 397454 700448 397460 700460
rect 59228 700420 397460 700448
rect 59228 700408 59234 700420
rect 397454 700408 397460 700420
rect 397512 700408 397518 700460
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 13078 700380 13084 700392
rect 8168 700352 13084 700380
rect 8168 700340 8174 700352
rect 13078 700340 13084 700352
rect 13136 700340 13142 700392
rect 59078 700340 59084 700392
rect 59136 700380 59142 700392
rect 413646 700380 413652 700392
rect 59136 700352 413652 700380
rect 59136 700340 59142 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 59262 700272 59268 700324
rect 59320 700312 59326 700324
rect 462314 700312 462320 700324
rect 59320 700284 462320 700312
rect 59320 700272 59326 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 58434 700204 58440 700256
rect 58492 700244 58498 700256
rect 89162 700244 89168 700256
rect 58492 700216 89168 700244
rect 58492 700204 58498 700216
rect 89162 700204 89168 700216
rect 89220 700204 89226 700256
rect 136450 700204 136456 700256
rect 136508 700244 136514 700256
rect 235166 700244 235172 700256
rect 136508 700216 235172 700244
rect 136508 700204 136514 700216
rect 235166 700204 235172 700216
rect 235224 700204 235230 700256
rect 58618 700136 58624 700188
rect 58676 700176 58682 700188
rect 154114 700176 154120 700188
rect 58676 700148 154120 700176
rect 58676 700136 58682 700148
rect 154114 700136 154120 700148
rect 154172 700136 154178 700188
rect 58710 700068 58716 700120
rect 58768 700108 58774 700120
rect 137830 700108 137836 700120
rect 58768 700080 137836 700108
rect 58768 700068 58774 700080
rect 137830 700068 137836 700080
rect 137888 700068 137894 700120
rect 58526 700000 58532 700052
rect 58584 700040 58590 700052
rect 72970 700040 72976 700052
rect 58584 700012 72976 700040
rect 58584 700000 58590 700012
rect 72970 700000 72976 700012
rect 73028 700000 73034 700052
rect 40494 699932 40500 699984
rect 40552 699972 40558 699984
rect 42058 699972 42064 699984
rect 40552 699944 42064 699972
rect 40552 699932 40558 699944
rect 42058 699932 42064 699944
rect 42116 699932 42122 699984
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 58158 696940 58164 696992
rect 58216 696980 58222 696992
rect 580166 696980 580172 696992
rect 58216 696952 580172 696980
rect 58216 696940 58222 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 429194 692792 429200 692844
rect 429252 692832 429258 692844
rect 429930 692832 429936 692844
rect 429252 692804 429936 692832
rect 429252 692792 429258 692804
rect 429930 692792 429936 692804
rect 429988 692792 429994 692844
rect 299658 688576 299664 688628
rect 299716 688616 299722 688628
rect 300118 688616 300124 688628
rect 299716 688588 300124 688616
rect 299716 688576 299722 688588
rect 300118 688576 300124 688588
rect 300176 688576 300182 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 299492 685936 301268 685964
rect 59354 685856 59360 685908
rect 59412 685896 59418 685908
rect 299492 685896 299520 685936
rect 59412 685868 299520 685896
rect 301240 685896 301268 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 301240 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 59412 685856 59418 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 299566 684428 299572 684480
rect 299624 684468 299630 684480
rect 299658 684468 299664 684480
rect 299624 684440 299664 684468
rect 299624 684428 299630 684440
rect 299658 684428 299664 684440
rect 299716 684428 299722 684480
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559098 684468 559104 684480
rect 559064 684440 559104 684468
rect 559064 684428 559070 684440
rect 559098 684428 559104 684440
rect 559156 684428 559162 684480
rect 299658 678988 299664 679040
rect 299716 678988 299722 679040
rect 559098 678988 559104 679040
rect 559156 678988 559162 679040
rect 299676 678904 299704 678988
rect 559116 678904 559144 678988
rect 299658 678852 299664 678904
rect 299716 678852 299722 678904
rect 559098 678852 559104 678904
rect 559156 678852 559162 678904
rect 560294 673888 560300 673940
rect 560352 673928 560358 673940
rect 565170 673928 565176 673940
rect 560352 673900 565176 673928
rect 560352 673888 560358 673900
rect 565170 673888 565176 673900
rect 565228 673888 565234 673940
rect 289814 673752 289820 673804
rect 289872 673792 289878 673804
rect 292666 673792 292672 673804
rect 289872 673764 292672 673792
rect 289872 673752 289878 673764
rect 292666 673752 292672 673764
rect 292724 673752 292730 673804
rect 540974 673752 540980 673804
rect 541032 673792 541038 673804
rect 548610 673792 548616 673804
rect 541032 673764 548616 673792
rect 541032 673752 541038 673764
rect 548610 673752 548616 673764
rect 548668 673752 548674 673804
rect 429194 673412 429200 673464
rect 429252 673452 429258 673464
rect 429470 673452 429476 673464
rect 429252 673424 429476 673452
rect 429252 673412 429258 673424
rect 429470 673412 429476 673424
rect 429528 673412 429534 673464
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 21358 667944 21364 667956
rect 3476 667916 21364 667944
rect 3476 667904 3482 667916
rect 21358 667904 21364 667916
rect 21416 667904 21422 667956
rect 299658 666544 299664 666596
rect 299716 666584 299722 666596
rect 299934 666584 299940 666596
rect 299716 666556 299940 666584
rect 299716 666544 299722 666556
rect 299934 666544 299940 666556
rect 299992 666544 299998 666596
rect 559098 666544 559104 666596
rect 559156 666584 559162 666596
rect 559374 666584 559380 666596
rect 559156 666556 559380 666584
rect 559156 666544 559162 666556
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 299658 661716 299664 661768
rect 299716 661756 299722 661768
rect 299934 661756 299940 661768
rect 299716 661728 299940 661756
rect 299716 661716 299722 661728
rect 299934 661716 299940 661728
rect 299992 661716 299998 661768
rect 559098 661716 559104 661768
rect 559156 661756 559162 661768
rect 559374 661756 559380 661768
rect 559156 661728 559380 661756
rect 559156 661716 559162 661728
rect 559374 661716 559380 661728
rect 559432 661716 559438 661768
rect 299658 656888 299664 656940
rect 299716 656928 299722 656940
rect 299750 656928 299756 656940
rect 299716 656900 299756 656928
rect 299716 656888 299722 656900
rect 299750 656888 299756 656900
rect 299808 656888 299814 656940
rect 559098 656888 559104 656940
rect 559156 656928 559162 656940
rect 559190 656928 559196 656940
rect 559156 656900 559196 656928
rect 559156 656888 559162 656900
rect 559190 656888 559196 656900
rect 559248 656888 559254 656940
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 14458 652780 14464 652792
rect 3108 652752 14464 652780
rect 3108 652740 3114 652752
rect 14458 652740 14464 652752
rect 14516 652740 14522 652792
rect 560294 650360 560300 650412
rect 560352 650400 560358 650412
rect 565170 650400 565176 650412
rect 560352 650372 565176 650400
rect 560352 650360 560358 650372
rect 565170 650360 565176 650372
rect 565228 650360 565234 650412
rect 425054 650224 425060 650276
rect 425112 650264 425118 650276
rect 434530 650264 434536 650276
rect 425112 650236 434536 650264
rect 425112 650224 425118 650236
rect 434530 650224 434536 650236
rect 434588 650224 434594 650276
rect 540974 650224 540980 650276
rect 541032 650264 541038 650276
rect 548610 650264 548616 650276
rect 541032 650236 548616 650264
rect 541032 650224 541038 650236
rect 548610 650224 548616 650236
rect 548668 650224 548674 650276
rect 299658 647232 299664 647284
rect 299716 647272 299722 647284
rect 299750 647272 299756 647284
rect 299716 647244 299756 647272
rect 299716 647232 299722 647244
rect 299750 647232 299756 647244
rect 299808 647232 299814 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 299658 640364 299664 640416
rect 299716 640404 299722 640416
rect 299750 640404 299756 640416
rect 299716 640376 299756 640404
rect 299716 640364 299722 640376
rect 299750 640364 299756 640376
rect 299808 640364 299814 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 59630 638936 59636 638988
rect 59688 638976 59694 638988
rect 580166 638976 580172 638988
rect 59688 638948 580172 638976
rect 59688 638936 59694 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 299750 630680 299756 630692
rect 299624 630652 299756 630680
rect 299624 630640 299630 630652
rect 299750 630640 299756 630652
rect 299808 630640 299814 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 560294 626968 560300 627020
rect 560352 627008 560358 627020
rect 565170 627008 565176 627020
rect 560352 626980 565176 627008
rect 560352 626968 560358 626980
rect 565170 626968 565176 626980
rect 565228 626968 565234 627020
rect 289814 626832 289820 626884
rect 289872 626872 289878 626884
rect 292666 626872 292672 626884
rect 289872 626844 292672 626872
rect 289872 626832 289878 626844
rect 292666 626832 292672 626844
rect 292724 626832 292730 626884
rect 425054 626832 425060 626884
rect 425112 626872 425118 626884
rect 427906 626872 427912 626884
rect 425112 626844 427912 626872
rect 425112 626832 425118 626844
rect 427906 626832 427912 626844
rect 427964 626832 427970 626884
rect 540974 626832 540980 626884
rect 541032 626872 541038 626884
rect 548610 626872 548616 626884
rect 541032 626844 548616 626872
rect 541032 626832 541038 626844
rect 548610 626832 548616 626844
rect 548668 626832 548674 626884
rect 4062 623772 4068 623824
rect 4120 623812 4126 623824
rect 4982 623812 4988 623824
rect 4120 623784 4988 623812
rect 4120 623772 4126 623784
rect 4982 623772 4988 623784
rect 5040 623772 5046 623824
rect 429470 618196 429476 618248
rect 429528 618236 429534 618248
rect 429654 618236 429660 618248
rect 429528 618208 429660 618236
rect 429528 618196 429534 618208
rect 429654 618196 429660 618208
rect 429712 618196 429718 618248
rect 559190 618196 559196 618248
rect 559248 618236 559254 618248
rect 559374 618236 559380 618248
rect 559248 618208 559380 618236
rect 559248 618196 559254 618208
rect 559374 618196 559380 618208
rect 559432 618196 559438 618248
rect 299566 611328 299572 611380
rect 299624 611368 299630 611380
rect 299750 611368 299756 611380
rect 299624 611340 299756 611368
rect 299624 611328 299630 611340
rect 299750 611328 299756 611340
rect 299808 611328 299814 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 28258 610008 28264 610020
rect 3476 609980 28264 610008
rect 3476 609968 3482 609980
rect 28258 609968 28264 609980
rect 28316 609968 28322 610020
rect 429286 608608 429292 608660
rect 429344 608648 429350 608660
rect 429654 608648 429660 608660
rect 429344 608620 429660 608648
rect 429344 608608 429350 608620
rect 429654 608608 429660 608620
rect 429712 608608 429718 608660
rect 559098 608540 559104 608592
rect 559156 608580 559162 608592
rect 559466 608580 559472 608592
rect 559156 608552 559472 608580
rect 559156 608540 559162 608552
rect 559466 608540 559472 608552
rect 559524 608540 559530 608592
rect 429194 608472 429200 608524
rect 429252 608512 429258 608524
rect 429286 608512 429292 608524
rect 429252 608484 429292 608512
rect 429252 608472 429258 608484
rect 429286 608472 429292 608484
rect 429344 608472 429350 608524
rect 560294 603440 560300 603492
rect 560352 603480 560358 603492
rect 565170 603480 565176 603492
rect 560352 603452 565176 603480
rect 560352 603440 560358 603452
rect 565170 603440 565176 603452
rect 565228 603440 565234 603492
rect 289814 603304 289820 603356
rect 289872 603344 289878 603356
rect 292666 603344 292672 603356
rect 289872 603316 292672 603344
rect 289872 603304 289878 603316
rect 292666 603304 292672 603316
rect 292724 603304 292730 603356
rect 425054 603304 425060 603356
rect 425112 603344 425118 603356
rect 429930 603344 429936 603356
rect 425112 603316 429936 603344
rect 425112 603304 425118 603316
rect 429930 603304 429936 603316
rect 429988 603304 429994 603356
rect 540974 603304 540980 603356
rect 541032 603344 541038 603356
rect 548610 603344 548616 603356
rect 541032 603316 548616 603344
rect 541032 603304 541038 603316
rect 548610 603304 548616 603316
rect 548668 603304 548674 603356
rect 299658 599020 299664 599072
rect 299716 599060 299722 599072
rect 299842 599060 299848 599072
rect 299716 599032 299848 599060
rect 299716 599020 299722 599032
rect 299842 599020 299848 599032
rect 299900 599020 299906 599072
rect 429194 598952 429200 599004
rect 429252 598992 429258 599004
rect 429378 598992 429384 599004
rect 429252 598964 429384 598992
rect 429252 598952 429258 598964
rect 429378 598952 429384 598964
rect 429436 598952 429442 599004
rect 299658 598884 299664 598936
rect 299716 598924 299722 598936
rect 299842 598924 299848 598936
rect 299716 598896 299848 598924
rect 299716 598884 299722 598896
rect 299842 598884 299848 598896
rect 299900 598884 299906 598936
rect 429194 598816 429200 598868
rect 429252 598856 429258 598868
rect 429378 598856 429384 598868
rect 429252 598828 429384 598856
rect 429252 598816 429258 598828
rect 429378 598816 429384 598828
rect 429436 598816 429442 598868
rect 559190 597524 559196 597576
rect 559248 597564 559254 597576
rect 559374 597564 559380 597576
rect 559248 597536 559380 597564
rect 559248 597524 559254 597536
rect 559374 597524 559380 597536
rect 559432 597524 559438 597576
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 17310 594844 17316 594856
rect 3292 594816 17316 594844
rect 3292 594804 3298 594816
rect 17310 594804 17316 594816
rect 17368 594804 17374 594856
rect 59722 592016 59728 592068
rect 59780 592056 59786 592068
rect 580166 592056 580172 592068
rect 59780 592028 580172 592056
rect 59780 592016 59786 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 299658 589296 299664 589348
rect 299716 589336 299722 589348
rect 299934 589336 299940 589348
rect 299716 589308 299940 589336
rect 299716 589296 299722 589308
rect 299934 589296 299940 589308
rect 299992 589296 299998 589348
rect 429194 589296 429200 589348
rect 429252 589336 429258 589348
rect 429470 589336 429476 589348
rect 429252 589308 429476 589336
rect 429252 589296 429258 589308
rect 429470 589296 429476 589308
rect 429528 589296 429534 589348
rect 559190 589296 559196 589348
rect 559248 589336 559254 589348
rect 559374 589336 559380 589348
rect 559248 589308 559380 589336
rect 559248 589296 559254 589308
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 299934 582468 299940 582480
rect 299860 582440 299940 582468
rect 299860 582344 299888 582440
rect 299934 582428 299940 582440
rect 299992 582428 299998 582480
rect 559374 582468 559380 582480
rect 559300 582440 559380 582468
rect 559300 582344 559328 582440
rect 559374 582428 559380 582440
rect 559432 582428 559438 582480
rect 299842 582292 299848 582344
rect 299900 582292 299906 582344
rect 559282 582292 559288 582344
rect 559340 582292 559346 582344
rect 58342 579640 58348 579692
rect 58400 579680 58406 579692
rect 580166 579680 580172 579692
rect 58400 579652 580172 579680
rect 58400 579640 58406 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 429378 579572 429384 579624
rect 429436 579612 429442 579624
rect 429562 579612 429568 579624
rect 429436 579584 429568 579612
rect 429436 579572 429442 579584
rect 429562 579572 429568 579584
rect 429620 579572 429626 579624
rect 429378 569916 429384 569968
rect 429436 569956 429442 569968
rect 429654 569956 429660 569968
rect 429436 569928 429660 569956
rect 429436 569916 429442 569928
rect 429654 569916 429660 569928
rect 429712 569916 429718 569968
rect 429470 563728 429476 563780
rect 429528 563768 429534 563780
rect 429654 563768 429660 563780
rect 429528 563740 429660 563768
rect 429528 563728 429534 563740
rect 429654 563728 429660 563740
rect 429712 563728 429718 563780
rect 299566 563116 299572 563168
rect 299624 563116 299630 563168
rect 559006 563116 559012 563168
rect 559064 563116 559070 563168
rect 299584 563032 299612 563116
rect 559024 563032 559052 563116
rect 299566 562980 299572 563032
rect 299624 562980 299630 563032
rect 559006 562980 559012 563032
rect 559064 562980 559070 563032
rect 429286 560192 429292 560244
rect 429344 560232 429350 560244
rect 429470 560232 429476 560244
rect 429344 560204 429476 560232
rect 429344 560192 429350 560204
rect 429470 560192 429476 560204
rect 429528 560192 429534 560244
rect 58250 556180 58256 556232
rect 58308 556220 58314 556232
rect 580166 556220 580172 556232
rect 58308 556192 580172 556220
rect 58308 556180 58314 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 263778 554004 263784 554056
rect 263836 554044 263842 554056
rect 378502 554044 378508 554056
rect 263836 554016 378508 554044
rect 263836 554004 263842 554016
rect 378502 554004 378508 554016
rect 378560 554004 378566 554056
rect 507854 554004 507860 554056
rect 507912 554044 507918 554056
rect 513374 554044 513380 554056
rect 507912 554016 513380 554044
rect 507912 554004 507918 554016
rect 513374 554004 513380 554016
rect 513432 554004 513438 554056
rect 299566 553500 299572 553512
rect 299492 553472 299572 553500
rect 133690 553392 133696 553444
rect 133748 553432 133754 553444
rect 139578 553432 139584 553444
rect 133748 553404 139584 553432
rect 133748 553392 133754 553404
rect 139578 553392 139584 553404
rect 139636 553432 139642 553444
rect 259178 553432 259184 553444
rect 139636 553404 259184 553432
rect 139636 553392 139642 553404
rect 259178 553392 259184 553404
rect 259236 553432 259242 553444
rect 263778 553432 263784 553444
rect 259236 553404 263784 553432
rect 259236 553392 259242 553404
rect 263778 553392 263784 553404
rect 263836 553392 263842 553444
rect 299492 553376 299520 553472
rect 299566 553460 299572 553472
rect 299624 553460 299630 553512
rect 378502 553392 378508 553444
rect 378560 553432 378566 553444
rect 382918 553432 382924 553444
rect 378560 553404 382924 553432
rect 378560 553392 378566 553404
rect 382918 553392 382924 553404
rect 382976 553432 382982 553444
rect 389358 553432 389364 553444
rect 382976 553404 389364 553432
rect 382976 553392 382982 553404
rect 389358 553392 389364 553404
rect 389416 553432 389422 553444
rect 507854 553432 507860 553444
rect 389416 553404 507860 553432
rect 389416 553392 389422 553404
rect 507854 553392 507860 553404
rect 507912 553392 507918 553444
rect 558914 553392 558920 553444
rect 558972 553432 558978 553444
rect 558972 553404 559052 553432
rect 558972 553392 558978 553404
rect 559024 553376 559052 553404
rect 299474 553324 299480 553376
rect 299532 553324 299538 553376
rect 559006 553324 559012 553376
rect 559064 553324 559070 553376
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 32398 552072 32404 552084
rect 3200 552044 32404 552072
rect 3200 552032 3206 552044
rect 32398 552032 32404 552044
rect 32456 552032 32462 552084
rect 429286 550604 429292 550656
rect 429344 550644 429350 550656
rect 429562 550644 429568 550656
rect 429344 550616 429568 550644
rect 429344 550604 429350 550616
rect 429562 550604 429568 550616
rect 429620 550604 429626 550656
rect 558914 550604 558920 550656
rect 558972 550644 558978 550656
rect 559006 550644 559012 550656
rect 558972 550616 559012 550644
rect 558972 550604 558978 550616
rect 559006 550604 559012 550616
rect 559064 550604 559070 550656
rect 139394 550264 139400 550316
rect 139452 550304 139458 550316
rect 266446 550304 266452 550316
rect 139452 550276 266452 550304
rect 139452 550264 139458 550276
rect 266446 550264 266452 550276
rect 266504 550264 266510 550316
rect 302234 550264 302240 550316
rect 302292 550304 302298 550316
rect 389174 550304 389180 550316
rect 302292 550276 389180 550304
rect 302292 550264 302298 550276
rect 389174 550264 389180 550276
rect 389232 550304 389238 550316
rect 516410 550304 516416 550316
rect 389232 550276 516416 550304
rect 389232 550264 389238 550276
rect 516410 550264 516416 550276
rect 516468 550264 516474 550316
rect 270402 549244 270408 549296
rect 270460 549284 270466 549296
rect 302234 549284 302240 549296
rect 270460 549256 302240 549284
rect 270460 549244 270466 549256
rect 302234 549244 302240 549256
rect 302292 549244 302298 549296
rect 299474 549176 299480 549228
rect 299532 549216 299538 549228
rect 299566 549216 299572 549228
rect 299532 549188 299572 549216
rect 299532 549176 299538 549188
rect 299566 549176 299572 549188
rect 299624 549176 299630 549228
rect 150342 546456 150348 546508
rect 150400 546496 150406 546508
rect 187694 546496 187700 546508
rect 150400 546468 187700 546496
rect 150400 546456 150406 546468
rect 187694 546456 187700 546468
rect 187752 546456 187758 546508
rect 399478 546456 399484 546508
rect 399536 546496 399542 546508
rect 437474 546496 437480 546508
rect 399536 546468 437480 546496
rect 399536 546456 399542 546468
rect 437474 546456 437480 546468
rect 437532 546456 437538 546508
rect 147582 545096 147588 545148
rect 147640 545136 147646 545148
rect 187694 545136 187700 545148
rect 147640 545108 187700 545136
rect 147640 545096 147646 545108
rect 187694 545096 187700 545108
rect 187752 545096 187758 545148
rect 304442 545096 304448 545148
rect 304500 545136 304506 545148
rect 307662 545136 307668 545148
rect 304500 545108 307668 545136
rect 304500 545096 304506 545108
rect 307662 545096 307668 545108
rect 307720 545096 307726 545148
rect 398098 545096 398104 545148
rect 398156 545136 398162 545148
rect 437474 545136 437480 545148
rect 398156 545108 437480 545136
rect 398156 545096 398162 545108
rect 437474 545096 437480 545108
rect 437532 545096 437538 545148
rect 144822 543736 144828 543788
rect 144880 543776 144886 543788
rect 187694 543776 187700 543788
rect 144880 543748 187700 543776
rect 144880 543736 144886 543748
rect 187694 543736 187700 543748
rect 187752 543736 187758 543788
rect 299566 543736 299572 543788
rect 299624 543736 299630 543788
rect 395338 543736 395344 543788
rect 395396 543776 395402 543788
rect 437474 543776 437480 543788
rect 395396 543748 437480 543776
rect 395396 543736 395402 543748
rect 437474 543736 437480 543748
rect 437532 543736 437538 543788
rect 558914 543736 558920 543788
rect 558972 543736 558978 543788
rect 299584 543652 299612 543736
rect 299566 543600 299572 543652
rect 299624 543600 299630 543652
rect 558932 543640 558960 543736
rect 559006 543640 559012 543652
rect 558932 543612 559012 543640
rect 559006 543600 559012 543612
rect 559064 543600 559070 543652
rect 143442 542376 143448 542428
rect 143500 542416 143506 542428
rect 187694 542416 187700 542428
rect 143500 542388 187700 542416
rect 143500 542376 143506 542388
rect 187694 542376 187700 542388
rect 187752 542376 187758 542428
rect 304350 542376 304356 542428
rect 304408 542416 304414 542428
rect 307202 542416 307208 542428
rect 304408 542388 307208 542416
rect 304408 542376 304414 542388
rect 307202 542376 307208 542388
rect 307260 542376 307266 542428
rect 393958 542376 393964 542428
rect 394016 542416 394022 542428
rect 437474 542416 437480 542428
rect 394016 542388 437480 542416
rect 394016 542376 394022 542388
rect 437474 542376 437480 542388
rect 437532 542376 437538 542428
rect 140682 539656 140688 539708
rect 140740 539696 140746 539708
rect 187786 539696 187792 539708
rect 140740 539668 187792 539696
rect 140740 539656 140746 539668
rect 187786 539656 187792 539668
rect 187844 539656 187850 539708
rect 392578 539656 392584 539708
rect 392636 539696 392642 539708
rect 437566 539696 437572 539708
rect 392636 539668 437572 539696
rect 392636 539656 392642 539668
rect 437566 539656 437572 539668
rect 437624 539656 437630 539708
rect 139302 539588 139308 539640
rect 139360 539628 139366 539640
rect 187694 539628 187700 539640
rect 139360 539600 187700 539628
rect 139360 539588 139366 539600
rect 187694 539588 187700 539600
rect 187752 539588 187758 539640
rect 304258 539588 304264 539640
rect 304316 539628 304322 539640
rect 307662 539628 307668 539640
rect 304316 539600 307668 539628
rect 304316 539588 304322 539600
rect 307662 539588 307668 539600
rect 307720 539588 307726 539640
rect 391198 539588 391204 539640
rect 391256 539628 391262 539640
rect 437474 539628 437480 539640
rect 391256 539600 437480 539628
rect 391256 539588 391262 539600
rect 437474 539588 437480 539600
rect 437532 539588 437538 539640
rect 388438 536800 388444 536852
rect 388496 536840 388502 536852
rect 437474 536840 437480 536852
rect 388496 536812 437480 536840
rect 388496 536800 388502 536812
rect 437474 536800 437480 536812
rect 437532 536800 437538 536852
rect 559006 534012 559012 534064
rect 559064 534052 559070 534064
rect 559190 534052 559196 534064
rect 559064 534024 559196 534052
rect 559064 534012 559070 534024
rect 559190 534012 559196 534024
rect 559248 534012 559254 534064
rect 299566 531292 299572 531344
rect 299624 531332 299630 531344
rect 299658 531332 299664 531344
rect 299624 531304 299664 531332
rect 299624 531292 299630 531304
rect 299658 531292 299664 531304
rect 299716 531292 299722 531344
rect 429194 531292 429200 531344
rect 429252 531332 429258 531344
rect 429470 531332 429476 531344
rect 429252 531304 429476 531332
rect 429252 531292 429258 531304
rect 429470 531292 429476 531304
rect 429528 531292 429534 531344
rect 429470 524424 429476 524476
rect 429528 524424 429534 524476
rect 559190 524424 559196 524476
rect 559248 524424 559254 524476
rect 429488 524396 429516 524424
rect 429562 524396 429568 524408
rect 429488 524368 429568 524396
rect 429562 524356 429568 524368
rect 429620 524356 429626 524408
rect 559208 524396 559236 524424
rect 559282 524396 559288 524408
rect 559208 524368 559288 524396
rect 559282 524356 559288 524368
rect 559340 524356 559346 524408
rect 299474 521636 299480 521688
rect 299532 521676 299538 521688
rect 299750 521676 299756 521688
rect 299532 521648 299756 521676
rect 299532 521636 299538 521648
rect 299750 521636 299756 521648
rect 299808 521636 299814 521688
rect 429378 511980 429384 512032
rect 429436 512020 429442 512032
rect 429654 512020 429660 512032
rect 429436 511992 429660 512020
rect 429436 511980 429442 511992
rect 429654 511980 429660 511992
rect 429712 511980 429718 512032
rect 559098 511980 559104 512032
rect 559156 512020 559162 512032
rect 559374 512020 559380 512032
rect 559156 511992 559380 512020
rect 559156 511980 559162 511992
rect 559374 511980 559380 511992
rect 559432 511980 559438 512032
rect 299474 502324 299480 502376
rect 299532 502364 299538 502376
rect 299750 502364 299756 502376
rect 299532 502336 299756 502364
rect 299532 502324 299538 502336
rect 299750 502324 299756 502336
rect 299808 502324 299814 502376
rect 429470 502324 429476 502376
rect 429528 502364 429534 502376
rect 429654 502364 429660 502376
rect 429528 502336 429660 502364
rect 429528 502324 429534 502336
rect 429654 502324 429660 502336
rect 429712 502324 429718 502376
rect 559190 502324 559196 502376
rect 559248 502364 559254 502376
rect 559374 502364 559380 502376
rect 559248 502336 559380 502364
rect 559248 502324 559254 502336
rect 559374 502324 559380 502336
rect 559432 502324 559438 502376
rect 299474 492600 299480 492652
rect 299532 492640 299538 492652
rect 299658 492640 299664 492652
rect 299532 492612 299664 492640
rect 299532 492600 299538 492612
rect 299658 492600 299664 492612
rect 299716 492600 299722 492652
rect 559098 492600 559104 492652
rect 559156 492640 559162 492652
rect 559190 492640 559196 492652
rect 559156 492612 559196 492640
rect 559156 492600 559162 492612
rect 559190 492600 559196 492612
rect 559248 492600 559254 492652
rect 429470 485800 429476 485852
rect 429528 485800 429534 485852
rect 429488 485772 429516 485800
rect 429562 485772 429568 485784
rect 429488 485744 429568 485772
rect 429562 485732 429568 485744
rect 429620 485732 429626 485784
rect 559098 485732 559104 485784
rect 559156 485772 559162 485784
rect 559190 485772 559196 485784
rect 559156 485744 559196 485772
rect 559156 485732 559162 485744
rect 559190 485732 559196 485744
rect 559248 485732 559254 485784
rect 269114 484372 269120 484424
rect 269172 484412 269178 484424
rect 302878 484412 302884 484424
rect 269172 484384 302884 484412
rect 269172 484372 269178 484384
rect 302878 484372 302884 484384
rect 302936 484372 302942 484424
rect 429562 482944 429568 482996
rect 429620 482984 429626 482996
rect 429654 482984 429660 482996
rect 429620 482956 429660 482984
rect 429620 482944 429626 482956
rect 429654 482944 429660 482956
rect 429712 482944 429718 482996
rect 2958 480224 2964 480276
rect 3016 480264 3022 480276
rect 20070 480264 20076 480276
rect 3016 480236 20076 480264
rect 3016 480224 3022 480236
rect 20070 480224 20076 480236
rect 20128 480224 20134 480276
rect 402238 480224 402244 480276
rect 402296 480264 402302 480276
rect 437474 480264 437480 480276
rect 402296 480236 437480 480264
rect 402296 480224 402302 480236
rect 437474 480224 437480 480236
rect 437532 480224 437538 480276
rect 302970 477504 302976 477556
rect 303028 477544 303034 477556
rect 307110 477544 307116 477556
rect 303028 477516 307116 477544
rect 303028 477504 303034 477516
rect 307110 477504 307116 477516
rect 307168 477504 307174 477556
rect 429654 476116 429660 476128
rect 429580 476088 429660 476116
rect 429580 476060 429608 476088
rect 429654 476076 429660 476088
rect 429712 476076 429718 476128
rect 559006 476076 559012 476128
rect 559064 476116 559070 476128
rect 559190 476116 559196 476128
rect 559064 476088 559196 476116
rect 559064 476076 559070 476088
rect 559190 476076 559196 476088
rect 559248 476076 559254 476128
rect 429562 476008 429568 476060
rect 429620 476008 429626 476060
rect 559098 473288 559104 473340
rect 559156 473328 559162 473340
rect 559190 473328 559196 473340
rect 559156 473300 559196 473328
rect 559156 473288 559162 473300
rect 559190 473288 559196 473300
rect 559248 473288 559254 473340
rect 299658 466420 299664 466472
rect 299716 466420 299722 466472
rect 559190 466460 559196 466472
rect 559116 466432 559196 466460
rect 299676 466392 299704 466420
rect 559116 466404 559144 466432
rect 559190 466420 559196 466432
rect 559248 466420 559254 466472
rect 299750 466392 299756 466404
rect 299676 466364 299756 466392
rect 299750 466352 299756 466364
rect 299808 466352 299814 466404
rect 559098 466352 559104 466404
rect 559156 466352 559162 466404
rect 299750 463632 299756 463684
rect 299808 463672 299814 463684
rect 299842 463672 299848 463684
rect 299808 463644 299848 463672
rect 299808 463632 299814 463644
rect 299842 463632 299848 463644
rect 299900 463632 299906 463684
rect 188890 460164 188896 460216
rect 188948 460204 188954 460216
rect 302970 460204 302976 460216
rect 188948 460176 302976 460204
rect 188948 460164 188954 460176
rect 302970 460164 302976 460176
rect 303028 460164 303034 460216
rect 59814 459484 59820 459536
rect 59872 459524 59878 459536
rect 188890 459524 188896 459536
rect 59872 459496 188896 459524
rect 59872 459484 59878 459496
rect 188890 459484 188896 459496
rect 188948 459484 188954 459536
rect 302970 459484 302976 459536
rect 303028 459524 303034 459536
rect 438118 459524 438124 459536
rect 303028 459496 438124 459524
rect 303028 459484 303034 459496
rect 438118 459484 438124 459496
rect 438176 459484 438182 459536
rect 302878 459416 302884 459468
rect 302936 459456 302942 459468
rect 389174 459456 389180 459468
rect 302936 459428 389180 459456
rect 302936 459416 302942 459428
rect 389174 459416 389180 459428
rect 389232 459416 389238 459468
rect 77294 458124 77300 458176
rect 77352 458164 77358 458176
rect 86310 458164 86316 458176
rect 77352 458136 86316 458164
rect 77352 458124 77358 458136
rect 86310 458124 86316 458136
rect 86368 458164 86374 458176
rect 86862 458164 86868 458176
rect 86368 458136 86868 458164
rect 86368 458124 86374 458136
rect 86862 458124 86868 458136
rect 86920 458124 86926 458176
rect 99374 458124 99380 458176
rect 99432 458164 99438 458176
rect 105354 458164 105360 458176
rect 99432 458136 105360 458164
rect 99432 458124 99438 458136
rect 105354 458124 105360 458136
rect 105412 458124 105418 458176
rect 122742 458124 122748 458176
rect 122800 458164 122806 458176
rect 127066 458164 127072 458176
rect 122800 458136 127072 458164
rect 122800 458124 122806 458136
rect 127066 458124 127072 458136
rect 127124 458124 127130 458176
rect 142062 458124 142068 458176
rect 142120 458164 142126 458176
rect 146938 458164 146944 458176
rect 142120 458136 146944 458164
rect 142120 458124 142126 458136
rect 146938 458124 146944 458136
rect 146996 458124 147002 458176
rect 161382 458124 161388 458176
rect 161440 458164 161446 458176
rect 190454 458164 190460 458176
rect 161440 458136 190460 458164
rect 161440 458124 161446 458136
rect 190454 458124 190460 458136
rect 190512 458124 190518 458176
rect 200022 458124 200028 458176
rect 200080 458164 200086 458176
rect 209774 458164 209780 458176
rect 200080 458136 209780 458164
rect 200080 458124 200086 458136
rect 209774 458124 209780 458136
rect 209832 458124 209838 458176
rect 215294 458124 215300 458176
rect 215352 458164 215358 458176
rect 217226 458164 217232 458176
rect 215352 458136 217232 458164
rect 215352 458124 215358 458136
rect 217226 458124 217232 458136
rect 217284 458124 217290 458176
rect 219342 458124 219348 458176
rect 219400 458164 219406 458176
rect 226334 458164 226340 458176
rect 219400 458136 226340 458164
rect 219400 458124 219406 458136
rect 226334 458124 226340 458136
rect 226392 458124 226398 458176
rect 335354 458124 335360 458176
rect 335412 458164 335418 458176
rect 344738 458164 344744 458176
rect 335412 458136 344744 458164
rect 335412 458124 335418 458136
rect 344738 458124 344744 458136
rect 344796 458164 344802 458176
rect 353294 458164 353300 458176
rect 344796 458136 353300 458164
rect 344796 458124 344802 458136
rect 353294 458124 353300 458136
rect 353352 458124 353358 458176
rect 354030 458124 354036 458176
rect 354088 458164 354094 458176
rect 484394 458164 484400 458176
rect 354088 458136 484400 458164
rect 354088 458124 354094 458136
rect 484394 458124 484400 458136
rect 484452 458124 484458 458176
rect 79962 458056 79968 458108
rect 80020 458096 80026 458108
rect 89070 458096 89076 458108
rect 80020 458068 89076 458096
rect 80020 458056 80026 458068
rect 89070 458056 89076 458068
rect 89128 458056 89134 458108
rect 91094 458056 91100 458108
rect 91152 458096 91158 458108
rect 100570 458096 100576 458108
rect 91152 458068 100576 458096
rect 91152 458056 91158 458068
rect 100570 458056 100576 458068
rect 100628 458056 100634 458108
rect 107654 458056 107660 458108
rect 107712 458096 107718 458108
rect 223574 458096 223580 458108
rect 107712 458068 223580 458096
rect 107712 458056 107718 458068
rect 223574 458056 223580 458068
rect 223632 458056 223638 458108
rect 223666 458056 223672 458108
rect 223724 458096 223730 458108
rect 231854 458096 231860 458108
rect 223724 458068 231860 458096
rect 223724 458056 223730 458068
rect 231854 458056 231860 458068
rect 231912 458056 231918 458108
rect 329098 458056 329104 458108
rect 329156 458096 329162 458108
rect 338022 458096 338028 458108
rect 329156 458068 338028 458096
rect 329156 458056 329162 458068
rect 338022 458056 338028 458068
rect 338080 458056 338086 458108
rect 344370 458056 344376 458108
rect 344428 458096 344434 458108
rect 351914 458096 351920 458108
rect 344428 458068 351920 458096
rect 344428 458056 344434 458068
rect 351914 458056 351920 458068
rect 351972 458056 351978 458108
rect 352742 458056 352748 458108
rect 352800 458096 352806 458108
rect 483014 458096 483020 458108
rect 352800 458068 483020 458096
rect 352800 458056 352806 458068
rect 483014 458056 483020 458068
rect 483072 458056 483078 458108
rect 75822 457988 75828 458040
rect 75880 458028 75886 458040
rect 84194 458028 84200 458040
rect 75880 458000 84200 458028
rect 75880 457988 75886 458000
rect 84194 457988 84200 458000
rect 84252 458028 84258 458040
rect 93578 458028 93584 458040
rect 84252 458000 93584 458028
rect 84252 457988 84258 458000
rect 93578 457988 93584 458000
rect 93636 458028 93642 458040
rect 102778 458028 102784 458040
rect 93636 458000 102784 458028
rect 93636 457988 93642 458000
rect 102778 457988 102784 458000
rect 102836 457988 102842 458040
rect 106274 457988 106280 458040
rect 106332 458028 106338 458040
rect 220814 458028 220820 458040
rect 106332 458000 220820 458028
rect 106332 457988 106338 458000
rect 220814 457988 220820 458000
rect 220872 457988 220878 458040
rect 224310 457988 224316 458040
rect 224368 458028 224374 458040
rect 233234 458028 233240 458040
rect 224368 458000 233240 458028
rect 224368 457988 224374 458000
rect 233234 457988 233240 458000
rect 233292 457988 233298 458040
rect 343542 457988 343548 458040
rect 343600 458028 343606 458040
rect 351822 458028 351828 458040
rect 343600 458000 351828 458028
rect 343600 457988 343606 458000
rect 351822 457988 351828 458000
rect 351880 457988 351886 458040
rect 353938 457988 353944 458040
rect 353996 458028 354002 458040
rect 483198 458028 483204 458040
rect 353996 458000 483204 458028
rect 353996 457988 354002 458000
rect 483198 457988 483204 458000
rect 483256 457988 483262 458040
rect 86862 457920 86868 457972
rect 86920 457960 86926 457972
rect 95786 457960 95792 457972
rect 86920 457932 95792 457960
rect 86920 457920 86926 457932
rect 95786 457920 95792 457932
rect 95844 457960 95850 457972
rect 99374 457960 99380 457972
rect 95844 457932 99380 457960
rect 95844 457920 95850 457932
rect 99374 457920 99380 457932
rect 99432 457920 99438 457972
rect 108758 457920 108764 457972
rect 108816 457960 108822 457972
rect 122742 457960 122748 457972
rect 108816 457932 122748 457960
rect 108816 457920 108822 457932
rect 122742 457920 122748 457932
rect 122800 457920 122806 457972
rect 127066 457920 127072 457972
rect 127124 457960 127130 457972
rect 142062 457960 142068 457972
rect 127124 457932 142068 457960
rect 127124 457920 127130 457932
rect 142062 457920 142068 457932
rect 142120 457920 142126 457972
rect 146938 457920 146944 457972
rect 146996 457960 147002 457972
rect 161382 457960 161388 457972
rect 146996 457932 161388 457960
rect 146996 457920 147002 457932
rect 161382 457920 161388 457932
rect 161440 457920 161446 457972
rect 190454 457920 190460 457972
rect 190512 457960 190518 457972
rect 200022 457960 200028 457972
rect 190512 457932 200028 457960
rect 190512 457920 190518 457932
rect 200022 457920 200028 457932
rect 200080 457920 200086 457972
rect 224954 457920 224960 457972
rect 225012 457960 225018 457972
rect 225874 457960 225880 457972
rect 225012 457932 225880 457960
rect 225012 457920 225018 457932
rect 225874 457920 225880 457932
rect 225932 457960 225938 457972
rect 234614 457960 234620 457972
rect 225932 457932 234620 457960
rect 225932 457920 225938 457932
rect 234614 457920 234620 457932
rect 234672 457920 234678 457972
rect 336550 457920 336556 457972
rect 336608 457960 336614 457972
rect 345934 457960 345940 457972
rect 336608 457932 345940 457960
rect 336608 457920 336614 457932
rect 345934 457920 345940 457932
rect 345992 457960 345998 457972
rect 353662 457960 353668 457972
rect 345992 457932 353668 457960
rect 345992 457920 345998 457932
rect 353662 457920 353668 457932
rect 353720 457920 353726 457972
rect 471790 457920 471796 457972
rect 471848 457960 471854 457972
rect 480438 457960 480444 457972
rect 471848 457932 480444 457960
rect 471848 457920 471854 457932
rect 480438 457920 480444 457932
rect 480496 457920 480502 457972
rect 81342 457852 81348 457904
rect 81400 457892 81406 457904
rect 90174 457892 90180 457904
rect 81400 457864 90180 457892
rect 81400 457852 81406 457864
rect 90174 457852 90180 457864
rect 90232 457892 90238 457904
rect 99466 457892 99472 457904
rect 90232 457864 99472 457892
rect 90232 457852 90238 457864
rect 99466 457852 99472 457864
rect 99524 457892 99530 457904
rect 108776 457892 108804 457920
rect 99524 457864 108804 457892
rect 99524 457852 99530 457864
rect 208210 457852 208216 457904
rect 208268 457892 208274 457904
rect 216674 457892 216680 457904
rect 208268 457864 216680 457892
rect 208268 457852 208274 457864
rect 216674 457852 216680 457864
rect 216732 457892 216738 457904
rect 217134 457892 217140 457904
rect 216732 457864 217140 457892
rect 216732 457852 216738 457864
rect 217134 457852 217140 457864
rect 217192 457852 217198 457904
rect 217226 457852 217232 457904
rect 217284 457892 217290 457904
rect 224310 457892 224316 457904
rect 217284 457864 224316 457892
rect 217284 457852 217290 457864
rect 224310 457852 224316 457864
rect 224368 457852 224374 457904
rect 331306 457852 331312 457904
rect 331364 457892 331370 457904
rect 331858 457892 331864 457904
rect 331364 457864 331864 457892
rect 331364 457852 331370 457864
rect 331858 457852 331864 457864
rect 331916 457892 331922 457904
rect 341242 457892 341248 457904
rect 331916 457864 341248 457892
rect 331916 457852 331922 457864
rect 341242 457852 341248 457864
rect 341300 457892 341306 457904
rect 350534 457892 350540 457904
rect 341300 457864 350540 457892
rect 341300 457852 341306 457864
rect 350534 457852 350540 457864
rect 350592 457852 350598 457904
rect 350626 457852 350632 457904
rect 350684 457892 350690 457904
rect 356054 457892 356060 457904
rect 350684 457864 356060 457892
rect 350684 457852 350690 457864
rect 356054 457852 356060 457864
rect 356112 457852 356118 457904
rect 460198 457852 460204 457904
rect 460256 457892 460262 457904
rect 468754 457892 468760 457904
rect 460256 457864 468760 457892
rect 460256 457852 460262 457864
rect 468754 457852 468760 457864
rect 468812 457892 468818 457904
rect 478322 457892 478328 457904
rect 468812 457864 478328 457892
rect 468812 457852 468818 457864
rect 478322 457852 478328 457864
rect 478380 457892 478386 457904
rect 487154 457892 487160 457904
rect 478380 457864 487160 457892
rect 478380 457852 478386 457864
rect 487154 457852 487160 457864
rect 487212 457852 487218 457904
rect 78582 457784 78588 457836
rect 78640 457824 78646 457836
rect 87874 457824 87880 457836
rect 78640 457796 87880 457824
rect 78640 457784 78646 457796
rect 87874 457784 87880 457796
rect 87932 457824 87938 457836
rect 97166 457824 97172 457836
rect 87932 457796 97172 457824
rect 87932 457784 87938 457796
rect 97166 457784 97172 457796
rect 97224 457824 97230 457836
rect 97902 457824 97908 457836
rect 97224 457796 97908 457824
rect 97224 457784 97230 457796
rect 97902 457784 97908 457796
rect 97960 457784 97966 457836
rect 213086 457784 213092 457836
rect 213144 457824 213150 457836
rect 222562 457824 222568 457836
rect 213144 457796 222568 457824
rect 213144 457784 213150 457796
rect 222562 457784 222568 457796
rect 222620 457824 222626 457836
rect 231854 457824 231860 457836
rect 222620 457796 231860 457824
rect 222620 457784 222626 457796
rect 231854 457784 231860 457796
rect 231912 457784 231918 457836
rect 339034 457784 339040 457836
rect 339092 457824 339098 457836
rect 340874 457824 340880 457836
rect 339092 457796 340880 457824
rect 339092 457784 339098 457796
rect 340874 457784 340880 457796
rect 340932 457784 340938 457836
rect 464982 457784 464988 457836
rect 465040 457824 465046 457836
rect 465040 457796 471468 457824
rect 465040 457784 465046 457796
rect 89070 457716 89076 457768
rect 89128 457756 89134 457768
rect 98546 457756 98552 457768
rect 89128 457728 98552 457756
rect 89128 457716 89134 457728
rect 98546 457716 98552 457728
rect 98604 457756 98610 457768
rect 107654 457756 107660 457768
rect 98604 457728 107660 457756
rect 98604 457716 98610 457728
rect 107654 457716 107660 457728
rect 107712 457716 107718 457768
rect 214006 457716 214012 457768
rect 214064 457756 214070 457768
rect 223666 457756 223672 457768
rect 214064 457728 223672 457756
rect 214064 457716 214070 457728
rect 223666 457716 223672 457728
rect 223724 457716 223730 457768
rect 226426 457716 226432 457768
rect 226484 457756 226490 457768
rect 227162 457756 227168 457768
rect 226484 457728 227168 457756
rect 226484 457716 226490 457728
rect 227162 457716 227168 457728
rect 227220 457756 227226 457768
rect 235994 457756 236000 457768
rect 227220 457728 236000 457756
rect 227220 457716 227226 457728
rect 235994 457716 236000 457728
rect 236052 457716 236058 457768
rect 332594 457716 332600 457768
rect 332652 457756 332658 457768
rect 333146 457756 333152 457768
rect 332652 457728 333152 457756
rect 332652 457716 332658 457728
rect 333146 457716 333152 457728
rect 333204 457756 333210 457768
rect 342530 457756 342536 457768
rect 333204 457728 342536 457756
rect 333204 457716 333210 457728
rect 342530 457716 342536 457728
rect 342588 457756 342594 457768
rect 343542 457756 343548 457768
rect 342588 457728 343548 457756
rect 342588 457716 342594 457728
rect 343542 457716 343548 457728
rect 343600 457716 343606 457768
rect 349246 457716 349252 457768
rect 349304 457756 349310 457768
rect 349304 457728 349660 457756
rect 349304 457716 349310 457728
rect 73062 457648 73068 457700
rect 73120 457688 73126 457700
rect 81894 457688 81900 457700
rect 73120 457660 81900 457688
rect 73120 457648 73126 457660
rect 81894 457648 81900 457660
rect 81952 457688 81958 457700
rect 91094 457688 91100 457700
rect 81952 457660 91100 457688
rect 81952 457648 81958 457660
rect 91094 457648 91100 457660
rect 91152 457648 91158 457700
rect 97902 457648 97908 457700
rect 97960 457688 97966 457700
rect 106274 457688 106280 457700
rect 97960 457660 106280 457688
rect 97960 457648 97966 457660
rect 106274 457648 106280 457660
rect 106332 457648 106338 457700
rect 176562 457648 176568 457700
rect 176620 457688 176626 457700
rect 201494 457688 201500 457700
rect 176620 457660 201500 457688
rect 176620 457648 176626 457660
rect 201494 457648 201500 457660
rect 201552 457648 201558 457700
rect 207750 457648 207756 457700
rect 207808 457688 207814 457700
rect 209682 457688 209688 457700
rect 207808 457660 209688 457688
rect 207808 457648 207814 457660
rect 209682 457648 209688 457660
rect 209740 457688 209746 457700
rect 218882 457688 218888 457700
rect 209740 457660 218888 457688
rect 209740 457648 209746 457660
rect 218882 457648 218888 457660
rect 218940 457688 218946 457700
rect 228358 457688 228364 457700
rect 218940 457660 228364 457688
rect 218940 457648 218946 457660
rect 228358 457648 228364 457660
rect 228416 457688 228422 457700
rect 237374 457688 237380 457700
rect 228416 457660 237380 457688
rect 228416 457648 228422 457660
rect 237374 457648 237380 457660
rect 237432 457648 237438 457700
rect 338022 457648 338028 457700
rect 338080 457688 338086 457700
rect 346854 457688 346860 457700
rect 338080 457660 346860 457688
rect 338080 457648 338086 457660
rect 346854 457648 346860 457660
rect 346912 457688 346918 457700
rect 349632 457688 349660 457728
rect 349706 457716 349712 457768
rect 349764 457756 349770 457768
rect 349764 457728 353616 457756
rect 349764 457716 349770 457728
rect 353588 457688 353616 457728
rect 453482 457716 453488 457768
rect 453540 457756 453546 457768
rect 463050 457756 463056 457768
rect 453540 457728 463056 457756
rect 453540 457716 453546 457728
rect 463050 457716 463056 457728
rect 463108 457756 463114 457768
rect 471330 457756 471336 457768
rect 463108 457728 471336 457756
rect 463108 457716 463114 457728
rect 471330 457716 471336 457728
rect 471388 457716 471394 457768
rect 471440 457756 471468 457796
rect 471514 457784 471520 457836
rect 471572 457824 471578 457836
rect 475470 457824 475476 457836
rect 471572 457796 475476 457824
rect 471572 457784 471578 457796
rect 475470 457784 475476 457796
rect 475528 457824 475534 457836
rect 484394 457824 484400 457836
rect 475528 457796 484400 457824
rect 475528 457784 475534 457796
rect 484394 457784 484400 457796
rect 484452 457784 484458 457836
rect 473446 457756 473452 457768
rect 471440 457728 473452 457756
rect 473446 457716 473452 457728
rect 473504 457756 473510 457768
rect 480254 457756 480260 457768
rect 473504 457728 480260 457756
rect 473504 457716 473510 457728
rect 480254 457716 480260 457728
rect 480312 457716 480318 457768
rect 357434 457688 357440 457700
rect 346912 457660 349384 457688
rect 349632 457660 353524 457688
rect 353588 457660 357440 457688
rect 346912 457648 346918 457660
rect 74166 457580 74172 457632
rect 74224 457620 74230 457632
rect 82814 457620 82820 457632
rect 74224 457592 82820 457620
rect 74224 457580 74230 457592
rect 82814 457580 82820 457592
rect 82872 457620 82878 457632
rect 92474 457620 92480 457632
rect 82872 457592 92480 457620
rect 82872 457580 82878 457592
rect 92474 457580 92480 457592
rect 92532 457620 92538 457632
rect 101858 457620 101864 457632
rect 92532 457592 101864 457620
rect 92532 457580 92538 457592
rect 101858 457580 101864 457592
rect 101916 457580 101922 457632
rect 175182 457580 175188 457632
rect 175240 457620 175246 457632
rect 200206 457620 200212 457632
rect 175240 457592 200212 457620
rect 175240 457580 175246 457592
rect 200206 457580 200212 457592
rect 200264 457580 200270 457632
rect 209130 457580 209136 457632
rect 209188 457620 209194 457632
rect 210510 457620 210516 457632
rect 209188 457592 210516 457620
rect 209188 457580 209194 457592
rect 210510 457580 210516 457592
rect 210568 457620 210574 457632
rect 220170 457620 220176 457632
rect 210568 457592 220176 457620
rect 210568 457580 210574 457592
rect 220170 457580 220176 457592
rect 220228 457620 220234 457632
rect 229554 457620 229560 457632
rect 220228 457592 229560 457620
rect 220228 457580 220234 457592
rect 229554 457580 229560 457592
rect 229612 457620 229618 457632
rect 238754 457620 238760 457632
rect 229612 457592 238760 457620
rect 229612 457580 229618 457592
rect 238754 457580 238760 457592
rect 238812 457580 238818 457632
rect 339862 457580 339868 457632
rect 339920 457620 339926 457632
rect 349246 457620 349252 457632
rect 339920 457592 349252 457620
rect 339920 457580 339926 457592
rect 349246 457580 349252 457592
rect 349304 457580 349310 457632
rect 349356 457620 349384 457660
rect 350626 457620 350632 457632
rect 349356 457592 350632 457620
rect 350626 457580 350632 457592
rect 350684 457580 350690 457632
rect 353496 457620 353524 457660
rect 357434 457648 357440 457660
rect 357492 457648 357498 457700
rect 359458 457648 359464 457700
rect 359516 457688 359522 457700
rect 458174 457688 458180 457700
rect 359516 457660 458180 457688
rect 359516 457648 359522 457660
rect 458174 457648 458180 457660
rect 458232 457648 458238 457700
rect 460382 457648 460388 457700
rect 460440 457688 460446 457700
rect 469950 457688 469956 457700
rect 460440 457660 469956 457688
rect 460440 457648 460446 457660
rect 469950 457648 469956 457660
rect 470008 457688 470014 457700
rect 479426 457688 479432 457700
rect 470008 457660 479432 457688
rect 470008 457648 470014 457660
rect 479426 457648 479432 457660
rect 479484 457688 479490 457700
rect 488534 457688 488540 457700
rect 479484 457660 488540 457688
rect 479484 457648 479490 457660
rect 488534 457648 488540 457660
rect 488592 457648 488598 457700
rect 358814 457620 358820 457632
rect 353496 457592 358820 457620
rect 358814 457580 358820 457592
rect 358872 457580 358878 457632
rect 453298 457580 453304 457632
rect 453356 457620 453362 457632
rect 461762 457620 461768 457632
rect 453356 457592 461768 457620
rect 453356 457580 453362 457592
rect 461762 457580 461768 457592
rect 461820 457620 461826 457632
rect 471790 457620 471796 457632
rect 461820 457592 471796 457620
rect 461820 457580 461826 457592
rect 471790 457580 471796 457592
rect 471848 457580 471854 457632
rect 472250 457620 472256 457632
rect 471900 457592 472256 457620
rect 77202 457512 77208 457564
rect 77260 457552 77266 457564
rect 85482 457552 85488 457564
rect 77260 457524 85488 457552
rect 77260 457512 77266 457524
rect 85482 457512 85488 457524
rect 85540 457552 85546 457564
rect 94774 457552 94780 457564
rect 85540 457524 94780 457552
rect 85540 457512 85546 457524
rect 94774 457512 94780 457524
rect 94832 457552 94838 457564
rect 104250 457552 104256 457564
rect 94832 457524 104256 457552
rect 94832 457512 94838 457524
rect 104250 457512 104256 457524
rect 104308 457512 104314 457564
rect 172422 457512 172428 457564
rect 172480 457552 172486 457564
rect 198734 457552 198740 457564
rect 172480 457524 198740 457552
rect 172480 457512 172486 457524
rect 198734 457512 198740 457524
rect 198792 457512 198798 457564
rect 212442 457512 212448 457564
rect 212500 457552 212506 457564
rect 221366 457552 221372 457564
rect 212500 457524 221372 457552
rect 212500 457512 212506 457524
rect 221366 457512 221372 457524
rect 221424 457552 221430 457564
rect 230474 457552 230480 457564
rect 221424 457524 230480 457552
rect 221424 457512 221430 457524
rect 230474 457512 230480 457524
rect 230532 457512 230538 457564
rect 334066 457512 334072 457564
rect 334124 457552 334130 457564
rect 344370 457552 344376 457564
rect 334124 457524 344376 457552
rect 334124 457512 334130 457524
rect 344370 457512 344376 457524
rect 344428 457512 344434 457564
rect 353662 457512 353668 457564
rect 353720 457552 353726 457564
rect 355042 457552 355048 457564
rect 353720 457524 355048 457552
rect 353720 457512 353726 457524
rect 355042 457512 355048 457524
rect 355100 457512 355106 457564
rect 358078 457512 358084 457564
rect 358136 457552 358142 457564
rect 456794 457552 456800 457564
rect 358136 457524 456800 457552
rect 358136 457512 358142 457524
rect 456794 457512 456800 457524
rect 456852 457512 456858 457564
rect 465166 457512 465172 457564
rect 465224 457552 465230 457564
rect 471238 457552 471244 457564
rect 465224 457524 471244 457552
rect 465224 457512 465230 457524
rect 471238 457512 471244 457524
rect 471296 457512 471302 457564
rect 471330 457512 471336 457564
rect 471388 457552 471394 457564
rect 471900 457552 471928 457592
rect 472250 457580 472256 457592
rect 472308 457620 472314 457632
rect 481634 457620 481640 457632
rect 472308 457592 481640 457620
rect 472308 457580 472314 457592
rect 481634 457580 481640 457592
rect 481692 457580 481698 457632
rect 471388 457524 471928 457552
rect 471388 457512 471394 457524
rect 476298 457512 476304 457564
rect 476356 457552 476362 457564
rect 476942 457552 476948 457564
rect 476356 457524 476948 457552
rect 476356 457512 476362 457524
rect 476942 457512 476948 457524
rect 477000 457552 477006 457564
rect 485774 457552 485780 457564
rect 477000 457524 485780 457552
rect 477000 457512 477006 457524
rect 485774 457512 485780 457524
rect 485832 457512 485838 457564
rect 60734 457444 60740 457496
rect 60792 457484 60798 457496
rect 63678 457484 63684 457496
rect 60792 457456 63684 457484
rect 60792 457444 60798 457456
rect 63678 457444 63684 457456
rect 63736 457484 63742 457496
rect 193858 457484 193864 457496
rect 63736 457456 193864 457484
rect 63736 457444 63742 457456
rect 193858 457444 193864 457456
rect 193916 457484 193922 457496
rect 313734 457484 313740 457496
rect 193916 457456 313740 457484
rect 193916 457444 193922 457456
rect 313734 457444 313740 457456
rect 313792 457484 313798 457496
rect 442994 457484 443000 457496
rect 313792 457456 443000 457484
rect 313792 457444 313798 457456
rect 442994 457444 443000 457456
rect 443052 457444 443058 457496
rect 443638 457444 443644 457496
rect 443696 457484 443702 457496
rect 459554 457484 459560 457496
rect 443696 457456 459560 457484
rect 443696 457444 443702 457456
rect 459554 457444 459560 457456
rect 459612 457444 459618 457496
rect 465718 457444 465724 457496
rect 465776 457484 465782 457496
rect 487154 457484 487160 457496
rect 465776 457456 487160 457484
rect 465776 457444 465782 457456
rect 487154 457444 487160 457456
rect 487212 457444 487218 457496
rect 171042 457376 171048 457428
rect 171100 457416 171106 457428
rect 197354 457416 197360 457428
rect 171100 457388 197360 457416
rect 171100 457376 171106 457388
rect 197354 457376 197360 457388
rect 197412 457376 197418 457428
rect 209038 457376 209044 457428
rect 209096 457416 209102 457428
rect 209096 457388 215708 457416
rect 209096 457376 209102 457388
rect 133782 457308 133788 457360
rect 133840 457348 133846 457360
rect 195974 457348 195980 457360
rect 133840 457320 195980 457348
rect 133840 457308 133846 457320
rect 195974 457308 195980 457320
rect 196032 457308 196038 457360
rect 202138 457308 202144 457360
rect 202196 457348 202202 457360
rect 212442 457348 212448 457360
rect 202196 457320 212448 457348
rect 202196 457308 202202 457320
rect 212442 457308 212448 457320
rect 212500 457308 212506 457360
rect 215680 457348 215708 457388
rect 217134 457376 217140 457428
rect 217192 457416 217198 457428
rect 224954 457416 224960 457428
rect 217192 457388 224960 457416
rect 217192 457376 217198 457388
rect 224954 457376 224960 457388
rect 225012 457376 225018 457428
rect 309778 457376 309784 457428
rect 309836 457416 309842 457428
rect 331214 457416 331220 457428
rect 309836 457388 331220 457416
rect 309836 457376 309842 457388
rect 331214 457376 331220 457388
rect 331272 457376 331278 457428
rect 340874 457376 340880 457428
rect 340932 457416 340938 457428
rect 348234 457416 348240 457428
rect 340932 457388 348240 457416
rect 340932 457376 340938 457388
rect 348234 457376 348240 457388
rect 348292 457416 348298 457428
rect 349706 457416 349712 457428
rect 348292 457388 349712 457416
rect 348292 457376 348298 457388
rect 349706 457376 349712 457388
rect 349764 457376 349770 457428
rect 355318 457376 355324 457428
rect 355376 457416 355382 457428
rect 454034 457416 454040 457428
rect 355376 457388 454040 457416
rect 355376 457376 355382 457388
rect 454034 457376 454040 457388
rect 454092 457376 454098 457428
rect 454678 457376 454684 457428
rect 454736 457416 454742 457428
rect 464982 457416 464988 457428
rect 454736 457388 464988 457416
rect 454736 457376 454742 457388
rect 464982 457376 464988 457388
rect 465040 457376 465046 457428
rect 467098 457376 467104 457428
rect 467156 457416 467162 457428
rect 488534 457416 488540 457428
rect 467156 457388 488540 457416
rect 467156 457376 467162 457388
rect 488534 457376 488540 457388
rect 488592 457376 488598 457428
rect 217594 457348 217600 457360
rect 215680 457320 217600 457348
rect 217594 457308 217600 457320
rect 217652 457348 217658 457360
rect 226426 457348 226432 457360
rect 217652 457320 226432 457348
rect 217652 457308 217658 457320
rect 226426 457308 226432 457320
rect 226484 457308 226490 457360
rect 322198 457308 322204 457360
rect 322256 457348 322262 457360
rect 331306 457348 331312 457360
rect 322256 457320 331312 457348
rect 322256 457308 322262 457320
rect 331306 457308 331312 457320
rect 331364 457308 331370 457360
rect 342898 457308 342904 457360
rect 342956 457348 342962 457360
rect 452654 457348 452660 457360
rect 342956 457320 452660 457348
rect 342956 457308 342962 457320
rect 452654 457308 452660 457320
rect 452712 457308 452718 457360
rect 464338 457308 464344 457360
rect 464396 457348 464402 457360
rect 485774 457348 485780 457360
rect 464396 457320 485780 457348
rect 464396 457308 464402 457320
rect 485774 457308 485780 457320
rect 485832 457308 485838 457360
rect 100570 457240 100576 457292
rect 100628 457280 100634 457292
rect 209774 457280 209780 457292
rect 100628 457252 209780 457280
rect 100628 457240 100634 457252
rect 209774 457240 209780 457252
rect 209832 457240 209838 457292
rect 209866 457240 209872 457292
rect 209924 457280 209930 457292
rect 219342 457280 219348 457292
rect 209924 457252 219348 457280
rect 209924 457240 209930 457252
rect 219342 457240 219348 457252
rect 219400 457240 219406 457292
rect 312538 457240 312544 457292
rect 312596 457280 312602 457292
rect 329834 457280 329840 457292
rect 312596 457252 329840 457280
rect 312596 457240 312602 457252
rect 329834 457240 329840 457252
rect 329892 457240 329898 457292
rect 349798 457240 349804 457292
rect 349856 457280 349862 457292
rect 477494 457280 477500 457292
rect 349856 457252 477500 457280
rect 349856 457240 349862 457252
rect 477494 457240 477500 457252
rect 477552 457240 477558 457292
rect 480254 457240 480260 457292
rect 480312 457280 480318 457292
rect 483106 457280 483112 457292
rect 480312 457252 483112 457280
rect 480312 457240 480318 457252
rect 483106 457240 483112 457252
rect 483164 457240 483170 457292
rect 101858 457172 101864 457224
rect 101916 457212 101922 457224
rect 212534 457212 212540 457224
rect 101916 457184 212540 457212
rect 101916 457172 101922 457184
rect 212534 457172 212540 457184
rect 212592 457172 212598 457224
rect 327902 457172 327908 457224
rect 327960 457212 327966 457224
rect 336550 457212 336556 457224
rect 327960 457184 336556 457212
rect 327960 457172 327966 457184
rect 336550 457172 336556 457184
rect 336608 457172 336614 457224
rect 351178 457172 351184 457224
rect 351236 457212 351242 457224
rect 478874 457212 478880 457224
rect 351236 457184 478880 457212
rect 351236 457172 351242 457184
rect 478874 457172 478880 457184
rect 478932 457172 478938 457224
rect 63402 457104 63408 457156
rect 63460 457144 63466 457156
rect 73154 457144 73160 457156
rect 63460 457116 73160 457144
rect 63460 457104 63466 457116
rect 73154 457104 73160 457116
rect 73212 457104 73218 457156
rect 102778 457104 102784 457156
rect 102836 457144 102842 457156
rect 213914 457144 213920 457156
rect 102836 457116 213920 457144
rect 102836 457104 102842 457116
rect 213914 457104 213920 457116
rect 213972 457104 213978 457156
rect 215202 457104 215208 457156
rect 215260 457144 215266 457156
rect 246298 457144 246304 457156
rect 215260 457116 246304 457144
rect 215260 457104 215266 457116
rect 246298 457104 246304 457116
rect 246356 457104 246362 457156
rect 315298 457104 315304 457156
rect 315356 457144 315362 457156
rect 328454 457144 328460 457156
rect 315356 457116 328460 457144
rect 315356 457104 315362 457116
rect 328454 457104 328460 457116
rect 328512 457104 328518 457156
rect 329282 457104 329288 457156
rect 329340 457144 329346 457156
rect 339034 457144 339040 457156
rect 329340 457116 339040 457144
rect 329340 457104 329346 457116
rect 339034 457104 339040 457116
rect 339092 457104 339098 457156
rect 352558 457104 352564 457156
rect 352616 457144 352622 457156
rect 480530 457144 480536 457156
rect 352616 457116 480536 457144
rect 352616 457104 352622 457116
rect 480530 457104 480536 457116
rect 480588 457104 480594 457156
rect 70302 457036 70308 457088
rect 70360 457076 70366 457088
rect 77294 457076 77300 457088
rect 70360 457048 77300 457076
rect 70360 457036 70366 457048
rect 77294 457036 77300 457048
rect 77352 457036 77358 457088
rect 104250 457036 104256 457088
rect 104308 457076 104314 457088
rect 216674 457076 216680 457088
rect 104308 457048 216680 457076
rect 104308 457036 104314 457048
rect 216674 457036 216680 457048
rect 216732 457036 216738 457088
rect 323578 457036 323584 457088
rect 323636 457076 323642 457088
rect 332594 457076 332600 457088
rect 323636 457048 332600 457076
rect 323636 457036 323642 457048
rect 332594 457036 332600 457048
rect 332652 457036 332658 457088
rect 352650 457036 352656 457088
rect 352708 457076 352714 457088
rect 481634 457076 481640 457088
rect 352708 457048 481640 457076
rect 352708 457036 352714 457048
rect 481634 457036 481640 457048
rect 481692 457036 481698 457088
rect 68922 456968 68928 457020
rect 68980 457008 68986 457020
rect 75914 457008 75920 457020
rect 68980 456980 75920 457008
rect 68980 456968 68986 456980
rect 75914 456968 75920 456980
rect 75972 456968 75978 457020
rect 105354 456968 105360 457020
rect 105412 457008 105418 457020
rect 219434 457008 219440 457020
rect 105412 456980 219440 457008
rect 105412 456968 105418 456980
rect 219434 456968 219440 456980
rect 219492 456968 219498 457020
rect 308398 456968 308404 457020
rect 308456 457008 308462 457020
rect 317414 457008 317420 457020
rect 308456 456980 317420 457008
rect 308456 456968 308462 456980
rect 317414 456968 317420 456980
rect 317472 456968 317478 457020
rect 347038 456968 347044 457020
rect 347096 457008 347102 457020
rect 476114 457008 476120 457020
rect 347096 456980 476120 457008
rect 347096 456968 347102 456980
rect 476114 456968 476120 456980
rect 476172 456968 476178 457020
rect 66162 456900 66168 456952
rect 66220 456940 66226 456952
rect 74718 456940 74724 456952
rect 66220 456912 74724 456940
rect 66220 456900 66226 456912
rect 74718 456900 74724 456912
rect 74776 456900 74782 456952
rect 206830 456900 206836 456952
rect 206888 456940 206894 456952
rect 215294 456940 215300 456952
rect 206888 456912 215300 456940
rect 206888 456900 206894 456912
rect 215294 456900 215300 456912
rect 215352 456900 215358 456952
rect 324958 456900 324964 456952
rect 325016 456940 325022 456952
rect 334066 456940 334072 456952
rect 325016 456912 334072 456940
rect 325016 456900 325022 456912
rect 334066 456900 334072 456912
rect 334124 456900 334130 456952
rect 459370 456900 459376 456952
rect 459428 456940 459434 456952
rect 468018 456940 468024 456952
rect 459428 456912 468024 456940
rect 459428 456900 459434 456912
rect 468018 456900 468024 456912
rect 468076 456940 468082 456952
rect 476298 456940 476304 456952
rect 468076 456912 476304 456940
rect 468076 456900 468082 456912
rect 476298 456900 476304 456912
rect 476356 456900 476362 456952
rect 73062 456832 73068 456884
rect 73120 456872 73126 456884
rect 78766 456872 78772 456884
rect 73120 456844 78772 456872
rect 73120 456832 73126 456844
rect 78766 456832 78772 456844
rect 78824 456832 78830 456884
rect 205450 456832 205456 456884
rect 205508 456872 205514 456884
rect 214006 456872 214012 456884
rect 205508 456844 214012 456872
rect 205508 456832 205514 456844
rect 214006 456832 214012 456844
rect 214064 456832 214070 456884
rect 216582 456832 216588 456884
rect 216640 456872 216646 456884
rect 244918 456872 244924 456884
rect 216640 456844 244924 456872
rect 216640 456832 216646 456844
rect 244918 456832 244924 456844
rect 244976 456832 244982 456884
rect 326338 456832 326344 456884
rect 326396 456872 326402 456884
rect 335446 456872 335452 456884
rect 326396 456844 335452 456872
rect 326396 456832 326402 456844
rect 335446 456832 335452 456844
rect 335504 456832 335510 456884
rect 356698 456832 356704 456884
rect 356756 456872 356762 456884
rect 455414 456872 455420 456884
rect 356756 456844 455420 456872
rect 356756 456832 356762 456844
rect 455414 456832 455420 456844
rect 455472 456832 455478 456884
rect 456702 456832 456708 456884
rect 456760 456872 456766 456884
rect 465166 456872 465172 456884
rect 456760 456844 465172 456872
rect 456760 456832 456766 456844
rect 465166 456832 465172 456844
rect 465224 456832 465230 456884
rect 466638 456872 466644 456884
rect 466012 456844 466644 456872
rect 62022 456764 62028 456816
rect 62080 456804 62086 456816
rect 71774 456804 71780 456816
rect 62080 456776 71780 456804
rect 62080 456764 62086 456776
rect 71774 456764 71780 456776
rect 71832 456764 71838 456816
rect 76558 456764 76564 456816
rect 76616 456804 76622 456816
rect 78674 456804 78680 456816
rect 76616 456776 78680 456804
rect 76616 456764 76622 456776
rect 78674 456764 78680 456776
rect 78732 456764 78738 456816
rect 203518 456764 203524 456816
rect 203576 456804 203582 456816
rect 213086 456804 213092 456816
rect 203576 456776 213092 456804
rect 203576 456764 203582 456776
rect 213086 456764 213092 456776
rect 213144 456764 213150 456816
rect 217962 456764 217968 456816
rect 218020 456804 218026 456816
rect 242158 456804 242164 456816
rect 218020 456776 242164 456804
rect 218020 456764 218026 456776
rect 242158 456764 242164 456776
rect 242216 456764 242222 456816
rect 299842 456804 299848 456816
rect 299768 456776 299848 456804
rect 299768 456748 299796 456776
rect 299842 456764 299848 456776
rect 299900 456764 299906 456816
rect 316678 456764 316684 456816
rect 316736 456804 316742 456816
rect 324314 456804 324320 456816
rect 316736 456776 324320 456804
rect 316736 456764 316742 456776
rect 324314 456764 324320 456776
rect 324372 456764 324378 456816
rect 330478 456764 330484 456816
rect 330536 456804 330542 456816
rect 339862 456804 339868 456816
rect 330536 456776 339868 456804
rect 330536 456764 330542 456776
rect 339862 456764 339868 456776
rect 339920 456764 339926 456816
rect 458082 456764 458088 456816
rect 458140 456804 458146 456816
rect 466012 456804 466040 456844
rect 466638 456832 466644 456844
rect 466696 456872 466702 456884
rect 471146 456872 471152 456884
rect 466696 456844 471152 456872
rect 466696 456832 466702 456844
rect 471146 456832 471152 456844
rect 471204 456832 471210 456884
rect 471238 456832 471244 456884
rect 471296 456872 471302 456884
rect 474826 456872 474832 456884
rect 471296 456844 474832 456872
rect 471296 456832 471302 456844
rect 474826 456832 474832 456844
rect 474884 456872 474890 456884
rect 483014 456872 483020 456884
rect 474884 456844 483020 456872
rect 474884 456832 474890 456844
rect 483014 456832 483020 456844
rect 483072 456832 483078 456884
rect 458140 456776 466040 456804
rect 458140 456764 458146 456776
rect 559006 456764 559012 456816
rect 559064 456804 559070 456816
rect 559190 456804 559196 456816
rect 559064 456776 559196 456804
rect 559064 456764 559070 456776
rect 559190 456764 559196 456776
rect 559248 456764 559254 456816
rect 299750 456696 299756 456748
rect 299808 456696 299814 456748
rect 57606 451256 57612 451308
rect 57664 451296 57670 451308
rect 580166 451296 580172 451308
rect 57664 451268 580172 451296
rect 57664 451256 57670 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 429470 447176 429476 447228
rect 429528 447176 429534 447228
rect 559190 447176 559196 447228
rect 559248 447176 559254 447228
rect 429488 447092 429516 447176
rect 559208 447092 559236 447176
rect 429470 447040 429476 447092
rect 429528 447040 429534 447092
rect 559190 447040 559196 447092
rect 559248 447040 559254 447092
rect 299658 444388 299664 444440
rect 299716 444428 299722 444440
rect 299842 444428 299848 444440
rect 299716 444400 299848 444428
rect 299716 444388 299722 444400
rect 299842 444388 299848 444400
rect 299900 444388 299906 444440
rect 327626 444388 327632 444440
rect 327684 444428 327690 444440
rect 327718 444428 327724 444440
rect 327684 444400 327724 444428
rect 327684 444388 327690 444400
rect 327718 444388 327724 444400
rect 327776 444388 327782 444440
rect 429378 444388 429384 444440
rect 429436 444428 429442 444440
rect 429470 444428 429476 444440
rect 429436 444400 429476 444428
rect 429436 444388 429442 444400
rect 429470 444388 429476 444400
rect 429528 444388 429534 444440
rect 559098 444388 559104 444440
rect 559156 444428 559162 444440
rect 559190 444428 559196 444440
rect 559156 444400 559196 444428
rect 559156 444388 559162 444400
rect 559190 444388 559196 444400
rect 559248 444388 559254 444440
rect 242342 443232 242348 443284
rect 242400 443272 242406 443284
rect 245102 443272 245108 443284
rect 242400 443244 245108 443272
rect 242400 443232 242406 443244
rect 245102 443232 245108 443244
rect 245160 443232 245166 443284
rect 61102 442892 61108 442944
rect 61160 442932 61166 442944
rect 62022 442932 62028 442944
rect 61160 442904 62028 442932
rect 61160 442892 61166 442904
rect 62022 442892 62028 442904
rect 62080 442892 62086 442944
rect 67818 442892 67824 442944
rect 67876 442932 67882 442944
rect 68922 442932 68928 442944
rect 67876 442904 68928 442932
rect 67876 442892 67882 442904
rect 68922 442892 68928 442904
rect 68980 442892 68986 442944
rect 74626 442892 74632 442944
rect 74684 442932 74690 442944
rect 76558 442932 76564 442944
rect 74684 442904 76564 442932
rect 74684 442892 74690 442904
rect 76558 442892 76564 442904
rect 76616 442892 76622 442944
rect 76926 442892 76932 442944
rect 76984 442932 76990 442944
rect 80054 442932 80060 442944
rect 76984 442904 80060 442932
rect 76984 442892 76990 442904
rect 80054 442892 80060 442904
rect 80112 442892 80118 442944
rect 81434 442892 81440 442944
rect 81492 442932 81498 442944
rect 82814 442932 82820 442944
rect 81492 442904 82820 442932
rect 81492 442892 81498 442904
rect 82814 442892 82820 442904
rect 82872 442892 82878 442944
rect 86862 442892 86868 442944
rect 86920 442932 86926 442944
rect 87966 442932 87972 442944
rect 86920 442904 87972 442932
rect 86920 442892 86926 442904
rect 87966 442892 87972 442904
rect 88024 442892 88030 442944
rect 88242 442892 88248 442944
rect 88300 442932 88306 442944
rect 90450 442932 90456 442944
rect 88300 442904 90456 442932
rect 88300 442892 88306 442904
rect 90450 442892 90456 442904
rect 90508 442892 90514 442944
rect 92382 442892 92388 442944
rect 92440 442932 92446 442944
rect 97258 442932 97264 442944
rect 92440 442904 97264 442932
rect 92440 442892 92446 442904
rect 97258 442892 97264 442904
rect 97316 442892 97322 442944
rect 97902 442892 97908 442944
rect 97960 442932 97966 442944
rect 108574 442932 108580 442944
rect 97960 442904 108580 442932
rect 97960 442892 97966 442904
rect 108574 442892 108580 442904
rect 108632 442892 108638 442944
rect 110322 442892 110328 442944
rect 110380 442932 110386 442944
rect 131298 442932 131304 442944
rect 110380 442904 131304 442932
rect 110380 442892 110386 442904
rect 131298 442892 131304 442904
rect 131356 442892 131362 442944
rect 138014 442892 138020 442944
rect 138072 442932 138078 442944
rect 139302 442932 139308 442944
rect 138072 442904 139308 442932
rect 138072 442892 138078 442904
rect 139302 442892 139308 442904
rect 139360 442892 139366 442944
rect 139394 442892 139400 442944
rect 139452 442932 139458 442944
rect 188338 442932 188344 442944
rect 139452 442904 188344 442932
rect 139452 442892 139458 442904
rect 188338 442892 188344 442904
rect 188396 442892 188402 442944
rect 206002 442892 206008 442944
rect 206060 442932 206066 442944
rect 207750 442932 207756 442944
rect 206060 442904 207756 442932
rect 206060 442892 206066 442904
rect 207750 442892 207756 442904
rect 207808 442892 207814 442944
rect 208210 442892 208216 442944
rect 208268 442932 208274 442944
rect 209130 442932 209136 442944
rect 208268 442904 209136 442932
rect 208268 442892 208274 442904
rect 209130 442892 209136 442904
rect 209188 442892 209194 442944
rect 224862 442892 224868 442944
rect 224920 442932 224926 442944
rect 269390 442932 269396 442944
rect 224920 442904 269396 442932
rect 224920 442892 224926 442904
rect 269390 442892 269396 442904
rect 269448 442892 269454 442944
rect 67542 442824 67548 442876
rect 67600 442864 67606 442876
rect 142522 442864 142528 442876
rect 67600 442836 142528 442864
rect 67600 442824 67606 442836
rect 142522 442824 142528 442836
rect 142580 442824 142586 442876
rect 142614 442824 142620 442876
rect 142672 442864 142678 442876
rect 143442 442864 143448 442876
rect 142672 442836 143448 442864
rect 142672 442824 142678 442836
rect 143442 442824 143448 442836
rect 143500 442824 143506 442876
rect 149330 442824 149336 442876
rect 149388 442864 149394 442876
rect 150342 442864 150348 442876
rect 149388 442836 150348 442864
rect 149388 442824 149394 442836
rect 150342 442824 150348 442836
rect 150400 442824 150406 442876
rect 226242 442824 226248 442876
rect 226300 442864 226306 442876
rect 271690 442864 271696 442876
rect 226300 442836 271696 442864
rect 226300 442824 226306 442836
rect 271690 442824 271696 442836
rect 271748 442824 271754 442876
rect 57054 442756 57060 442808
rect 57112 442796 57118 442808
rect 153930 442796 153936 442808
rect 57112 442768 153936 442796
rect 57112 442756 57118 442768
rect 153930 442756 153936 442768
rect 153988 442756 153994 442808
rect 201494 442756 201500 442808
rect 201552 442796 201558 442808
rect 207658 442796 207664 442808
rect 201552 442768 207664 442796
rect 201552 442756 201558 442768
rect 207658 442756 207664 442768
rect 207716 442756 207722 442808
rect 226150 442756 226156 442808
rect 226208 442796 226214 442808
rect 273898 442796 273904 442808
rect 226208 442768 273904 442796
rect 226208 442756 226214 442768
rect 273898 442756 273904 442768
rect 273956 442756 273962 442808
rect 57146 442688 57152 442740
rect 57204 442728 57210 442740
rect 156138 442728 156144 442740
rect 57204 442700 156144 442728
rect 57204 442688 57210 442700
rect 156138 442688 156144 442700
rect 156196 442688 156202 442740
rect 227622 442688 227628 442740
rect 227680 442728 227686 442740
rect 276198 442728 276204 442740
rect 227680 442700 276204 442728
rect 227680 442688 227686 442700
rect 276198 442688 276204 442700
rect 276256 442688 276262 442740
rect 56778 442620 56784 442672
rect 56836 442660 56842 442672
rect 158438 442660 158444 442672
rect 56836 442632 158444 442660
rect 56836 442620 56842 442632
rect 158438 442620 158444 442632
rect 158496 442620 158502 442672
rect 199194 442620 199200 442672
rect 199252 442660 199258 442672
rect 206278 442660 206284 442672
rect 199252 442632 206284 442660
rect 199252 442620 199258 442632
rect 206278 442620 206284 442632
rect 206336 442620 206342 442672
rect 229002 442620 229008 442672
rect 229060 442660 229066 442672
rect 278406 442660 278412 442672
rect 229060 442632 278412 442660
rect 229060 442620 229066 442632
rect 278406 442620 278412 442632
rect 278464 442620 278470 442672
rect 57330 442552 57336 442604
rect 57388 442592 57394 442604
rect 160646 442592 160652 442604
rect 57388 442564 160652 442592
rect 57388 442552 57394 442564
rect 160646 442552 160652 442564
rect 160704 442552 160710 442604
rect 187878 442552 187884 442604
rect 187936 442592 187942 442604
rect 188982 442592 188988 442604
rect 187936 442564 188988 442592
rect 187936 442552 187942 442564
rect 188982 442552 188988 442564
rect 189040 442552 189046 442604
rect 202782 442552 202788 442604
rect 202840 442592 202846 442604
rect 228634 442592 228640 442604
rect 202840 442564 228640 442592
rect 202840 442552 202846 442564
rect 228634 442552 228640 442564
rect 228692 442552 228698 442604
rect 230382 442552 230388 442604
rect 230440 442592 230446 442604
rect 280706 442592 280712 442604
rect 230440 442564 280712 442592
rect 230440 442552 230446 442564
rect 280706 442552 280712 442564
rect 280764 442552 280770 442604
rect 68830 442484 68836 442536
rect 68888 442524 68894 442536
rect 178770 442524 178776 442536
rect 68888 442496 178776 442524
rect 68888 442484 68894 442496
rect 178770 442484 178776 442496
rect 178828 442484 178834 442536
rect 204162 442484 204168 442536
rect 204220 442524 204226 442536
rect 230842 442524 230848 442536
rect 204220 442496 230848 442524
rect 204220 442484 204226 442496
rect 230842 442484 230848 442496
rect 230900 442484 230906 442536
rect 231762 442484 231768 442536
rect 231820 442524 231826 442536
rect 283006 442524 283012 442536
rect 231820 442496 283012 442524
rect 231820 442484 231826 442496
rect 283006 442484 283012 442496
rect 283064 442484 283070 442536
rect 70118 442416 70124 442468
rect 70176 442456 70182 442468
rect 181070 442456 181076 442468
rect 70176 442428 181076 442456
rect 70176 442416 70182 442428
rect 181070 442416 181076 442428
rect 181128 442416 181134 442468
rect 205542 442416 205548 442468
rect 205600 442456 205606 442468
rect 232774 442456 232780 442468
rect 205600 442428 232780 442456
rect 205600 442416 205606 442428
rect 232774 442416 232780 442428
rect 232832 442416 232838 442468
rect 233050 442416 233056 442468
rect 233108 442456 233114 442468
rect 285214 442456 285220 442468
rect 233108 442428 285220 442456
rect 233108 442416 233114 442428
rect 285214 442416 285220 442428
rect 285272 442416 285278 442468
rect 70210 442348 70216 442400
rect 70268 442388 70274 442400
rect 183370 442388 183376 442400
rect 70268 442360 183376 442388
rect 70268 442348 70274 442360
rect 183370 442348 183376 442360
rect 183428 442348 183434 442400
rect 194686 442348 194692 442400
rect 194744 442388 194750 442400
rect 203518 442388 203524 442400
rect 194744 442360 203524 442388
rect 194744 442348 194750 442360
rect 203518 442348 203524 442360
rect 203576 442348 203582 442400
rect 206922 442348 206928 442400
rect 206980 442388 206986 442400
rect 235442 442388 235448 442400
rect 206980 442360 235448 442388
rect 206980 442348 206986 442360
rect 235442 442348 235448 442360
rect 235500 442348 235506 442400
rect 235902 442348 235908 442400
rect 235960 442388 235966 442400
rect 292022 442388 292028 442400
rect 235960 442360 292028 442388
rect 235960 442348 235966 442360
rect 292022 442348 292028 442360
rect 292080 442348 292086 442400
rect 71682 442280 71688 442332
rect 71740 442320 71746 442332
rect 185578 442320 185584 442332
rect 71740 442292 185584 442320
rect 71740 442280 71746 442292
rect 185578 442280 185584 442292
rect 185636 442280 185642 442332
rect 196894 442280 196900 442332
rect 196952 442320 196958 442332
rect 204898 442320 204904 442332
rect 196952 442292 204904 442320
rect 196952 442280 196958 442292
rect 204898 442280 204904 442292
rect 204956 442280 204962 442332
rect 208302 442280 208308 442332
rect 208360 442320 208366 442332
rect 237650 442320 237656 442332
rect 208360 442292 237656 442320
rect 208360 442280 208366 442292
rect 237650 442280 237656 442292
rect 237708 442280 237714 442332
rect 238662 442280 238668 442332
rect 238720 442320 238726 442332
rect 296530 442320 296536 442332
rect 238720 442292 296536 442320
rect 238720 442280 238726 442292
rect 296530 442280 296536 442292
rect 296588 442280 296594 442332
rect 56962 442212 56968 442264
rect 57020 442252 57026 442264
rect 190086 442252 190092 442264
rect 57020 442224 190092 442252
rect 57020 442212 57026 442224
rect 190086 442212 190092 442224
rect 190144 442212 190150 442264
rect 192386 442212 192392 442264
rect 192444 442252 192450 442264
rect 202138 442252 202144 442264
rect 192444 442224 202144 442252
rect 192444 442212 192450 442224
rect 202138 442212 202144 442224
rect 202196 442212 202202 442264
rect 209682 442212 209688 442264
rect 209740 442252 209746 442264
rect 239950 442252 239956 442264
rect 209740 442224 239956 442252
rect 209740 442212 209746 442224
rect 239950 442212 239956 442224
rect 240008 442212 240014 442264
rect 242066 442212 242072 442264
rect 242124 442252 242130 442264
rect 246206 442252 246212 442264
rect 242124 442224 246212 442252
rect 242124 442212 242130 442224
rect 246206 442212 246212 442224
rect 246264 442212 246270 442264
rect 246298 442212 246304 442264
rect 246356 442252 246362 442264
rect 251266 442252 251272 442264
rect 246356 442224 251272 442252
rect 246356 442212 246362 442224
rect 251266 442212 251272 442224
rect 251324 442212 251330 442264
rect 251358 442212 251364 442264
rect 251416 442252 251422 442264
rect 298830 442252 298836 442264
rect 251416 442224 298836 442252
rect 251416 442212 251422 442224
rect 298830 442212 298836 442224
rect 298888 442212 298894 442264
rect 79134 442144 79140 442196
rect 79192 442184 79198 442196
rect 81342 442184 81348 442196
rect 79192 442156 81348 442184
rect 79192 442144 79198 442156
rect 81342 442144 81348 442156
rect 81400 442144 81406 442196
rect 89622 442144 89628 442196
rect 89680 442184 89686 442196
rect 92750 442184 92756 442196
rect 89680 442156 92756 442184
rect 89680 442144 89686 442156
rect 92750 442144 92756 442156
rect 92808 442144 92814 442196
rect 96522 442144 96528 442196
rect 96580 442184 96586 442196
rect 106366 442184 106372 442196
rect 96580 442156 106372 442184
rect 96580 442144 96586 442156
rect 106366 442144 106372 442156
rect 106424 442144 106430 442196
rect 108942 442144 108948 442196
rect 109000 442184 109006 442196
rect 128998 442184 129004 442196
rect 109000 442156 129004 442184
rect 109000 442144 109006 442156
rect 128998 442144 129004 442156
rect 129056 442144 129062 442196
rect 135806 442144 135812 442196
rect 135864 442184 135870 442196
rect 139394 442184 139400 442196
rect 135864 442156 139400 442184
rect 135864 442144 135870 442156
rect 139394 442144 139400 442156
rect 139452 442144 139458 442196
rect 142522 442144 142528 442196
rect 142580 442184 142586 442196
rect 151630 442184 151636 442196
rect 142580 442156 151636 442184
rect 142580 442144 142586 442156
rect 151630 442144 151636 442156
rect 151688 442144 151694 442196
rect 174262 442144 174268 442196
rect 174320 442184 174326 442196
rect 175182 442184 175188 442196
rect 174320 442156 175188 442184
rect 174320 442144 174326 442156
rect 175182 442144 175188 442156
rect 175240 442144 175246 442196
rect 223482 442144 223488 442196
rect 223540 442184 223546 442196
rect 267090 442184 267096 442196
rect 223540 442156 267096 442184
rect 223540 442144 223546 442156
rect 267090 442144 267096 442156
rect 267148 442144 267154 442196
rect 95142 442076 95148 442128
rect 95200 442116 95206 442128
rect 104066 442116 104072 442128
rect 95200 442088 104072 442116
rect 95200 442076 95206 442088
rect 104066 442076 104072 442088
rect 104124 442076 104130 442128
rect 106182 442076 106188 442128
rect 106240 442116 106246 442128
rect 124490 442116 124496 442128
rect 106240 442088 124496 442116
rect 106240 442076 106246 442088
rect 124490 442076 124496 442088
rect 124548 442076 124554 442128
rect 220722 442076 220728 442128
rect 220780 442116 220786 442128
rect 262582 442116 262588 442128
rect 220780 442088 262588 442116
rect 220780 442076 220786 442088
rect 262582 442076 262588 442088
rect 262640 442076 262646 442128
rect 93670 442008 93676 442060
rect 93728 442048 93734 442060
rect 101858 442048 101864 442060
rect 93728 442020 101864 442048
rect 93728 442008 93734 442020
rect 101858 442008 101864 442020
rect 101916 442008 101922 442060
rect 107562 442008 107568 442060
rect 107620 442048 107626 442060
rect 126698 442048 126704 442060
rect 107620 442020 126704 442048
rect 107620 442008 107626 442020
rect 126698 442008 126704 442020
rect 126756 442008 126762 442060
rect 222102 442008 222108 442060
rect 222160 442048 222166 442060
rect 264882 442048 264888 442060
rect 222160 442020 264888 442048
rect 222160 442008 222166 442020
rect 264882 442008 264888 442020
rect 264940 442008 264946 442060
rect 93762 441940 93768 441992
rect 93820 441980 93826 441992
rect 99558 441980 99564 441992
rect 93820 441952 99564 441980
rect 93820 441940 93826 441952
rect 99558 441940 99564 441952
rect 99616 441940 99622 441992
rect 104802 441940 104808 441992
rect 104860 441980 104866 441992
rect 122190 441980 122196 441992
rect 104860 441952 122196 441980
rect 104860 441940 104866 441952
rect 122190 441940 122196 441952
rect 122248 441940 122254 441992
rect 169754 441940 169760 441992
rect 169812 441980 169818 441992
rect 171042 441980 171048 441992
rect 169812 441952 171048 441980
rect 169812 441940 169818 441952
rect 171042 441940 171048 441952
rect 171100 441940 171106 441992
rect 217870 441940 217876 441992
rect 217928 441980 217934 441992
rect 258074 441980 258080 441992
rect 217928 441952 258080 441980
rect 217928 441940 217934 441952
rect 258074 441940 258080 441952
rect 258132 441940 258138 441992
rect 101950 441872 101956 441924
rect 102008 441912 102014 441924
rect 117682 441912 117688 441924
rect 102008 441884 117688 441912
rect 102008 441872 102014 441884
rect 117682 441872 117688 441884
rect 117740 441872 117746 441924
rect 203702 441872 203708 441924
rect 203760 441912 203766 441924
rect 209038 441912 209044 441924
rect 203760 441884 209044 441912
rect 203760 441872 203766 441884
rect 209038 441872 209044 441884
rect 209096 441872 209102 441924
rect 219342 441872 219348 441924
rect 219400 441912 219406 441924
rect 260282 441912 260288 441924
rect 219400 441884 260288 441912
rect 219400 441872 219406 441884
rect 260282 441872 260288 441884
rect 260340 441872 260346 441924
rect 103422 441804 103428 441856
rect 103480 441844 103486 441856
rect 119890 441844 119896 441856
rect 103480 441816 119896 441844
rect 103480 441804 103486 441816
rect 119890 441804 119896 441816
rect 119948 441804 119954 441856
rect 213822 441804 213828 441856
rect 213880 441844 213886 441856
rect 213880 441816 244872 441844
rect 213880 441804 213886 441816
rect 91002 441736 91008 441788
rect 91060 441776 91066 441788
rect 95050 441776 95056 441788
rect 91060 441748 95056 441776
rect 91060 441736 91066 441748
rect 95050 441736 95056 441748
rect 95108 441736 95114 441788
rect 100662 441736 100668 441788
rect 100720 441776 100726 441788
rect 113174 441776 113180 441788
rect 100720 441748 113180 441776
rect 100720 441736 100726 441748
rect 113174 441736 113180 441748
rect 113232 441736 113238 441788
rect 211062 441736 211068 441788
rect 211120 441776 211126 441788
rect 244458 441776 244464 441788
rect 211120 441748 244464 441776
rect 211120 441736 211126 441748
rect 244458 441736 244464 441748
rect 244516 441736 244522 441788
rect 244844 441776 244872 441816
rect 244918 441804 244924 441856
rect 244976 441844 244982 441856
rect 253566 441844 253572 441856
rect 244976 441816 253572 441844
rect 244976 441804 244982 441816
rect 253566 441804 253572 441816
rect 253624 441804 253630 441856
rect 248598 441776 248604 441788
rect 244844 441748 248604 441776
rect 248598 441736 248604 441748
rect 248656 441736 248662 441788
rect 248690 441736 248696 441788
rect 248748 441776 248754 441788
rect 251358 441776 251364 441788
rect 248748 441748 251364 441776
rect 248748 441736 248754 441748
rect 251358 441736 251364 441748
rect 251416 441736 251422 441788
rect 102042 441668 102048 441720
rect 102100 441708 102106 441720
rect 115382 441708 115388 441720
rect 102100 441680 115388 441708
rect 102100 441668 102106 441680
rect 115382 441668 115388 441680
rect 115440 441668 115446 441720
rect 212442 441668 212448 441720
rect 212500 441708 212506 441720
rect 242066 441708 242072 441720
rect 212500 441680 242072 441708
rect 212500 441668 212506 441680
rect 242066 441668 242072 441680
rect 242124 441668 242130 441720
rect 99282 441600 99288 441652
rect 99340 441640 99346 441652
rect 110874 441640 110880 441652
rect 99340 441612 110880 441640
rect 99340 441600 99346 441612
rect 110874 441600 110880 441612
rect 110932 441600 110938 441652
rect 210970 441600 210976 441652
rect 211028 441640 211034 441652
rect 242250 441640 242256 441652
rect 211028 441612 242256 441640
rect 211028 441600 211034 441612
rect 242250 441600 242256 441612
rect 242308 441600 242314 441652
rect 245102 441600 245108 441652
rect 245160 441640 245166 441652
rect 255774 441640 255780 441652
rect 245160 441612 255780 441640
rect 245160 441600 245166 441612
rect 255774 441600 255780 441612
rect 255832 441600 255838 441652
rect 56962 439832 56968 439884
rect 57020 439872 57026 439884
rect 136358 439872 136364 439884
rect 57020 439844 136364 439872
rect 57020 439832 57026 439844
rect 136358 439832 136364 439844
rect 136416 439832 136422 439884
rect 56778 439764 56784 439816
rect 56836 439804 56842 439816
rect 136450 439804 136456 439816
rect 56836 439776 136456 439804
rect 56836 439764 56842 439776
rect 136450 439764 136456 439776
rect 136508 439764 136514 439816
rect 56870 439696 56876 439748
rect 56928 439736 56934 439748
rect 299658 439736 299664 439748
rect 56928 439708 299664 439736
rect 56928 439696 56934 439708
rect 299658 439696 299664 439708
rect 299716 439696 299722 439748
rect 57054 439628 57060 439680
rect 57112 439668 57118 439680
rect 429378 439668 429384 439680
rect 57112 439640 429384 439668
rect 57112 439628 57118 439640
rect 429378 439628 429384 439640
rect 429436 439628 429442 439680
rect 57974 439560 57980 439612
rect 58032 439600 58038 439612
rect 580350 439600 580356 439612
rect 58032 439572 580356 439600
rect 58032 439560 58038 439572
rect 580350 439560 580356 439572
rect 580408 439560 580414 439612
rect 58066 439492 58072 439544
rect 58124 439532 58130 439544
rect 580718 439532 580724 439544
rect 58124 439504 580724 439532
rect 58124 439492 58130 439504
rect 580718 439492 580724 439504
rect 580776 439492 580782 439544
rect 58158 438948 58164 439000
rect 58216 438988 58222 439000
rect 580074 438988 580080 439000
rect 58216 438960 580080 438988
rect 58216 438948 58222 438960
rect 580074 438948 580080 438960
rect 580132 438948 580138 439000
rect 48958 438880 48964 438932
rect 49016 438920 49022 438932
rect 56594 438920 56600 438932
rect 49016 438892 56600 438920
rect 49016 438880 49022 438892
rect 56594 438880 56600 438892
rect 56652 438880 56658 438932
rect 57514 438880 57520 438932
rect 57572 438920 57578 438932
rect 580626 438920 580632 438932
rect 57572 438892 580632 438920
rect 57572 438880 57578 438892
rect 580626 438880 580632 438892
rect 580684 438880 580690 438932
rect 57238 438268 57244 438320
rect 57296 438308 57302 438320
rect 580534 438308 580540 438320
rect 57296 438280 580540 438308
rect 57296 438268 57302 438280
rect 580534 438268 580540 438280
rect 580592 438268 580598 438320
rect 57330 438200 57336 438252
rect 57388 438240 57394 438252
rect 580810 438240 580816 438252
rect 57388 438212 580816 438240
rect 57388 438200 57394 438212
rect 580810 438200 580816 438212
rect 580868 438200 580874 438252
rect 56686 438132 56692 438184
rect 56744 438172 56750 438184
rect 580258 438172 580264 438184
rect 56744 438144 580264 438172
rect 56744 438132 56750 438144
rect 580258 438132 580264 438144
rect 580316 438132 580322 438184
rect 59998 437996 60004 438048
rect 60056 438036 60062 438048
rect 580350 438036 580356 438048
rect 60056 438008 580356 438036
rect 60056 437996 60062 438008
rect 580350 437996 580356 438008
rect 580408 437996 580414 438048
rect 57422 437928 57428 437980
rect 57480 437968 57486 437980
rect 580442 437968 580448 437980
rect 57480 437940 580448 437968
rect 57480 437928 57486 437940
rect 580442 437928 580448 437940
rect 580500 437928 580506 437980
rect 302786 437384 302792 437436
rect 302844 437424 302850 437436
rect 467098 437424 467104 437436
rect 302844 437396 467104 437424
rect 302844 437384 302850 437396
rect 467098 437384 467104 437396
rect 467156 437384 467162 437436
rect 51718 436092 51724 436144
rect 51776 436132 51782 436144
rect 56594 436132 56600 436144
rect 51776 436104 56600 436132
rect 51776 436092 51782 436104
rect 56594 436092 56600 436104
rect 56652 436092 56658 436144
rect 15838 434732 15844 434784
rect 15896 434772 15902 434784
rect 56686 434772 56692 434784
rect 15896 434744 56692 434772
rect 15896 434732 15902 434744
rect 56686 434732 56692 434744
rect 56744 434732 56750 434784
rect 302786 434664 302792 434716
rect 302844 434704 302850 434716
rect 323486 434704 323492 434716
rect 302844 434676 323492 434704
rect 302844 434664 302850 434676
rect 323486 434664 323492 434676
rect 323544 434664 323550 434716
rect 327534 434664 327540 434716
rect 327592 434704 327598 434716
rect 327626 434704 327632 434716
rect 327592 434676 327632 434704
rect 327592 434664 327598 434676
rect 327626 434664 327632 434676
rect 327684 434664 327690 434716
rect 327718 434664 327724 434716
rect 327776 434704 327782 434716
rect 465718 434704 465724 434716
rect 327776 434676 465724 434704
rect 327776 434664 327782 434676
rect 465718 434664 465724 434676
rect 465776 434664 465782 434716
rect 323486 434460 323492 434512
rect 323544 434500 323550 434512
rect 327718 434500 327724 434512
rect 323544 434472 327724 434500
rect 323544 434460 323550 434472
rect 327718 434460 327724 434472
rect 327776 434460 327782 434512
rect 302786 433236 302792 433288
rect 302844 433276 302850 433288
rect 464338 433276 464344 433288
rect 302844 433248 464344 433276
rect 302844 433236 302850 433248
rect 464338 433236 464344 433248
rect 464396 433236 464402 433288
rect 39298 431944 39304 431996
rect 39356 431984 39362 431996
rect 56686 431984 56692 431996
rect 39356 431956 56692 431984
rect 39356 431944 39362 431956
rect 56686 431944 56692 431956
rect 56744 431944 56750 431996
rect 302786 430516 302792 430568
rect 302844 430556 302850 430568
rect 354030 430556 354036 430568
rect 302844 430528 354036 430556
rect 302844 430516 302850 430528
rect 354030 430516 354036 430528
rect 354088 430516 354094 430568
rect 46198 429156 46204 429208
rect 46256 429196 46262 429208
rect 57146 429196 57152 429208
rect 46256 429168 57152 429196
rect 46256 429156 46262 429168
rect 57146 429156 57152 429168
rect 57204 429156 57210 429208
rect 302786 429088 302792 429140
rect 302844 429128 302850 429140
rect 353938 429128 353944 429140
rect 302844 429100 353944 429128
rect 302844 429088 302850 429100
rect 353938 429088 353944 429100
rect 353996 429088 354002 429140
rect 10318 427796 10324 427848
rect 10376 427836 10382 427848
rect 57146 427836 57152 427848
rect 10376 427808 57152 427836
rect 10376 427796 10382 427808
rect 57146 427796 57152 427808
rect 57204 427796 57210 427848
rect 302786 426368 302792 426420
rect 302844 426408 302850 426420
rect 352742 426408 352748 426420
rect 302844 426380 352748 426408
rect 302844 426368 302850 426380
rect 352742 426368 352748 426380
rect 352800 426368 352806 426420
rect 17218 425076 17224 425128
rect 17276 425116 17282 425128
rect 57146 425116 57152 425128
rect 17276 425088 57152 425116
rect 17276 425076 17282 425088
rect 57146 425076 57152 425088
rect 57204 425076 57210 425128
rect 43438 423648 43444 423700
rect 43496 423688 43502 423700
rect 57146 423688 57152 423700
rect 43496 423660 57152 423688
rect 43496 423648 43502 423660
rect 57146 423648 57152 423660
rect 57204 423648 57210 423700
rect 327534 423648 327540 423700
rect 327592 423688 327598 423700
rect 327626 423688 327632 423700
rect 327592 423660 327632 423688
rect 327592 423648 327598 423660
rect 327626 423648 327632 423660
rect 327684 423648 327690 423700
rect 302786 423580 302792 423632
rect 302844 423620 302850 423632
rect 352650 423620 352656 423632
rect 302844 423592 352656 423620
rect 302844 423580 302850 423592
rect 352650 423580 352656 423592
rect 352708 423580 352714 423632
rect 302786 422220 302792 422272
rect 302844 422260 302850 422272
rect 352558 422260 352564 422272
rect 302844 422232 352564 422260
rect 302844 422220 302850 422232
rect 352558 422220 352564 422232
rect 352616 422220 352622 422272
rect 4890 420928 4896 420980
rect 4948 420968 4954 420980
rect 57146 420968 57152 420980
rect 4948 420940 57152 420968
rect 4948 420928 4954 420940
rect 57146 420928 57152 420940
rect 57204 420928 57210 420980
rect 19978 419500 19984 419552
rect 20036 419540 20042 419552
rect 57146 419540 57152 419552
rect 20036 419512 57152 419540
rect 20036 419500 20042 419512
rect 57146 419500 57152 419512
rect 57204 419500 57210 419552
rect 302786 419432 302792 419484
rect 302844 419472 302850 419484
rect 351178 419472 351184 419484
rect 302844 419444 351184 419472
rect 302844 419432 302850 419444
rect 351178 419432 351184 419444
rect 351236 419432 351242 419484
rect 302786 418072 302792 418124
rect 302844 418112 302850 418124
rect 349798 418112 349804 418124
rect 302844 418084 349804 418112
rect 302844 418072 302850 418084
rect 349798 418072 349804 418084
rect 349856 418072 349862 418124
rect 33778 416780 33784 416832
rect 33836 416820 33842 416832
rect 57146 416820 57152 416832
rect 33836 416792 57152 416820
rect 33836 416780 33842 416792
rect 57146 416780 57152 416792
rect 57204 416780 57210 416832
rect 5074 415420 5080 415472
rect 5132 415460 5138 415472
rect 57146 415460 57152 415472
rect 5132 415432 57152 415460
rect 5132 415420 5138 415432
rect 57146 415420 57152 415432
rect 57204 415420 57210 415472
rect 302786 415352 302792 415404
rect 302844 415392 302850 415404
rect 347038 415392 347044 415404
rect 302844 415364 347044 415392
rect 302844 415352 302850 415364
rect 347038 415352 347044 415364
rect 347096 415352 347102 415404
rect 327534 413924 327540 413976
rect 327592 413964 327598 413976
rect 327718 413964 327724 413976
rect 327592 413936 327724 413964
rect 327592 413924 327598 413936
rect 327718 413924 327724 413936
rect 327776 413924 327782 413976
rect 53098 412632 53104 412684
rect 53156 412672 53162 412684
rect 57146 412672 57152 412684
rect 53156 412644 57152 412672
rect 53156 412632 53162 412644
rect 57146 412632 57152 412644
rect 57204 412632 57210 412684
rect 302786 412564 302792 412616
rect 302844 412604 302850 412616
rect 476206 412604 476212 412616
rect 302844 412576 476212 412604
rect 302844 412564 302850 412576
rect 476206 412564 476212 412576
rect 476264 412564 476270 412616
rect 31018 411272 31024 411324
rect 31076 411312 31082 411324
rect 57146 411312 57152 411324
rect 31076 411284 57152 411312
rect 31076 411272 31082 411284
rect 57146 411272 57152 411284
rect 57204 411272 57210 411324
rect 302786 411204 302792 411256
rect 302844 411244 302850 411256
rect 474734 411244 474740 411256
rect 302844 411216 474740 411244
rect 302844 411204 302850 411216
rect 474734 411204 474740 411216
rect 474792 411204 474798 411256
rect 3510 408484 3516 408536
rect 3568 408524 3574 408536
rect 57146 408524 57152 408536
rect 3568 408496 57152 408524
rect 3568 408484 3574 408496
rect 57146 408484 57152 408496
rect 57204 408484 57210 408536
rect 302786 408416 302792 408468
rect 302844 408456 302850 408468
rect 473354 408456 473360 408468
rect 302844 408428 473360 408456
rect 302844 408416 302850 408428
rect 473354 408416 473360 408428
rect 473412 408416 473418 408468
rect 37918 407124 37924 407176
rect 37976 407164 37982 407176
rect 57146 407164 57152 407176
rect 37976 407136 57152 407164
rect 37976 407124 37982 407136
rect 57146 407124 57152 407136
rect 57204 407124 57210 407176
rect 302786 407056 302792 407108
rect 302844 407096 302850 407108
rect 471974 407096 471980 407108
rect 302844 407068 471980 407096
rect 302844 407056 302850 407068
rect 471974 407056 471980 407068
rect 472032 407056 472038 407108
rect 5166 404336 5172 404388
rect 5224 404376 5230 404388
rect 57146 404376 57152 404388
rect 5224 404348 57152 404376
rect 5224 404336 5230 404348
rect 57146 404336 57152 404348
rect 57204 404336 57210 404388
rect 327534 404336 327540 404388
rect 327592 404376 327598 404388
rect 327718 404376 327724 404388
rect 327592 404348 327724 404376
rect 327592 404336 327598 404348
rect 327718 404336 327724 404348
rect 327776 404336 327782 404388
rect 302694 404268 302700 404320
rect 302752 404308 302758 404320
rect 470594 404308 470600 404320
rect 302752 404280 470600 404308
rect 302752 404268 302758 404280
rect 470594 404268 470600 404280
rect 470652 404268 470658 404320
rect 302786 401548 302792 401600
rect 302844 401588 302850 401600
rect 469214 401588 469220 401600
rect 302844 401560 469220 401588
rect 302844 401548 302850 401560
rect 469214 401548 469220 401560
rect 469272 401548 469278 401600
rect 35158 400188 35164 400240
rect 35216 400228 35222 400240
rect 56686 400228 56692 400240
rect 35216 400200 56692 400228
rect 35216 400188 35222 400200
rect 56686 400188 56692 400200
rect 56744 400188 56750 400240
rect 302786 400120 302792 400172
rect 302844 400160 302850 400172
rect 467926 400160 467932 400172
rect 302844 400132 467932 400160
rect 302844 400120 302850 400132
rect 467926 400120 467932 400132
rect 467984 400120 467990 400172
rect 5258 398828 5264 398880
rect 5316 398868 5322 398880
rect 56686 398868 56692 398880
rect 5316 398840 56692 398868
rect 5316 398828 5322 398840
rect 56686 398828 56692 398840
rect 56744 398828 56750 398880
rect 302786 397400 302792 397452
rect 302844 397440 302850 397452
rect 467834 397440 467840 397452
rect 302844 397412 467840 397440
rect 302844 397400 302850 397412
rect 467834 397400 467840 397412
rect 467892 397400 467898 397452
rect 302510 395972 302516 396024
rect 302568 396012 302574 396024
rect 466454 396012 466460 396024
rect 302568 395984 466460 396012
rect 302568 395972 302574 395984
rect 466454 395972 466460 395984
rect 466512 395972 466518 396024
rect 2774 394748 2780 394800
rect 2832 394788 2838 394800
rect 5350 394788 5356 394800
rect 2832 394760 5356 394788
rect 2832 394748 2838 394760
rect 5350 394748 5356 394760
rect 5408 394748 5414 394800
rect 4062 394680 4068 394732
rect 4120 394720 4126 394732
rect 56502 394720 56508 394732
rect 4120 394692 56508 394720
rect 4120 394680 4126 394692
rect 56502 394680 56508 394692
rect 56560 394680 56566 394732
rect 327534 394612 327540 394664
rect 327592 394652 327598 394664
rect 327626 394652 327632 394664
rect 327592 394624 327632 394652
rect 327592 394612 327598 394624
rect 327626 394612 327632 394624
rect 327684 394612 327690 394664
rect 302694 393252 302700 393304
rect 302752 393292 302758 393304
rect 465074 393292 465080 393304
rect 302752 393264 465080 393292
rect 302752 393252 302758 393264
rect 465074 393252 465080 393264
rect 465132 393252 465138 393304
rect 3878 391960 3884 392012
rect 3936 392000 3942 392012
rect 56594 392000 56600 392012
rect 3936 391972 56600 392000
rect 3936 391960 3942 391972
rect 56594 391960 56600 391972
rect 56652 391960 56658 392012
rect 302786 390464 302792 390516
rect 302844 390504 302850 390516
rect 463694 390504 463700 390516
rect 302844 390476 463700 390504
rect 302844 390464 302850 390476
rect 463694 390464 463700 390476
rect 463752 390464 463758 390516
rect 3234 389172 3240 389224
rect 3292 389212 3298 389224
rect 56594 389212 56600 389224
rect 3292 389184 56600 389212
rect 3292 389172 3298 389184
rect 56594 389172 56600 389184
rect 56652 389172 56658 389224
rect 302786 389104 302792 389156
rect 302844 389144 302850 389156
rect 462314 389144 462320 389156
rect 302844 389116 462320 389144
rect 302844 389104 302850 389116
rect 462314 389104 462320 389116
rect 462372 389104 462378 389156
rect 302510 386316 302516 386368
rect 302568 386356 302574 386368
rect 461026 386356 461032 386368
rect 302568 386328 461032 386356
rect 302568 386316 302574 386328
rect 461026 386316 461032 386328
rect 461084 386316 461090 386368
rect 3050 385024 3056 385076
rect 3108 385064 3114 385076
rect 56594 385064 56600 385076
rect 3108 385036 56600 385064
rect 3108 385024 3114 385036
rect 56594 385024 56600 385036
rect 56652 385024 56658 385076
rect 327626 385024 327632 385076
rect 327684 385064 327690 385076
rect 327810 385064 327816 385076
rect 327684 385036 327816 385064
rect 327684 385024 327690 385036
rect 327810 385024 327816 385036
rect 327868 385024 327874 385076
rect 302510 384956 302516 385008
rect 302568 384996 302574 385008
rect 460934 384996 460940 385008
rect 302568 384968 460940 384996
rect 302568 384956 302574 384968
rect 460934 384956 460940 384968
rect 460992 384956 460998 385008
rect 22094 384888 22100 384940
rect 22152 384928 22158 384940
rect 38654 384928 38660 384940
rect 22152 384900 38660 384928
rect 22152 384888 22158 384900
rect 38654 384888 38660 384900
rect 38712 384888 38718 384940
rect 42886 384888 42892 384940
rect 42944 384928 42950 384940
rect 42944 384900 51028 384928
rect 42944 384888 42950 384900
rect 5350 384820 5356 384872
rect 5408 384860 5414 384872
rect 19334 384860 19340 384872
rect 5408 384832 19340 384860
rect 5408 384820 5414 384832
rect 19334 384820 19340 384832
rect 19392 384820 19398 384872
rect 51000 384792 51028 384900
rect 56594 384792 56600 384804
rect 51000 384764 56600 384792
rect 56594 384752 56600 384764
rect 56652 384752 56658 384804
rect 3326 382168 3332 382220
rect 3384 382208 3390 382220
rect 56594 382208 56600 382220
rect 3384 382180 56600 382208
rect 3384 382168 3390 382180
rect 56594 382168 56600 382180
rect 56652 382168 56658 382220
rect 302786 382168 302792 382220
rect 302844 382208 302850 382220
rect 443638 382208 443644 382220
rect 302844 382180 443644 382208
rect 302844 382168 302850 382180
rect 443638 382168 443644 382180
rect 443696 382168 443702 382220
rect 302602 380808 302608 380860
rect 302660 380848 302666 380860
rect 359458 380848 359464 380860
rect 302660 380820 359464 380848
rect 302660 380808 302666 380820
rect 359458 380808 359464 380820
rect 359516 380808 359522 380860
rect 3326 380740 3332 380792
rect 3384 380780 3390 380792
rect 56594 380780 56600 380792
rect 3384 380752 56600 380780
rect 3384 380740 3390 380752
rect 56594 380740 56600 380752
rect 56652 380740 56658 380792
rect 3142 380604 3148 380656
rect 3200 380644 3206 380656
rect 56594 380644 56600 380656
rect 3200 380616 56600 380644
rect 3200 380604 3206 380616
rect 56594 380604 56600 380616
rect 56652 380604 56658 380656
rect 3970 378088 3976 378140
rect 4028 378128 4034 378140
rect 56594 378128 56600 378140
rect 4028 378100 56600 378128
rect 4028 378088 4034 378100
rect 56594 378088 56600 378100
rect 56652 378088 56658 378140
rect 302786 378088 302792 378140
rect 302844 378128 302850 378140
rect 358078 378128 358084 378140
rect 302844 378100 358084 378128
rect 302844 378088 302850 378100
rect 358078 378088 358084 378100
rect 358136 378088 358142 378140
rect 327626 376728 327632 376780
rect 327684 376768 327690 376780
rect 327810 376768 327816 376780
rect 327684 376740 327816 376768
rect 327684 376728 327690 376740
rect 327810 376728 327816 376740
rect 327868 376728 327874 376780
rect 3786 376660 3792 376712
rect 3844 376700 3850 376712
rect 56594 376700 56600 376712
rect 3844 376672 56600 376700
rect 3844 376660 3850 376672
rect 56594 376660 56600 376672
rect 56652 376660 56658 376712
rect 302786 375300 302792 375352
rect 302844 375340 302850 375352
rect 356698 375340 356704 375352
rect 302844 375312 356704 375340
rect 302844 375300 302850 375312
rect 356698 375300 356704 375312
rect 356756 375300 356762 375352
rect 20070 373940 20076 373992
rect 20128 373980 20134 373992
rect 56594 373980 56600 373992
rect 20128 373952 56600 373980
rect 20128 373940 20134 373952
rect 56594 373940 56600 373952
rect 56652 373940 56658 373992
rect 302786 373940 302792 373992
rect 302844 373980 302850 373992
rect 355318 373980 355324 373992
rect 302844 373952 355324 373980
rect 302844 373940 302850 373952
rect 355318 373940 355324 373952
rect 355376 373940 355382 373992
rect 3694 372512 3700 372564
rect 3752 372552 3758 372564
rect 56594 372552 56600 372564
rect 3752 372524 56600 372552
rect 3752 372512 3758 372524
rect 56594 372512 56600 372524
rect 56652 372512 56658 372564
rect 302326 371152 302332 371204
rect 302384 371192 302390 371204
rect 342898 371192 342904 371204
rect 302384 371164 342904 371192
rect 302384 371152 302390 371164
rect 342898 371152 342904 371164
rect 342956 371152 342962 371204
rect 32398 369792 32404 369844
rect 32456 369832 32462 369844
rect 56594 369832 56600 369844
rect 32456 369804 56600 369832
rect 32456 369792 32462 369804
rect 56594 369792 56600 369804
rect 56652 369792 56658 369844
rect 302602 369792 302608 369844
rect 302660 369832 302666 369844
rect 452746 369832 452752 369844
rect 302660 369804 452752 369832
rect 302660 369792 302666 369804
rect 452746 369792 452752 369804
rect 452804 369792 452810 369844
rect 3602 368432 3608 368484
rect 3660 368472 3666 368484
rect 56594 368472 56600 368484
rect 3660 368444 56600 368472
rect 3660 368432 3666 368444
rect 56594 368432 56600 368444
rect 56652 368432 56658 368484
rect 302786 367004 302792 367056
rect 302844 367044 302850 367056
rect 330478 367044 330484 367056
rect 302844 367016 330484 367044
rect 302844 367004 302850 367016
rect 330478 367004 330484 367016
rect 330536 367004 330542 367056
rect 3418 365644 3424 365696
rect 3476 365684 3482 365696
rect 56594 365684 56600 365696
rect 3476 365656 56600 365684
rect 3476 365644 3482 365656
rect 56594 365644 56600 365656
rect 56652 365644 56658 365696
rect 28258 364284 28264 364336
rect 28316 364324 28322 364336
rect 56594 364324 56600 364336
rect 28316 364296 56600 364324
rect 28316 364284 28322 364296
rect 56594 364284 56600 364296
rect 56652 364284 56658 364336
rect 302510 364284 302516 364336
rect 302568 364324 302574 364336
rect 329282 364324 329288 364336
rect 302568 364296 329288 364324
rect 302568 364284 302574 364296
rect 329282 364284 329288 364296
rect 329340 364284 329346 364336
rect 302418 362856 302424 362908
rect 302476 362896 302482 362908
rect 329098 362896 329104 362908
rect 302476 362868 329104 362896
rect 302476 362856 302482 362868
rect 329098 362856 329104 362868
rect 329156 362856 329162 362908
rect 17310 361496 17316 361548
rect 17368 361536 17374 361548
rect 56594 361536 56600 361548
rect 17368 361508 56600 361536
rect 17368 361496 17374 361508
rect 56594 361496 56600 361508
rect 56652 361496 56658 361548
rect 4982 360136 4988 360188
rect 5040 360176 5046 360188
rect 56594 360176 56600 360188
rect 5040 360148 56600 360176
rect 5040 360136 5046 360148
rect 56594 360136 56600 360148
rect 56652 360136 56658 360188
rect 302326 360136 302332 360188
rect 302384 360176 302390 360188
rect 328086 360176 328092 360188
rect 302384 360148 328092 360176
rect 302384 360136 302390 360148
rect 328086 360136 328092 360148
rect 328144 360136 328150 360188
rect 302510 358708 302516 358760
rect 302568 358748 302574 358760
rect 326338 358748 326344 358760
rect 302568 358720 326344 358748
rect 302568 358708 302574 358720
rect 326338 358708 326344 358720
rect 326396 358708 326402 358760
rect 21358 357348 21364 357400
rect 21416 357388 21422 357400
rect 56594 357388 56600 357400
rect 21416 357360 56600 357388
rect 21416 357348 21422 357360
rect 56594 357348 56600 357360
rect 56652 357348 56658 357400
rect 14458 355988 14464 356040
rect 14516 356028 14522 356040
rect 56594 356028 56600 356040
rect 14516 356000 56600 356028
rect 14516 355988 14522 356000
rect 56594 355988 56600 356000
rect 56652 355988 56658 356040
rect 302786 355988 302792 356040
rect 302844 356028 302850 356040
rect 324958 356028 324964 356040
rect 302844 356000 324964 356028
rect 302844 355988 302850 356000
rect 324958 355988 324964 356000
rect 325016 355988 325022 356040
rect 4798 353200 4804 353252
rect 4856 353240 4862 353252
rect 56594 353240 56600 353252
rect 4856 353212 56600 353240
rect 4856 353200 4862 353212
rect 56594 353200 56600 353212
rect 56652 353200 56658 353252
rect 302786 353200 302792 353252
rect 302844 353240 302850 353252
rect 323578 353240 323584 353252
rect 302844 353212 323584 353240
rect 302844 353200 302850 353212
rect 323578 353200 323584 353212
rect 323636 353200 323642 353252
rect 24762 351840 24768 351892
rect 24820 351880 24826 351892
rect 56594 351880 56600 351892
rect 24820 351852 56600 351880
rect 24820 351840 24826 351852
rect 56594 351840 56600 351852
rect 56652 351840 56658 351892
rect 302418 351840 302424 351892
rect 302476 351880 302482 351892
rect 322198 351880 322204 351892
rect 302476 351852 322204 351880
rect 302476 351840 302482 351852
rect 322198 351840 322204 351852
rect 322256 351840 322262 351892
rect 13078 349052 13084 349104
rect 13136 349092 13142 349104
rect 56594 349092 56600 349104
rect 13136 349064 56600 349092
rect 13136 349052 13142 349064
rect 56594 349052 56600 349064
rect 56652 349052 56658 349104
rect 302694 349052 302700 349104
rect 302752 349092 302758 349104
rect 460382 349092 460388 349104
rect 302752 349064 460388 349092
rect 302752 349052 302758 349064
rect 460382 349052 460388 349064
rect 460440 349052 460446 349104
rect 302510 347692 302516 347744
rect 302568 347732 302574 347744
rect 460198 347732 460204 347744
rect 302568 347704 460204 347732
rect 302568 347692 302574 347704
rect 460198 347692 460204 347704
rect 460256 347692 460262 347744
rect 42058 346332 42064 346384
rect 42116 346372 42122 346384
rect 56594 346372 56600 346384
rect 42116 346344 56600 346372
rect 42116 346332 42122 346344
rect 56594 346332 56600 346344
rect 56652 346332 56658 346384
rect 302786 344972 302792 345024
rect 302844 345012 302850 345024
rect 458818 345012 458824 345024
rect 302844 344984 458824 345012
rect 302844 344972 302850 344984
rect 458818 344972 458824 344984
rect 458876 344972 458882 345024
rect 302786 342184 302792 342236
rect 302844 342224 302850 342236
rect 457438 342224 457444 342236
rect 302844 342196 457444 342224
rect 302844 342184 302850 342196
rect 457438 342184 457444 342196
rect 457496 342184 457502 342236
rect 302418 340824 302424 340876
rect 302476 340864 302482 340876
rect 456058 340864 456064 340876
rect 302476 340836 456064 340864
rect 302476 340824 302482 340836
rect 456058 340824 456064 340836
rect 456116 340824 456122 340876
rect 302694 338036 302700 338088
rect 302752 338076 302758 338088
rect 454678 338076 454684 338088
rect 302752 338048 454684 338076
rect 302752 338036 302758 338048
rect 454678 338036 454684 338048
rect 454736 338036 454742 338088
rect 302510 336676 302516 336728
rect 302568 336716 302574 336728
rect 453482 336716 453488 336728
rect 302568 336688 453488 336716
rect 302568 336676 302574 336688
rect 453482 336676 453488 336688
rect 453540 336676 453546 336728
rect 302786 333888 302792 333940
rect 302844 333928 302850 333940
rect 453298 333928 453304 333940
rect 302844 333900 453304 333928
rect 302844 333888 302850 333900
rect 453298 333888 453304 333900
rect 453356 333888 453362 333940
rect 302510 331100 302516 331152
rect 302568 331140 302574 331152
rect 305822 331140 305828 331152
rect 302568 331112 305828 331140
rect 302568 331100 302574 331112
rect 305822 331100 305828 331112
rect 305880 331100 305886 331152
rect 302326 329400 302332 329452
rect 302384 329440 302390 329452
rect 304442 329440 304448 329452
rect 302384 329412 304448 329440
rect 302384 329400 302390 329412
rect 304442 329400 304448 329412
rect 304500 329400 304506 329452
rect 302510 326884 302516 326936
rect 302568 326924 302574 326936
rect 305730 326924 305736 326936
rect 302568 326896 305736 326924
rect 302568 326884 302574 326896
rect 305730 326884 305736 326896
rect 305788 326884 305794 326936
rect 302326 324436 302332 324488
rect 302384 324476 302390 324488
rect 304350 324476 304356 324488
rect 302384 324448 304356 324476
rect 302384 324436 302390 324448
rect 304350 324436 304356 324448
rect 304408 324436 304414 324488
rect 302326 322668 302332 322720
rect 302384 322708 302390 322720
rect 305638 322708 305644 322720
rect 302384 322680 305644 322708
rect 302384 322668 302390 322680
rect 305638 322668 305644 322680
rect 305696 322668 305702 322720
rect 302326 320084 302332 320136
rect 302384 320124 302390 320136
rect 304258 320124 304264 320136
rect 302384 320096 304264 320124
rect 302384 320084 302390 320096
rect 304258 320084 304264 320096
rect 304316 320084 304322 320136
rect 57790 319472 57796 319524
rect 57848 319512 57854 319524
rect 59998 319512 60004 319524
rect 57848 319484 60004 319512
rect 57848 319472 57854 319484
rect 59998 319472 60004 319484
rect 60056 319472 60062 319524
rect 302694 318316 302700 318368
rect 302752 318356 302758 318368
rect 307018 318356 307024 318368
rect 302752 318328 307024 318356
rect 302752 318316 302758 318328
rect 307018 318316 307024 318328
rect 307076 318316 307082 318368
rect 302786 315936 302792 315988
rect 302844 315976 302850 315988
rect 316034 315976 316040 315988
rect 302844 315948 316040 315976
rect 302844 315936 302850 315948
rect 316034 315936 316040 315948
rect 316092 315936 316098 315988
rect 302786 314576 302792 314628
rect 302844 314616 302850 314628
rect 399478 314616 399484 314628
rect 302844 314588 399484 314616
rect 302844 314576 302850 314588
rect 399478 314576 399484 314588
rect 399536 314576 399542 314628
rect 302694 311788 302700 311840
rect 302752 311828 302758 311840
rect 398098 311828 398104 311840
rect 302752 311800 398104 311828
rect 302752 311788 302758 311800
rect 398098 311788 398104 311800
rect 398156 311788 398162 311840
rect 302786 309068 302792 309120
rect 302844 309108 302850 309120
rect 395338 309108 395344 309120
rect 302844 309080 395344 309108
rect 302844 309068 302850 309080
rect 395338 309068 395344 309080
rect 395396 309068 395402 309120
rect 302786 307708 302792 307760
rect 302844 307748 302850 307760
rect 393958 307748 393964 307760
rect 302844 307720 393964 307748
rect 302844 307708 302850 307720
rect 393958 307708 393964 307720
rect 394016 307708 394022 307760
rect 302786 304920 302792 304972
rect 302844 304960 302850 304972
rect 392578 304960 392584 304972
rect 302844 304932 392584 304960
rect 302844 304920 302850 304932
rect 392578 304920 392584 304932
rect 392636 304920 392642 304972
rect 302786 303560 302792 303612
rect 302844 303600 302850 303612
rect 391198 303600 391204 303612
rect 302844 303572 391204 303600
rect 302844 303560 302850 303572
rect 391198 303560 391204 303572
rect 391256 303560 391262 303612
rect 302694 300772 302700 300824
rect 302752 300812 302758 300824
rect 388438 300812 388444 300824
rect 302752 300784 388444 300812
rect 302752 300772 302758 300784
rect 388438 300772 388444 300784
rect 388496 300772 388502 300824
rect 302786 298052 302792 298104
rect 302844 298092 302850 298104
rect 445754 298092 445760 298104
rect 302844 298064 445760 298092
rect 302844 298052 302850 298064
rect 445754 298052 445760 298064
rect 445812 298052 445818 298104
rect 302602 295876 302608 295928
rect 302660 295916 302666 295928
rect 305914 295916 305920 295928
rect 302660 295888 305920 295916
rect 302660 295876 302666 295888
rect 305914 295876 305920 295888
rect 305972 295876 305978 295928
rect 3050 295264 3056 295316
rect 3108 295304 3114 295316
rect 56686 295304 56692 295316
rect 3108 295276 56692 295304
rect 3108 295264 3114 295276
rect 56686 295264 56692 295276
rect 56744 295264 56750 295316
rect 302786 293904 302792 293956
rect 302844 293944 302850 293956
rect 402238 293944 402244 293956
rect 302844 293916 402244 293944
rect 302844 293904 302850 293916
rect 402238 293904 402244 293916
rect 402296 293904 402302 293956
rect 302510 292476 302516 292528
rect 302568 292516 302574 292528
rect 320266 292516 320272 292528
rect 302568 292488 320272 292516
rect 302568 292476 302574 292488
rect 320266 292476 320272 292488
rect 320324 292476 320330 292528
rect 302694 289756 302700 289808
rect 302752 289796 302758 289808
rect 320174 289796 320180 289808
rect 302752 289768 320180 289796
rect 302752 289756 302758 289768
rect 320174 289756 320180 289768
rect 320232 289756 320238 289808
rect 302786 286968 302792 287020
rect 302844 287008 302850 287020
rect 318794 287008 318800 287020
rect 302844 286980 318800 287008
rect 302844 286968 302850 286980
rect 318794 286968 318800 286980
rect 318852 286968 318858 287020
rect 302694 285268 302700 285320
rect 302752 285308 302758 285320
rect 308398 285308 308404 285320
rect 302752 285280 308404 285308
rect 302752 285268 302758 285280
rect 308398 285268 308404 285280
rect 308456 285268 308462 285320
rect 302510 282820 302516 282872
rect 302568 282860 302574 282872
rect 450538 282860 450544 282872
rect 302568 282832 450544 282860
rect 302568 282820 302574 282832
rect 450538 282820 450544 282832
rect 450596 282820 450602 282872
rect 302510 281460 302516 281512
rect 302568 281500 302574 281512
rect 449158 281500 449164 281512
rect 302568 281472 449164 281500
rect 302568 281460 302574 281472
rect 449158 281460 449164 281472
rect 449216 281460 449222 281512
rect 3418 280100 3424 280152
rect 3476 280140 3482 280152
rect 35158 280140 35164 280152
rect 3476 280112 35164 280140
rect 3476 280100 3482 280112
rect 35158 280100 35164 280112
rect 35216 280100 35222 280152
rect 302326 278672 302332 278724
rect 302384 278712 302390 278724
rect 447778 278712 447784 278724
rect 302384 278684 447784 278712
rect 302384 278672 302390 278684
rect 447778 278672 447784 278684
rect 447836 278672 447842 278724
rect 302602 277312 302608 277364
rect 302660 277352 302666 277364
rect 446398 277352 446404 277364
rect 302660 277324 446404 277352
rect 302660 277312 302666 277324
rect 446398 277312 446404 277324
rect 446456 277312 446462 277364
rect 302786 274592 302792 274644
rect 302844 274632 302850 274644
rect 358814 274632 358820 274644
rect 302844 274604 358820 274632
rect 302844 274592 302850 274604
rect 358814 274592 358820 274604
rect 358872 274592 358878 274644
rect 302510 271804 302516 271856
rect 302568 271844 302574 271856
rect 357434 271844 357440 271856
rect 302568 271816 357440 271844
rect 302568 271804 302574 271816
rect 357434 271804 357440 271816
rect 357492 271804 357498 271856
rect 302510 270444 302516 270496
rect 302568 270484 302574 270496
rect 356054 270484 356060 270496
rect 302568 270456 356060 270484
rect 302568 270444 302574 270456
rect 356054 270444 356060 270456
rect 356112 270444 356118 270496
rect 302326 267656 302332 267708
rect 302384 267696 302390 267708
rect 354674 267696 354680 267708
rect 302384 267668 354680 267696
rect 302384 267656 302390 267668
rect 354674 267656 354680 267668
rect 354732 267656 354738 267708
rect 302602 266296 302608 266348
rect 302660 266336 302666 266348
rect 353294 266336 353300 266348
rect 302660 266308 353300 266336
rect 302660 266296 302666 266308
rect 353294 266296 353300 266308
rect 353352 266296 353358 266348
rect 2774 266228 2780 266280
rect 2832 266268 2838 266280
rect 5258 266268 5264 266280
rect 2832 266240 5264 266268
rect 2832 266228 2838 266240
rect 5258 266228 5264 266240
rect 5316 266228 5322 266280
rect 302786 263508 302792 263560
rect 302844 263548 302850 263560
rect 352006 263548 352012 263560
rect 302844 263520 352012 263548
rect 302844 263508 302850 263520
rect 352006 263508 352012 263520
rect 352064 263508 352070 263560
rect 302510 260788 302516 260840
rect 302568 260828 302574 260840
rect 351914 260828 351920 260840
rect 302568 260800 351920 260828
rect 302568 260788 302574 260800
rect 351914 260788 351920 260800
rect 351972 260788 351978 260840
rect 302418 259360 302424 259412
rect 302476 259400 302482 259412
rect 350534 259400 350540 259412
rect 302476 259372 350540 259400
rect 302476 259360 302482 259372
rect 350534 259360 350540 259372
rect 350592 259360 350598 259412
rect 302326 256640 302332 256692
rect 302384 256680 302390 256692
rect 349154 256680 349160 256692
rect 302384 256652 349160 256680
rect 302384 256640 302390 256652
rect 349154 256640 349160 256652
rect 349212 256640 349218 256692
rect 302510 255212 302516 255264
rect 302568 255252 302574 255264
rect 347774 255252 347780 255264
rect 302568 255224 347780 255252
rect 302568 255212 302574 255224
rect 347774 255212 347780 255224
rect 347832 255212 347838 255264
rect 3418 252492 3424 252544
rect 3476 252532 3482 252544
rect 57146 252532 57152 252544
rect 3476 252504 57152 252532
rect 3476 252492 3482 252504
rect 57146 252492 57152 252504
rect 57204 252492 57210 252544
rect 302786 252492 302792 252544
rect 302844 252532 302850 252544
rect 346394 252532 346400 252544
rect 302844 252504 346400 252532
rect 302844 252492 302850 252504
rect 346394 252492 346400 252504
rect 346452 252492 346458 252544
rect 302786 249704 302792 249756
rect 302844 249744 302850 249756
rect 345014 249744 345020 249756
rect 302844 249716 345020 249744
rect 302844 249704 302850 249716
rect 345014 249704 345020 249716
rect 345072 249704 345078 249756
rect 302418 248344 302424 248396
rect 302476 248384 302482 248396
rect 343726 248384 343732 248396
rect 302476 248356 343732 248384
rect 302476 248344 302482 248356
rect 343726 248344 343732 248356
rect 343784 248344 343790 248396
rect 302694 245556 302700 245608
rect 302752 245596 302758 245608
rect 343634 245596 343640 245608
rect 302752 245568 343640 245596
rect 302752 245556 302758 245568
rect 343634 245556 343640 245568
rect 343692 245556 343698 245608
rect 302510 244196 302516 244248
rect 302568 244236 302574 244248
rect 342254 244236 342260 244248
rect 302568 244208 342260 244236
rect 302568 244196 302574 244208
rect 342254 244196 342260 244208
rect 342312 244196 342318 244248
rect 302786 241408 302792 241460
rect 302844 241448 302850 241460
rect 340874 241448 340880 241460
rect 302844 241420 340880 241448
rect 302844 241408 302850 241420
rect 340874 241408 340880 241420
rect 340932 241408 340938 241460
rect 302786 238688 302792 238740
rect 302844 238728 302850 238740
rect 339494 238728 339500 238740
rect 302844 238700 339500 238728
rect 302844 238688 302850 238700
rect 339494 238688 339500 238700
rect 339552 238688 339558 238740
rect 3418 237328 3424 237380
rect 3476 237368 3482 237380
rect 37918 237368 37924 237380
rect 3476 237340 37924 237368
rect 3476 237328 3482 237340
rect 37918 237328 37924 237340
rect 37976 237328 37982 237380
rect 302418 237328 302424 237380
rect 302476 237368 302482 237380
rect 338114 237368 338120 237380
rect 302476 237340 338120 237368
rect 302476 237328 302482 237340
rect 338114 237328 338120 237340
rect 338172 237328 338178 237380
rect 302694 234540 302700 234592
rect 302752 234580 302758 234592
rect 336826 234580 336832 234592
rect 302752 234552 336832 234580
rect 302752 234540 302758 234552
rect 336826 234540 336832 234552
rect 336884 234540 336890 234592
rect 302510 233180 302516 233232
rect 302568 233220 302574 233232
rect 336734 233220 336740 233232
rect 302568 233192 336740 233220
rect 302568 233180 302574 233192
rect 336734 233180 336740 233192
rect 336792 233180 336798 233232
rect 302786 230392 302792 230444
rect 302844 230432 302850 230444
rect 335354 230432 335360 230444
rect 302844 230404 335360 230432
rect 302844 230392 302850 230404
rect 335354 230392 335360 230404
rect 335412 230392 335418 230444
rect 302786 227672 302792 227724
rect 302844 227712 302850 227724
rect 333974 227712 333980 227724
rect 302844 227684 333980 227712
rect 302844 227672 302850 227684
rect 333974 227672 333980 227684
rect 334032 227672 334038 227724
rect 302786 226244 302792 226296
rect 302844 226284 302850 226296
rect 332594 226284 332600 226296
rect 302844 226256 332600 226284
rect 302844 226244 302850 226256
rect 332594 226244 332600 226256
rect 332652 226244 332658 226296
rect 302694 223524 302700 223576
rect 302752 223564 302758 223576
rect 309778 223564 309784 223576
rect 302752 223536 309784 223564
rect 302752 223524 302758 223536
rect 309778 223524 309784 223536
rect 309836 223524 309842 223576
rect 2774 223048 2780 223100
rect 2832 223088 2838 223100
rect 5166 223088 5172 223100
rect 2832 223060 5172 223088
rect 2832 223048 2838 223060
rect 5166 223048 5172 223060
rect 5224 223048 5230 223100
rect 302786 222096 302792 222148
rect 302844 222136 302850 222148
rect 329926 222136 329932 222148
rect 302844 222108 329932 222136
rect 302844 222096 302850 222108
rect 329926 222096 329932 222108
rect 329984 222096 329990 222148
rect 302786 219376 302792 219428
rect 302844 219416 302850 219428
rect 312538 219416 312544 219428
rect 302844 219388 312544 219416
rect 302844 219376 302850 219388
rect 312538 219376 312544 219388
rect 312596 219376 312602 219428
rect 302786 216588 302792 216640
rect 302844 216628 302850 216640
rect 315298 216628 315304 216640
rect 302844 216600 315304 216628
rect 302844 216588 302850 216600
rect 315298 216588 315304 216600
rect 315356 216588 315362 216640
rect 302786 215228 302792 215280
rect 302844 215268 302850 215280
rect 327074 215268 327080 215280
rect 302844 215240 327080 215268
rect 302844 215228 302850 215240
rect 327074 215228 327080 215240
rect 327132 215228 327138 215280
rect 302602 212440 302608 212492
rect 302660 212480 302666 212492
rect 325694 212480 325700 212492
rect 302660 212452 325700 212480
rect 302660 212440 302666 212452
rect 325694 212440 325700 212452
rect 325752 212440 325758 212492
rect 302786 211080 302792 211132
rect 302844 211120 302850 211132
rect 316678 211120 316684 211132
rect 302844 211092 316684 211120
rect 302844 211080 302850 211092
rect 316678 211080 316684 211092
rect 316736 211080 316742 211132
rect 302786 208292 302792 208344
rect 302844 208332 302850 208344
rect 322934 208332 322940 208344
rect 302844 208304 322940 208332
rect 302844 208292 302850 208304
rect 322934 208292 322940 208304
rect 322992 208292 322998 208344
rect 302786 205572 302792 205624
rect 302844 205612 302850 205624
rect 321554 205612 321560 205624
rect 302844 205584 321560 205612
rect 302844 205572 302850 205584
rect 321554 205572 321560 205584
rect 321612 205572 321618 205624
rect 56962 205504 56968 205556
rect 57020 205544 57026 205556
rect 57020 205516 57192 205544
rect 57020 205504 57026 205516
rect 57164 205216 57192 205516
rect 579890 205368 579896 205420
rect 579948 205408 579954 205420
rect 580166 205408 580172 205420
rect 579948 205380 580172 205408
rect 579948 205368 579954 205380
rect 580166 205368 580172 205380
rect 580224 205368 580230 205420
rect 57146 205164 57152 205216
rect 57204 205164 57210 205216
rect 57146 201600 57152 201612
rect 57072 201572 57152 201600
rect 57072 201396 57100 201572
rect 57146 201560 57152 201572
rect 57204 201560 57210 201612
rect 57514 201600 57520 201612
rect 57440 201572 57520 201600
rect 57146 201424 57152 201476
rect 57204 201464 57210 201476
rect 57440 201464 57468 201572
rect 57514 201560 57520 201572
rect 57572 201560 57578 201612
rect 57204 201436 57468 201464
rect 57204 201424 57210 201436
rect 57514 201424 57520 201476
rect 57572 201464 57578 201476
rect 57790 201464 57796 201476
rect 57572 201436 57796 201464
rect 57572 201424 57578 201436
rect 57790 201424 57796 201436
rect 57848 201424 57854 201476
rect 57974 201396 57980 201408
rect 57072 201368 57980 201396
rect 57974 201356 57980 201368
rect 58032 201356 58038 201408
rect 57054 200812 57060 200864
rect 57112 200852 57118 200864
rect 580810 200852 580816 200864
rect 57112 200824 580816 200852
rect 57112 200812 57118 200824
rect 580810 200812 580816 200824
rect 580868 200812 580874 200864
rect 56962 200744 56968 200796
rect 57020 200784 57026 200796
rect 579982 200784 579988 200796
rect 57020 200756 579988 200784
rect 57020 200744 57026 200756
rect 579982 200744 579988 200756
rect 580040 200744 580046 200796
rect 57698 200676 57704 200728
rect 57756 200716 57762 200728
rect 580534 200716 580540 200728
rect 57756 200688 580540 200716
rect 57756 200676 57762 200688
rect 580534 200676 580540 200688
rect 580592 200676 580598 200728
rect 57146 200608 57152 200660
rect 57204 200648 57210 200660
rect 580166 200648 580172 200660
rect 57204 200620 580172 200648
rect 57204 200608 57210 200620
rect 580166 200608 580172 200620
rect 580224 200608 580230 200660
rect 57514 200540 57520 200592
rect 57572 200580 57578 200592
rect 580074 200580 580080 200592
rect 57572 200552 580080 200580
rect 57572 200540 57578 200552
rect 580074 200540 580080 200552
rect 580132 200540 580138 200592
rect 57974 200472 57980 200524
rect 58032 200512 58038 200524
rect 579890 200512 579896 200524
rect 58032 200484 579896 200512
rect 58032 200472 58038 200484
rect 579890 200472 579896 200484
rect 579948 200472 579954 200524
rect 59814 200404 59820 200456
rect 59872 200444 59878 200456
rect 580350 200444 580356 200456
rect 59872 200416 580356 200444
rect 59872 200404 59878 200416
rect 580350 200404 580356 200416
rect 580408 200404 580414 200456
rect 57238 200064 57244 200116
rect 57296 200104 57302 200116
rect 580718 200104 580724 200116
rect 57296 200076 580724 200104
rect 57296 200064 57302 200076
rect 580718 200064 580724 200076
rect 580776 200064 580782 200116
rect 57606 199996 57612 200048
rect 57664 200036 57670 200048
rect 580902 200036 580908 200048
rect 57664 200008 580908 200036
rect 57664 199996 57670 200008
rect 580902 199996 580908 200008
rect 580960 199996 580966 200048
rect 56870 199928 56876 199980
rect 56928 199968 56934 199980
rect 580626 199968 580632 199980
rect 56928 199940 580632 199968
rect 56928 199928 56934 199940
rect 580626 199928 580632 199940
rect 580684 199928 580690 199980
rect 57882 199860 57888 199912
rect 57940 199900 57946 199912
rect 580442 199900 580448 199912
rect 57940 199872 580448 199900
rect 57940 199860 57946 199872
rect 580442 199860 580448 199872
rect 580500 199860 580506 199912
rect 71682 198636 71688 198688
rect 71740 198676 71746 198688
rect 186314 198676 186320 198688
rect 71740 198648 186320 198676
rect 71740 198636 71746 198648
rect 186314 198636 186320 198648
rect 186372 198636 186378 198688
rect 79962 198568 79968 198620
rect 80020 198608 80026 198620
rect 201126 198608 201132 198620
rect 80020 198580 201132 198608
rect 80020 198568 80026 198580
rect 201126 198568 201132 198580
rect 201184 198568 201190 198620
rect 78582 198500 78588 198552
rect 78640 198540 78646 198552
rect 199010 198540 199016 198552
rect 78640 198512 199016 198540
rect 78640 198500 78646 198512
rect 199010 198500 199016 198512
rect 199068 198500 199074 198552
rect 32398 198432 32404 198484
rect 32456 198472 32462 198484
rect 69474 198472 69480 198484
rect 32456 198444 69480 198472
rect 32456 198432 32462 198444
rect 69474 198432 69480 198444
rect 69532 198432 69538 198484
rect 85482 198432 85488 198484
rect 85540 198472 85546 198484
rect 211798 198472 211804 198484
rect 85540 198444 211804 198472
rect 85540 198432 85546 198444
rect 211798 198432 211804 198444
rect 211856 198432 211862 198484
rect 10962 198364 10968 198416
rect 11020 198404 11026 198416
rect 77938 198404 77944 198416
rect 11020 198376 77944 198404
rect 11020 198364 11026 198376
rect 77938 198364 77944 198376
rect 77996 198364 78002 198416
rect 86862 198364 86868 198416
rect 86920 198404 86926 198416
rect 213914 198404 213920 198416
rect 86920 198376 213920 198404
rect 86920 198364 86926 198376
rect 213914 198364 213920 198376
rect 213972 198364 213978 198416
rect 12342 198296 12348 198348
rect 12400 198336 12406 198348
rect 80054 198336 80060 198348
rect 12400 198308 80060 198336
rect 12400 198296 12406 198308
rect 80054 198296 80060 198308
rect 80112 198296 80118 198348
rect 92382 198296 92388 198348
rect 92440 198336 92446 198348
rect 224494 198336 224500 198348
rect 92440 198308 224500 198336
rect 92440 198296 92446 198308
rect 224494 198296 224500 198308
rect 224552 198296 224558 198348
rect 15102 198228 15108 198280
rect 15160 198268 15166 198280
rect 86494 198268 86500 198280
rect 15160 198240 86500 198268
rect 15160 198228 15166 198240
rect 86494 198228 86500 198240
rect 86552 198228 86558 198280
rect 93762 198228 93768 198280
rect 93820 198268 93826 198280
rect 226610 198268 226616 198280
rect 93820 198240 226616 198268
rect 93820 198228 93826 198240
rect 226610 198228 226616 198240
rect 226668 198228 226674 198280
rect 16482 198160 16488 198212
rect 16540 198200 16546 198212
rect 88610 198200 88616 198212
rect 16540 198172 88616 198200
rect 16540 198160 16546 198172
rect 88610 198160 88616 198172
rect 88668 198160 88674 198212
rect 99190 198160 99196 198212
rect 99248 198200 99254 198212
rect 237282 198200 237288 198212
rect 99248 198172 237288 198200
rect 99248 198160 99254 198172
rect 237282 198160 237288 198172
rect 237340 198160 237346 198212
rect 20622 198092 20628 198144
rect 20680 198132 20686 198144
rect 94958 198132 94964 198144
rect 20680 198104 94964 198132
rect 20680 198092 20686 198104
rect 94958 198092 94964 198104
rect 95016 198092 95022 198144
rect 100662 198092 100668 198144
rect 100720 198132 100726 198144
rect 239398 198132 239404 198144
rect 100720 198104 239404 198132
rect 100720 198092 100726 198104
rect 239398 198092 239404 198104
rect 239456 198092 239462 198144
rect 21910 198024 21916 198076
rect 21968 198064 21974 198076
rect 97074 198064 97080 198076
rect 21968 198036 97080 198064
rect 21968 198024 21974 198036
rect 97074 198024 97080 198036
rect 97132 198024 97138 198076
rect 107562 198024 107568 198076
rect 107620 198064 107626 198076
rect 249978 198064 249984 198076
rect 107620 198036 249984 198064
rect 107620 198024 107626 198036
rect 249978 198024 249984 198036
rect 250036 198024 250042 198076
rect 26142 197956 26148 198008
rect 26200 197996 26206 198008
rect 105538 197996 105544 198008
rect 26200 197968 105544 197996
rect 26200 197956 26206 197968
rect 105538 197956 105544 197968
rect 105596 197956 105602 198008
rect 107470 197956 107476 198008
rect 107528 197996 107534 198008
rect 252094 197996 252100 198008
rect 107528 197968 252100 197996
rect 107528 197956 107534 197968
rect 252094 197956 252100 197968
rect 252152 197956 252158 198008
rect 72970 197888 72976 197940
rect 73028 197928 73034 197940
rect 188430 197928 188436 197940
rect 73028 197900 188436 197928
rect 73028 197888 73034 197900
rect 188430 197888 188436 197900
rect 188488 197888 188494 197940
rect 64782 197820 64788 197872
rect 64840 197860 64846 197872
rect 175642 197860 175648 197872
rect 64840 197832 175648 197860
rect 64840 197820 64846 197832
rect 175642 197820 175648 197832
rect 175700 197820 175706 197872
rect 57882 197752 57888 197804
rect 57940 197792 57946 197804
rect 162946 197792 162952 197804
rect 57940 197764 162952 197792
rect 57940 197752 57946 197764
rect 162946 197752 162952 197764
rect 163004 197752 163010 197804
rect 55122 197684 55128 197736
rect 55180 197724 55186 197736
rect 156506 197724 156512 197736
rect 55180 197696 156512 197724
rect 55180 197684 55186 197696
rect 156506 197684 156512 197696
rect 156564 197684 156570 197736
rect 50982 197616 50988 197668
rect 51040 197656 51046 197668
rect 150158 197656 150164 197668
rect 51040 197628 150164 197656
rect 51040 197616 51046 197628
rect 150158 197616 150164 197628
rect 150216 197616 150222 197668
rect 48130 197548 48136 197600
rect 48188 197588 48194 197600
rect 143810 197588 143816 197600
rect 48188 197560 143816 197588
rect 48188 197548 48194 197560
rect 143810 197548 143816 197560
rect 143868 197548 143874 197600
rect 42702 197480 42708 197532
rect 42760 197520 42766 197532
rect 135346 197520 135352 197532
rect 42760 197492 135352 197520
rect 42760 197480 42766 197492
rect 135346 197480 135352 197492
rect 135404 197480 135410 197532
rect 39942 197412 39948 197464
rect 40000 197452 40006 197464
rect 130286 197452 130292 197464
rect 40000 197424 130292 197452
rect 40000 197412 40006 197424
rect 130286 197412 130292 197424
rect 130344 197412 130350 197464
rect 130378 197412 130384 197464
rect 130436 197452 130442 197464
rect 148042 197452 148048 197464
rect 130436 197424 148048 197452
rect 130436 197412 130442 197424
rect 148042 197412 148048 197424
rect 148100 197412 148106 197464
rect 127618 197344 127624 197396
rect 127676 197384 127682 197396
rect 160830 197384 160836 197396
rect 127676 197356 160836 197384
rect 127676 197344 127682 197356
rect 160830 197344 160836 197356
rect 160888 197344 160894 197396
rect 3142 194488 3148 194540
rect 3200 194528 3206 194540
rect 53098 194528 53104 194540
rect 3200 194500 53104 194528
rect 3200 194488 3206 194500
rect 53098 194488 53104 194500
rect 53156 194488 53162 194540
rect 92198 183540 92204 183592
rect 92256 183580 92262 183592
rect 92382 183580 92388 183592
rect 92256 183552 92388 183580
rect 92256 183540 92262 183552
rect 92382 183540 92388 183552
rect 92440 183540 92446 183592
rect 57330 182112 57336 182164
rect 57388 182152 57394 182164
rect 580166 182152 580172 182164
rect 57388 182124 580172 182152
rect 57388 182112 57394 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 31018 180792 31024 180804
rect 3292 180764 31024 180792
rect 3292 180752 3298 180764
rect 31018 180752 31024 180764
rect 31076 180752 31082 180804
rect 57422 171028 57428 171080
rect 57480 171068 57486 171080
rect 580166 171068 580172 171080
rect 57480 171040 580172 171068
rect 57480 171028 57486 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 2774 165452 2780 165504
rect 2832 165492 2838 165504
rect 5074 165492 5080 165504
rect 2832 165464 5080 165492
rect 2832 165452 2838 165464
rect 5074 165452 5080 165464
rect 5132 165452 5138 165504
rect 56778 158652 56784 158704
rect 56836 158692 56842 158704
rect 579798 158692 579804 158704
rect 56836 158664 579804 158692
rect 56836 158652 56842 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 92198 154504 92204 154556
rect 92256 154544 92262 154556
rect 92382 154544 92388 154556
rect 92256 154516 92388 154544
rect 92256 154504 92262 154516
rect 92382 154504 92388 154516
rect 92440 154504 92446 154556
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 19978 151756 19984 151768
rect 3200 151728 19984 151756
rect 3200 151716 3206 151728
rect 19978 151716 19984 151728
rect 20036 151716 20042 151768
rect 3234 136552 3240 136604
rect 3292 136592 3298 136604
rect 33778 136592 33784 136604
rect 3292 136564 33784 136592
rect 3292 136552 3298 136564
rect 33778 136552 33784 136564
rect 33836 136552 33842 136604
rect 56594 135192 56600 135244
rect 56652 135232 56658 135244
rect 580166 135232 580172 135244
rect 56652 135204 580172 135232
rect 56652 135192 56658 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 92106 135124 92112 135176
rect 92164 135164 92170 135176
rect 92382 135164 92388 135176
rect 92164 135136 92388 135164
rect 92164 135124 92170 135136
rect 92382 135124 92388 135136
rect 92440 135124 92446 135176
rect 56686 124108 56692 124160
rect 56744 124148 56750 124160
rect 580166 124148 580172 124160
rect 56744 124120 580172 124148
rect 56744 124108 56750 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 2774 122340 2780 122392
rect 2832 122380 2838 122392
rect 4890 122380 4896 122392
rect 2832 122352 4896 122380
rect 2832 122340 2838 122352
rect 4890 122340 4896 122352
rect 4948 122340 4954 122392
rect 92198 115880 92204 115932
rect 92256 115920 92262 115932
rect 92382 115920 92388 115932
rect 92256 115892 92388 115920
rect 92256 115880 92262 115892
rect 92382 115880 92388 115892
rect 92440 115880 92446 115932
rect 89622 110780 89628 110832
rect 89680 110820 89686 110832
rect 96522 110820 96528 110832
rect 89680 110792 96528 110820
rect 89680 110780 89686 110792
rect 96522 110780 96528 110792
rect 96580 110780 96586 110832
rect 147582 110644 147588 110696
rect 147640 110684 147646 110696
rect 154482 110684 154488 110696
rect 147640 110656 154488 110684
rect 147640 110644 147646 110656
rect 154482 110644 154488 110656
rect 154540 110644 154546 110696
rect 116026 110508 116032 110560
rect 116084 110548 116090 110560
rect 118786 110548 118792 110560
rect 116084 110520 118792 110548
rect 116084 110508 116090 110520
rect 118786 110508 118792 110520
rect 118844 110508 118850 110560
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 17218 108984 17224 108996
rect 3292 108956 17224 108984
rect 3292 108944 3298 108956
rect 17218 108944 17224 108956
rect 17276 108944 17282 108996
rect 92198 106292 92204 106344
rect 92256 106332 92262 106344
rect 92382 106332 92388 106344
rect 92256 106304 92388 106332
rect 92256 106292 92262 106304
rect 92382 106292 92388 106304
rect 92440 106292 92446 106344
rect 92382 96568 92388 96620
rect 92440 96608 92446 96620
rect 92566 96608 92572 96620
rect 92440 96580 92572 96608
rect 92440 96568 92446 96580
rect 92566 96568 92572 96580
rect 92624 96568 92630 96620
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 43438 93820 43444 93832
rect 3476 93792 43444 93820
rect 3476 93780 3482 93792
rect 43438 93780 43444 93792
rect 43496 93780 43502 93832
rect 89622 87252 89628 87304
rect 89680 87292 89686 87304
rect 96522 87292 96528 87304
rect 89680 87264 96528 87292
rect 89680 87252 89686 87264
rect 96522 87252 96528 87264
rect 96580 87252 96586 87304
rect 145558 87116 145564 87168
rect 145616 87156 145622 87168
rect 154482 87156 154488 87168
rect 145616 87128 154488 87156
rect 145616 87116 145622 87128
rect 154482 87116 154488 87128
rect 154540 87116 154546 87168
rect 92382 86980 92388 87032
rect 92440 87020 92446 87032
rect 92566 87020 92572 87032
rect 92440 86992 92572 87020
rect 92440 86980 92446 86992
rect 92566 86980 92572 86992
rect 92624 86980 92630 87032
rect 116026 86980 116032 87032
rect 116084 87020 116090 87032
rect 120810 87020 120816 87032
rect 116084 86992 120816 87020
rect 116084 86980 116090 86992
rect 120810 86980 120816 86992
rect 120868 86980 120874 87032
rect 3418 79976 3424 80028
rect 3476 80016 3482 80028
rect 10318 80016 10324 80028
rect 3476 79988 10324 80016
rect 3476 79976 3482 79988
rect 10318 79976 10324 79988
rect 10376 79976 10382 80028
rect 89622 76236 89628 76288
rect 89680 76276 89686 76288
rect 96522 76276 96528 76288
rect 89680 76248 96528 76276
rect 89680 76236 89686 76248
rect 96522 76236 96528 76248
rect 96580 76236 96586 76288
rect 147582 76100 147588 76152
rect 147640 76140 147646 76152
rect 154482 76140 154488 76152
rect 147640 76112 154488 76140
rect 147640 76100 147646 76112
rect 154482 76100 154488 76112
rect 154540 76100 154546 76152
rect 116026 75964 116032 76016
rect 116084 76004 116090 76016
rect 118786 76004 118792 76016
rect 116084 75976 118792 76004
rect 116084 75964 116090 75976
rect 118786 75964 118792 75976
rect 118844 75964 118850 76016
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 39298 64852 39304 64864
rect 3384 64824 39304 64852
rect 3384 64812 3390 64824
rect 39298 64812 39304 64824
rect 39356 64812 39362 64864
rect 88886 63860 88892 63912
rect 88944 63900 88950 63912
rect 96522 63900 96528 63912
rect 88944 63872 96528 63900
rect 88944 63860 88950 63872
rect 96522 63860 96528 63872
rect 96580 63860 96586 63912
rect 147582 63724 147588 63776
rect 147640 63764 147646 63776
rect 154482 63764 154488 63776
rect 147640 63736 154488 63764
rect 147640 63724 147646 63736
rect 154482 63724 154488 63736
rect 154540 63724 154546 63776
rect 116026 63588 116032 63640
rect 116084 63628 116090 63640
rect 118786 63628 118792 63640
rect 116084 63600 118792 63628
rect 116084 63588 116090 63600
rect 118786 63588 118792 63600
rect 118844 63588 118850 63640
rect 92198 57876 92204 57928
rect 92256 57916 92262 57928
rect 92382 57916 92388 57928
rect 92256 57888 92388 57916
rect 92256 57876 92262 57888
rect 92382 57876 92388 57888
rect 92440 57876 92446 57928
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 46198 51048 46204 51060
rect 3476 51020 46204 51048
rect 3476 51008 3482 51020
rect 46198 51008 46204 51020
rect 46256 51008 46262 51060
rect 92198 48288 92204 48340
rect 92256 48328 92262 48340
rect 92382 48328 92388 48340
rect 92256 48300 92388 48328
rect 92256 48288 92262 48300
rect 92382 48288 92388 48300
rect 92440 48288 92446 48340
rect 88886 40332 88892 40384
rect 88944 40372 88950 40384
rect 96522 40372 96528 40384
rect 88944 40344 96528 40372
rect 88944 40332 88950 40344
rect 96522 40332 96528 40344
rect 96580 40332 96586 40384
rect 147582 40196 147588 40248
rect 147640 40236 147646 40248
rect 154482 40236 154488 40248
rect 147640 40208 154488 40236
rect 147640 40196 147646 40208
rect 154482 40196 154488 40208
rect 154540 40196 154546 40248
rect 116026 40060 116032 40112
rect 116084 40100 116090 40112
rect 118786 40100 118792 40112
rect 116084 40072 118792 40100
rect 116084 40060 116090 40072
rect 118786 40060 118792 40072
rect 118844 40060 118850 40112
rect 92198 38564 92204 38616
rect 92256 38604 92262 38616
rect 92382 38604 92388 38616
rect 92256 38576 92388 38604
rect 92256 38564 92262 38576
rect 92382 38564 92388 38576
rect 92440 38564 92446 38616
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 15838 35884 15844 35896
rect 3476 35856 15844 35884
rect 3476 35844 3482 35856
rect 15838 35844 15844 35856
rect 15896 35844 15902 35896
rect 89622 29316 89628 29368
rect 89680 29356 89686 29368
rect 96522 29356 96528 29368
rect 89680 29328 96528 29356
rect 89680 29316 89686 29328
rect 96522 29316 96528 29328
rect 96580 29316 96586 29368
rect 116026 29044 116032 29096
rect 116084 29084 116090 29096
rect 120810 29084 120816 29096
rect 116084 29056 120816 29084
rect 116084 29044 116090 29056
rect 120810 29044 120816 29056
rect 120868 29044 120874 29096
rect 145006 29044 145012 29096
rect 145064 29084 145070 29096
rect 154482 29084 154488 29096
rect 145064 29056 154488 29084
rect 145064 29044 145070 29056
rect 154482 29044 154488 29056
rect 154540 29044 154546 29096
rect 92198 28976 92204 29028
rect 92256 29016 92262 29028
rect 92382 29016 92388 29028
rect 92256 28988 92388 29016
rect 92256 28976 92262 28988
rect 92382 28976 92388 28988
rect 92440 28976 92446 29028
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 48958 22080 48964 22092
rect 3200 22052 48964 22080
rect 3200 22040 3206 22052
rect 48958 22040 48964 22052
rect 49016 22040 49022 22092
rect 92198 19252 92204 19304
rect 92256 19292 92262 19304
rect 92382 19292 92388 19304
rect 92256 19264 92388 19292
rect 92256 19252 92262 19264
rect 92382 19252 92388 19264
rect 92440 19252 92446 19304
rect 57790 17892 57796 17944
rect 57848 17932 57854 17944
rect 579798 17932 579804 17944
rect 57848 17904 579804 17932
rect 57848 17892 57854 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 92198 9664 92204 9716
rect 92256 9704 92262 9716
rect 92382 9704 92388 9716
rect 92256 9676 92388 9704
rect 92256 9664 92262 9676
rect 92382 9664 92388 9676
rect 92440 9664 92446 9716
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 51718 8276 51724 8288
rect 3476 8248 51724 8276
rect 3476 8236 3482 8248
rect 51718 8236 51724 8248
rect 51776 8236 51782 8288
rect 52822 6672 52828 6724
rect 52880 6712 52886 6724
rect 153194 6712 153200 6724
rect 52880 6684 153200 6712
rect 52880 6672 52886 6684
rect 153194 6672 153200 6684
rect 153252 6672 153258 6724
rect 59998 6604 60004 6656
rect 60056 6644 60062 6656
rect 166994 6644 167000 6656
rect 60056 6616 167000 6644
rect 60056 6604 60062 6616
rect 166994 6604 167000 6616
rect 167052 6604 167058 6656
rect 63586 6536 63592 6588
rect 63644 6576 63650 6588
rect 172514 6576 172520 6588
rect 63644 6548 172520 6576
rect 63644 6536 63650 6548
rect 172514 6536 172520 6548
rect 172572 6536 172578 6588
rect 101582 6468 101588 6520
rect 101640 6508 101646 6520
rect 241514 6508 241520 6520
rect 101640 6480 241520 6508
rect 101640 6468 101646 6480
rect 241514 6468 241520 6480
rect 241572 6468 241578 6520
rect 108758 6400 108764 6452
rect 108816 6440 108822 6452
rect 253934 6440 253940 6452
rect 108816 6412 253940 6440
rect 108816 6400 108822 6412
rect 253934 6400 253940 6412
rect 253992 6400 253998 6452
rect 112346 6332 112352 6384
rect 112404 6372 112410 6384
rect 259454 6372 259460 6384
rect 112404 6344 259460 6372
rect 112404 6332 112410 6344
rect 259454 6332 259460 6344
rect 259512 6332 259518 6384
rect 116118 6264 116124 6316
rect 116176 6304 116182 6316
rect 266354 6304 266360 6316
rect 116176 6276 266360 6304
rect 116176 6264 116182 6276
rect 266354 6264 266360 6276
rect 266412 6264 266418 6316
rect 119430 6196 119436 6248
rect 119488 6236 119494 6248
rect 273254 6236 273260 6248
rect 119488 6208 273260 6236
rect 119488 6196 119494 6208
rect 273254 6196 273260 6208
rect 273312 6196 273318 6248
rect 123018 6128 123024 6180
rect 123076 6168 123082 6180
rect 278774 6168 278780 6180
rect 123076 6140 278780 6168
rect 123076 6128 123082 6140
rect 278774 6128 278780 6140
rect 278832 6128 278838 6180
rect 80054 5556 80060 5568
rect 76576 5528 80060 5556
rect 65518 5448 65524 5500
rect 65576 5488 65582 5500
rect 76576 5488 76604 5528
rect 80054 5516 80060 5528
rect 80112 5516 80118 5568
rect 103974 5516 103980 5568
rect 104032 5556 104038 5568
rect 109402 5556 109408 5568
rect 104032 5528 109408 5556
rect 104032 5516 104038 5528
rect 109402 5516 109408 5528
rect 109460 5516 109466 5568
rect 65576 5460 76604 5488
rect 65576 5448 65582 5460
rect 76650 5448 76656 5500
rect 76708 5488 76714 5500
rect 195974 5488 195980 5500
rect 76708 5460 195980 5488
rect 76708 5448 76714 5460
rect 195974 5448 195980 5460
rect 196032 5448 196038 5500
rect 12434 5380 12440 5432
rect 12492 5420 12498 5432
rect 81434 5420 81440 5432
rect 12492 5392 81440 5420
rect 12492 5380 12498 5392
rect 81434 5380 81440 5392
rect 81492 5380 81498 5432
rect 83826 5380 83832 5432
rect 83884 5420 83890 5432
rect 208394 5420 208400 5432
rect 83884 5392 208400 5420
rect 83884 5380 83890 5392
rect 208394 5380 208400 5392
rect 208452 5380 208458 5432
rect 80054 5312 80060 5364
rect 80112 5352 80118 5364
rect 80112 5324 91140 5352
rect 80112 5312 80118 5324
rect 17218 5244 17224 5296
rect 17276 5284 17282 5296
rect 89714 5284 89720 5296
rect 17276 5256 89720 5284
rect 17276 5244 17282 5256
rect 89714 5244 89720 5256
rect 89772 5244 89778 5296
rect 91112 5284 91140 5324
rect 91186 5312 91192 5364
rect 91244 5352 91250 5364
rect 222194 5352 222200 5364
rect 91244 5324 222200 5352
rect 91244 5312 91250 5324
rect 222194 5312 222200 5324
rect 222252 5312 222258 5364
rect 103974 5284 103980 5296
rect 91112 5256 103980 5284
rect 103974 5244 103980 5256
rect 104032 5244 104038 5296
rect 104250 5244 104256 5296
rect 104308 5284 104314 5296
rect 104308 5256 106412 5284
rect 104308 5244 104314 5256
rect 22002 5176 22008 5228
rect 22060 5216 22066 5228
rect 97994 5216 98000 5228
rect 22060 5188 98000 5216
rect 22060 5176 22066 5188
rect 97994 5176 98000 5188
rect 98052 5176 98058 5228
rect 98822 5176 98828 5228
rect 98880 5216 98886 5228
rect 106384 5216 106412 5256
rect 106458 5244 106464 5296
rect 106516 5284 106522 5296
rect 234614 5284 234620 5296
rect 106516 5256 234620 5284
rect 106516 5244 106522 5256
rect 234614 5244 234620 5256
rect 234672 5244 234678 5296
rect 107654 5216 107660 5228
rect 98880 5188 106320 5216
rect 106384 5188 107660 5216
rect 98880 5176 98886 5188
rect 106292 5160 106320 5188
rect 107654 5176 107660 5188
rect 107712 5176 107718 5228
rect 126606 5176 126612 5228
rect 126664 5216 126670 5228
rect 285674 5216 285680 5228
rect 126664 5188 285680 5216
rect 126664 5176 126670 5188
rect 285674 5176 285680 5188
rect 285732 5176 285738 5228
rect 26694 5108 26700 5160
rect 26752 5148 26758 5160
rect 104066 5148 104072 5160
rect 26752 5120 104072 5148
rect 26752 5108 26758 5120
rect 104066 5108 104072 5120
rect 104124 5108 104130 5160
rect 106274 5108 106280 5160
rect 106332 5108 106338 5160
rect 109402 5108 109408 5160
rect 109460 5148 109466 5160
rect 118602 5148 118608 5160
rect 109460 5120 118608 5148
rect 109460 5108 109466 5120
rect 118602 5108 118608 5120
rect 118660 5108 118666 5160
rect 127802 5108 127808 5160
rect 127860 5148 127866 5160
rect 287054 5148 287060 5160
rect 127860 5120 287060 5148
rect 127860 5108 127866 5120
rect 287054 5108 287060 5120
rect 287112 5108 287118 5160
rect 49326 5040 49332 5092
rect 49384 5080 49390 5092
rect 118510 5080 118516 5092
rect 49384 5052 118516 5080
rect 49384 5040 49390 5052
rect 118510 5040 118516 5052
rect 118568 5040 118574 5092
rect 118786 5040 118792 5092
rect 118844 5080 118850 5092
rect 130378 5080 130384 5092
rect 118844 5052 130384 5080
rect 118844 5040 118850 5052
rect 130378 5040 130384 5052
rect 130436 5040 130442 5092
rect 291194 5080 291200 5092
rect 130488 5052 291200 5080
rect 30282 4972 30288 5024
rect 30340 5012 30346 5024
rect 113174 5012 113180 5024
rect 30340 4984 113180 5012
rect 30340 4972 30346 4984
rect 113174 4972 113180 4984
rect 113232 4972 113238 5024
rect 114738 4972 114744 5024
rect 114796 5012 114802 5024
rect 115842 5012 115848 5024
rect 114796 4984 115848 5012
rect 114796 4972 114802 4984
rect 115842 4972 115848 4984
rect 115900 4972 115906 5024
rect 118878 4972 118884 5024
rect 118936 5012 118942 5024
rect 127618 5012 127624 5024
rect 118936 4984 127624 5012
rect 118936 4972 118942 4984
rect 127618 4972 127624 4984
rect 127676 4972 127682 5024
rect 130194 4972 130200 5024
rect 130252 5012 130258 5024
rect 130488 5012 130516 5052
rect 291194 5040 291200 5052
rect 291252 5040 291258 5092
rect 289814 5012 289820 5024
rect 130252 4984 130516 5012
rect 130580 4984 289820 5012
rect 130252 4972 130258 4984
rect 33870 4904 33876 4956
rect 33928 4944 33934 4956
rect 120074 4944 120080 4956
rect 33928 4916 120080 4944
rect 33928 4904 33934 4916
rect 120074 4904 120080 4916
rect 120132 4904 120138 4956
rect 128998 4904 129004 4956
rect 129056 4944 129062 4956
rect 130580 4944 130608 4984
rect 289814 4972 289820 4984
rect 289872 4972 289878 5024
rect 129056 4916 130608 4944
rect 129056 4904 129062 4916
rect 131390 4904 131396 4956
rect 131448 4944 131454 4956
rect 293954 4944 293960 4956
rect 131448 4916 293960 4944
rect 131448 4904 131454 4916
rect 293954 4904 293960 4916
rect 294012 4904 294018 4956
rect 37366 4836 37372 4888
rect 37424 4876 37430 4888
rect 125594 4876 125600 4888
rect 37424 4848 125600 4876
rect 37424 4836 37430 4848
rect 125594 4836 125600 4848
rect 125652 4836 125658 4888
rect 134886 4836 134892 4888
rect 134944 4876 134950 4888
rect 298094 4876 298100 4888
rect 134944 4848 298100 4876
rect 134944 4836 134950 4848
rect 298094 4836 298100 4848
rect 298152 4836 298158 4888
rect 40954 4768 40960 4820
rect 41012 4808 41018 4820
rect 132494 4808 132500 4820
rect 41012 4780 132500 4808
rect 41012 4768 41018 4780
rect 132494 4768 132500 4780
rect 132552 4768 132558 4820
rect 132586 4768 132592 4820
rect 132644 4808 132650 4820
rect 296714 4808 296720 4820
rect 132644 4780 296720 4808
rect 132644 4768 132650 4780
rect 296714 4768 296720 4780
rect 296772 4768 296778 4820
rect 56410 4700 56416 4752
rect 56468 4740 56474 4752
rect 65518 4740 65524 4752
rect 56468 4712 65524 4740
rect 56468 4700 56474 4712
rect 65518 4700 65524 4712
rect 65576 4700 65582 4752
rect 73062 4700 73068 4752
rect 73120 4740 73126 4752
rect 190454 4740 190460 4752
rect 73120 4712 190460 4740
rect 73120 4700 73126 4712
rect 190454 4700 190460 4712
rect 190512 4700 190518 4752
rect 69474 4632 69480 4684
rect 69532 4672 69538 4684
rect 183554 4672 183560 4684
rect 69532 4644 183560 4672
rect 69532 4632 69538 4644
rect 183554 4632 183560 4644
rect 183612 4632 183618 4684
rect 65978 4564 65984 4616
rect 66036 4604 66042 4616
rect 176654 4604 176660 4616
rect 66036 4576 176660 4604
rect 66036 4564 66042 4576
rect 176654 4564 176660 4576
rect 176712 4564 176718 4616
rect 62390 4496 62396 4548
rect 62448 4536 62454 4548
rect 171134 4536 171140 4548
rect 62448 4508 171140 4536
rect 62448 4496 62454 4508
rect 171134 4496 171140 4508
rect 171192 4496 171198 4548
rect 58802 4428 58808 4480
rect 58860 4468 58866 4480
rect 164234 4468 164240 4480
rect 58860 4440 164240 4468
rect 58860 4428 58866 4440
rect 164234 4428 164240 4440
rect 164292 4428 164298 4480
rect 55214 4360 55220 4412
rect 55272 4400 55278 4412
rect 158714 4400 158720 4412
rect 55272 4372 158720 4400
rect 55272 4360 55278 4372
rect 158714 4360 158720 4372
rect 158772 4360 158778 4412
rect 51626 4292 51632 4344
rect 51684 4332 51690 4344
rect 151814 4332 151820 4344
rect 51684 4304 151820 4332
rect 51684 4292 51690 4304
rect 151814 4292 151820 4304
rect 151872 4292 151878 4344
rect 48222 4224 48228 4276
rect 48280 4264 48286 4276
rect 144914 4264 144920 4276
rect 48280 4236 144920 4264
rect 48280 4224 48286 4236
rect 144914 4224 144920 4236
rect 144972 4224 144978 4276
rect 44542 4156 44548 4208
rect 44600 4196 44606 4208
rect 139394 4196 139400 4208
rect 44600 4168 139400 4196
rect 44600 4156 44606 4168
rect 139394 4156 139400 4168
rect 139452 4156 139458 4208
rect 8846 4088 8852 4140
rect 8904 4128 8910 4140
rect 65610 4128 65616 4140
rect 8904 4100 65616 4128
rect 8904 4088 8910 4100
rect 65610 4088 65616 4100
rect 65668 4088 65674 4140
rect 84194 4128 84200 4140
rect 79336 4100 84200 4128
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 79336 4060 79364 4100
rect 84194 4088 84200 4100
rect 84252 4088 84258 4140
rect 84930 4088 84936 4140
rect 84988 4128 84994 4140
rect 85482 4128 85488 4140
rect 84988 4100 85488 4128
rect 84988 4088 84994 4100
rect 85482 4088 85488 4100
rect 85540 4088 85546 4140
rect 86126 4088 86132 4140
rect 86184 4128 86190 4140
rect 86862 4128 86868 4140
rect 86184 4100 86868 4128
rect 86184 4088 86190 4100
rect 86862 4088 86868 4100
rect 86920 4088 86926 4140
rect 86954 4088 86960 4140
rect 87012 4128 87018 4140
rect 207014 4128 207020 4140
rect 87012 4100 207020 4128
rect 87012 4088 87018 4100
rect 207014 4088 207020 4100
rect 207072 4088 207078 4140
rect 92474 4060 92480 4072
rect 13688 4032 79364 4060
rect 82556 4032 92480 4060
rect 13688 4020 13694 4032
rect 18322 3952 18328 4004
rect 18380 3992 18386 4004
rect 82556 3992 82584 4032
rect 92474 4020 92480 4032
rect 92532 4020 92538 4072
rect 93302 4020 93308 4072
rect 93360 4060 93366 4072
rect 93762 4060 93768 4072
rect 93360 4032 93768 4060
rect 93360 4020 93366 4032
rect 93762 4020 93768 4032
rect 93820 4020 93826 4072
rect 218054 4060 218060 4072
rect 94516 4032 218060 4060
rect 18380 3964 82584 3992
rect 18380 3952 18386 3964
rect 82630 3952 82636 4004
rect 82688 3992 82694 4004
rect 86954 3992 86960 4004
rect 82688 3964 86960 3992
rect 82688 3952 82694 3964
rect 86954 3952 86960 3964
rect 87012 3952 87018 4004
rect 88518 3952 88524 4004
rect 88576 3992 88582 4004
rect 94516 3992 94544 4032
rect 218054 4020 218060 4032
rect 218112 4020 218118 4072
rect 88576 3964 94544 3992
rect 88576 3952 88582 3964
rect 95694 3952 95700 4004
rect 95752 3992 95758 4004
rect 230474 3992 230480 4004
rect 95752 3964 230480 3992
rect 95752 3952 95758 3964
rect 230474 3952 230480 3964
rect 230532 3952 230538 4004
rect 102134 3924 102140 3936
rect 27540 3896 102140 3924
rect 24302 3816 24308 3868
rect 24360 3856 24366 3868
rect 27540 3856 27568 3896
rect 102134 3884 102140 3896
rect 102192 3884 102198 3936
rect 102778 3884 102784 3936
rect 102836 3924 102842 3936
rect 106274 3924 106280 3936
rect 102836 3896 106280 3924
rect 102836 3884 102842 3896
rect 106274 3884 106280 3896
rect 106332 3884 106338 3936
rect 106366 3884 106372 3936
rect 106424 3924 106430 3936
rect 107562 3924 107568 3936
rect 106424 3896 107568 3924
rect 106424 3884 106430 3896
rect 107562 3884 107568 3896
rect 107620 3884 107626 3936
rect 115658 3884 115664 3936
rect 115716 3924 115722 3936
rect 242894 3924 242900 3936
rect 115716 3896 242900 3924
rect 115716 3884 115722 3896
rect 242894 3884 242900 3896
rect 242952 3884 242958 3936
rect 100754 3856 100760 3868
rect 24360 3828 27568 3856
rect 27632 3828 100760 3856
rect 24360 3816 24366 3828
rect 23106 3748 23112 3800
rect 23164 3788 23170 3800
rect 27632 3788 27660 3828
rect 100754 3816 100760 3828
rect 100812 3816 100818 3868
rect 103974 3816 103980 3868
rect 104032 3856 104038 3868
rect 245654 3856 245660 3868
rect 104032 3828 114784 3856
rect 104032 3816 104038 3828
rect 23164 3760 27660 3788
rect 23164 3748 23170 3760
rect 27890 3748 27896 3800
rect 27948 3788 27954 3800
rect 109034 3788 109040 3800
rect 27948 3760 109040 3788
rect 27948 3748 27954 3760
rect 109034 3748 109040 3760
rect 109092 3748 109098 3800
rect 109770 3748 109776 3800
rect 109828 3788 109834 3800
rect 114646 3788 114652 3800
rect 109828 3760 114652 3788
rect 109828 3748 109834 3760
rect 114646 3748 114652 3760
rect 114704 3748 114710 3800
rect 114756 3788 114784 3828
rect 115676 3828 245660 3856
rect 115676 3788 115704 3828
rect 245654 3816 245660 3828
rect 245712 3816 245718 3868
rect 114756 3760 115704 3788
rect 115842 3748 115848 3800
rect 115900 3788 115906 3800
rect 255314 3788 255320 3800
rect 115900 3760 255320 3788
rect 115900 3748 115906 3760
rect 255314 3748 255320 3760
rect 255372 3748 255378 3800
rect 29086 3680 29092 3732
rect 29144 3720 29150 3732
rect 111794 3720 111800 3732
rect 29144 3692 111800 3720
rect 29144 3680 29150 3692
rect 111794 3680 111800 3692
rect 111852 3680 111858 3732
rect 113542 3680 113548 3732
rect 113600 3720 113606 3732
rect 262214 3720 262220 3732
rect 113600 3692 262220 3720
rect 113600 3680 113606 3692
rect 262214 3680 262220 3692
rect 262272 3680 262278 3732
rect 31478 3612 31484 3664
rect 31536 3652 31542 3664
rect 31536 3624 111104 3652
rect 31536 3612 31542 3624
rect 32674 3544 32680 3596
rect 32732 3584 32738 3596
rect 109770 3584 109776 3596
rect 32732 3556 109776 3584
rect 32732 3544 32738 3556
rect 109770 3544 109776 3556
rect 109828 3544 109834 3596
rect 111076 3584 111104 3624
rect 118234 3612 118240 3664
rect 118292 3652 118298 3664
rect 270494 3652 270500 3664
rect 118292 3624 270500 3652
rect 118292 3612 118298 3624
rect 270494 3612 270500 3624
rect 270552 3612 270558 3664
rect 115934 3584 115940 3596
rect 111076 3556 115940 3584
rect 115934 3544 115940 3556
rect 115992 3544 115998 3596
rect 120626 3544 120632 3596
rect 120684 3584 120690 3596
rect 274634 3584 274640 3596
rect 120684 3556 274640 3584
rect 120684 3544 120690 3556
rect 274634 3544 274640 3556
rect 274692 3544 274698 3596
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10962 3516 10968 3528
rect 10100 3488 10968 3516
rect 10100 3476 10106 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 12342 3516 12348 3528
rect 11296 3488 12348 3516
rect 11296 3476 11302 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16482 3516 16488 3528
rect 16080 3488 16488 3516
rect 16080 3476 16086 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20622 3516 20628 3528
rect 19576 3488 20628 3516
rect 19576 3476 19582 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21910 3516 21916 3528
rect 20772 3488 21916 3516
rect 20772 3476 20778 3488
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 25498 3476 25504 3528
rect 25556 3516 25562 3528
rect 26142 3516 26148 3528
rect 25556 3488 26148 3516
rect 25556 3476 25562 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 34974 3476 34980 3528
rect 35032 3516 35038 3528
rect 121454 3516 121460 3528
rect 35032 3488 121460 3516
rect 35032 3476 35038 3488
rect 121454 3476 121460 3488
rect 121512 3476 121518 3528
rect 121822 3476 121828 3528
rect 121880 3516 121886 3528
rect 277394 3516 277400 3528
rect 121880 3488 277400 3516
rect 121880 3476 121886 3488
rect 277394 3476 277400 3488
rect 277452 3476 277458 3528
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 32398 3448 32404 3460
rect 5316 3420 32404 3448
rect 5316 3408 5322 3420
rect 32398 3408 32404 3420
rect 32456 3408 32462 3460
rect 42150 3408 42156 3460
rect 42208 3448 42214 3460
rect 42702 3448 42708 3460
rect 42208 3420 42708 3448
rect 42208 3408 42214 3420
rect 42702 3408 42708 3420
rect 42760 3408 42766 3460
rect 42794 3408 42800 3460
rect 42852 3448 42858 3460
rect 124122 3448 124128 3460
rect 42852 3420 124128 3448
rect 42852 3408 42858 3420
rect 124122 3408 124128 3420
rect 124180 3408 124186 3460
rect 124214 3408 124220 3460
rect 124272 3448 124278 3460
rect 281534 3448 281540 3460
rect 124272 3420 281540 3448
rect 124272 3408 124278 3420
rect 281534 3408 281540 3420
rect 281592 3408 281598 3460
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 65150 3380 65156 3392
rect 7708 3352 65156 3380
rect 7708 3340 7714 3352
rect 65150 3340 65156 3352
rect 65208 3340 65214 3392
rect 70486 3380 70492 3392
rect 65536 3352 70492 3380
rect 6454 3272 6460 3324
rect 6512 3312 6518 3324
rect 65536 3312 65564 3352
rect 70486 3340 70492 3352
rect 70544 3340 70550 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 71866 3340 71872 3392
rect 71924 3380 71930 3392
rect 72970 3380 72976 3392
rect 71924 3352 72976 3380
rect 71924 3340 71930 3352
rect 72970 3340 72976 3352
rect 73028 3340 73034 3392
rect 77846 3340 77852 3392
rect 77904 3380 77910 3392
rect 78582 3380 78588 3392
rect 77904 3352 78588 3380
rect 77904 3340 77910 3352
rect 78582 3340 78588 3352
rect 78640 3340 78646 3392
rect 79042 3340 79048 3392
rect 79100 3380 79106 3392
rect 79962 3380 79968 3392
rect 79100 3352 79968 3380
rect 79100 3340 79106 3352
rect 79962 3340 79968 3352
rect 80020 3340 80026 3392
rect 81434 3340 81440 3392
rect 81492 3380 81498 3392
rect 204254 3380 204260 3392
rect 81492 3352 204260 3380
rect 81492 3340 81498 3352
rect 204254 3340 204260 3352
rect 204312 3340 204318 3392
rect 6512 3284 65564 3312
rect 6512 3272 6518 3284
rect 65610 3272 65616 3324
rect 65668 3312 65674 3324
rect 74534 3312 74540 3324
rect 65668 3284 74540 3312
rect 65668 3272 65674 3284
rect 74534 3272 74540 3284
rect 74592 3272 74598 3324
rect 75454 3272 75460 3324
rect 75512 3312 75518 3324
rect 194594 3312 194600 3324
rect 75512 3284 194600 3312
rect 75512 3272 75518 3284
rect 194594 3272 194600 3284
rect 194652 3272 194658 3324
rect 4062 3204 4068 3256
rect 4120 3244 4126 3256
rect 4120 3216 65104 3244
rect 4120 3204 4126 3216
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 64966 3176 64972 3188
rect 2924 3148 64972 3176
rect 2924 3136 2930 3148
rect 64966 3136 64972 3148
rect 65024 3136 65030 3188
rect 65076 3176 65104 3216
rect 65150 3204 65156 3256
rect 65208 3244 65214 3256
rect 73154 3244 73160 3256
rect 65208 3216 73160 3244
rect 65208 3204 65214 3216
rect 73154 3204 73160 3216
rect 73212 3204 73218 3256
rect 74258 3204 74264 3256
rect 74316 3244 74322 3256
rect 191834 3244 191840 3256
rect 74316 3216 191840 3244
rect 74316 3204 74322 3216
rect 191834 3204 191840 3216
rect 191892 3204 191898 3256
rect 66254 3176 66260 3188
rect 65076 3148 66260 3176
rect 66254 3136 66260 3148
rect 66312 3136 66318 3188
rect 68278 3136 68284 3188
rect 68336 3176 68342 3188
rect 180794 3176 180800 3188
rect 68336 3148 180800 3176
rect 68336 3136 68342 3148
rect 180794 3136 180800 3148
rect 180852 3136 180858 3188
rect 566 3068 572 3120
rect 624 3108 630 3120
rect 60734 3108 60740 3120
rect 624 3080 60740 3108
rect 624 3068 630 3080
rect 60734 3068 60740 3080
rect 60792 3068 60798 3120
rect 62206 3108 62212 3120
rect 61120 3080 62212 3108
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 61120 3040 61148 3080
rect 62206 3068 62212 3080
rect 62264 3068 62270 3120
rect 67174 3068 67180 3120
rect 67232 3108 67238 3120
rect 179414 3108 179420 3120
rect 67232 3080 179420 3108
rect 67232 3068 67238 3080
rect 179414 3068 179420 3080
rect 179472 3068 179478 3120
rect 1728 3012 61148 3040
rect 1728 3000 1734 3012
rect 61194 3000 61200 3052
rect 61252 3040 61258 3052
rect 168374 3040 168380 3052
rect 61252 3012 168380 3040
rect 61252 3000 61258 3012
rect 168374 3000 168380 3012
rect 168432 3000 168438 3052
rect 36170 2932 36176 2984
rect 36228 2972 36234 2984
rect 42794 2972 42800 2984
rect 36228 2944 42800 2972
rect 36228 2932 36234 2944
rect 42794 2932 42800 2944
rect 42852 2932 42858 2984
rect 43346 2932 43352 2984
rect 43404 2972 43410 2984
rect 43404 2944 46888 2972
rect 43404 2932 43410 2944
rect 46860 2904 46888 2944
rect 46934 2932 46940 2984
rect 46992 2972 46998 2984
rect 48130 2972 48136 2984
rect 46992 2944 48136 2972
rect 46992 2932 46998 2944
rect 48130 2932 48136 2944
rect 48188 2932 48194 2984
rect 50522 2932 50528 2984
rect 50580 2972 50586 2984
rect 50982 2972 50988 2984
rect 50580 2944 50988 2972
rect 50580 2932 50586 2944
rect 50982 2932 50988 2944
rect 51040 2932 51046 2984
rect 54018 2932 54024 2984
rect 54076 2972 54082 2984
rect 55030 2972 55036 2984
rect 54076 2944 55036 2972
rect 54076 2932 54082 2944
rect 55030 2932 55036 2944
rect 55088 2932 55094 2984
rect 55122 2932 55128 2984
rect 55180 2972 55186 2984
rect 140774 2972 140780 2984
rect 55180 2944 140780 2972
rect 55180 2932 55186 2944
rect 140774 2932 140780 2944
rect 140832 2932 140838 2984
rect 136634 2904 136640 2916
rect 46860 2876 136640 2904
rect 136634 2864 136640 2876
rect 136692 2864 136698 2916
rect 38562 2796 38568 2848
rect 38620 2836 38626 2848
rect 128446 2836 128452 2848
rect 38620 2808 128452 2836
rect 38620 2796 38626 2808
rect 128446 2796 128452 2808
rect 128504 2796 128510 2848
rect 45738 2728 45744 2780
rect 45796 2768 45802 2780
rect 55122 2768 55128 2780
rect 45796 2740 55128 2768
rect 45796 2728 45802 2740
rect 55122 2728 55128 2740
rect 55180 2728 55186 2780
rect 109954 1912 109960 1964
rect 110012 1952 110018 1964
rect 115842 1952 115848 1964
rect 110012 1924 115848 1952
rect 110012 1912 110018 1924
rect 115842 1912 115848 1924
rect 115900 1912 115906 1964
rect 92106 552 92112 604
rect 92164 592 92170 604
rect 92474 592 92480 604
rect 92164 564 92480 592
rect 92164 552 92170 564
rect 92474 552 92480 564
rect 92532 552 92538 604
<< via1 >>
rect 57704 700952 57756 701004
rect 170312 700952 170364 701004
rect 58808 700884 58860 700936
rect 202788 700884 202840 700936
rect 57796 700816 57848 700868
rect 218980 700816 219032 700868
rect 58900 700748 58952 700800
rect 267648 700748 267700 700800
rect 59452 700680 59504 700732
rect 283840 700680 283892 700732
rect 59544 700612 59596 700664
rect 105452 700612 105504 700664
rect 136364 700612 136416 700664
rect 364984 700612 365036 700664
rect 58992 700544 59044 700596
rect 332508 700544 332560 700596
rect 57888 700476 57940 700528
rect 348792 700476 348844 700528
rect 59176 700408 59228 700460
rect 397460 700408 397512 700460
rect 8116 700340 8168 700392
rect 13084 700340 13136 700392
rect 59084 700340 59136 700392
rect 413652 700340 413704 700392
rect 59268 700272 59320 700324
rect 462320 700272 462372 700324
rect 58440 700204 58492 700256
rect 89168 700204 89220 700256
rect 136456 700204 136508 700256
rect 235172 700204 235224 700256
rect 58624 700136 58676 700188
rect 154120 700136 154172 700188
rect 58716 700068 58768 700120
rect 137836 700068 137888 700120
rect 58532 700000 58584 700052
rect 72976 700000 73028 700052
rect 40500 699932 40552 699984
rect 42064 699932 42116 699984
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 58164 696940 58216 696992
rect 580172 696940 580224 696992
rect 429200 692792 429252 692844
rect 429936 692792 429988 692844
rect 299664 688576 299716 688628
rect 300124 688576 300176 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 59360 685856 59412 685908
rect 580172 685856 580224 685908
rect 299572 684428 299624 684480
rect 299664 684428 299716 684480
rect 559012 684428 559064 684480
rect 559104 684428 559156 684480
rect 299664 678988 299716 679040
rect 559104 678988 559156 679040
rect 299664 678852 299716 678904
rect 559104 678852 559156 678904
rect 560300 673888 560352 673940
rect 565176 673888 565228 673940
rect 289820 673752 289872 673804
rect 292672 673752 292724 673804
rect 540980 673752 541032 673804
rect 548616 673752 548668 673804
rect 429200 673412 429252 673464
rect 429476 673412 429528 673464
rect 3424 667904 3476 667956
rect 21364 667904 21416 667956
rect 299664 666544 299716 666596
rect 299940 666544 299992 666596
rect 559104 666544 559156 666596
rect 559380 666544 559432 666596
rect 299664 661716 299716 661768
rect 299940 661716 299992 661768
rect 559104 661716 559156 661768
rect 559380 661716 559432 661768
rect 299664 656888 299716 656940
rect 299756 656888 299808 656940
rect 559104 656888 559156 656940
rect 559196 656888 559248 656940
rect 3056 652740 3108 652792
rect 14464 652740 14516 652792
rect 560300 650360 560352 650412
rect 565176 650360 565228 650412
rect 425060 650224 425112 650276
rect 434536 650224 434588 650276
rect 540980 650224 541032 650276
rect 548616 650224 548668 650276
rect 299664 647232 299716 647284
rect 299756 647232 299808 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 299664 640364 299716 640416
rect 299756 640364 299808 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 59636 638936 59688 638988
rect 580172 638936 580224 638988
rect 299572 630640 299624 630692
rect 299756 630640 299808 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 560300 626968 560352 627020
rect 565176 626968 565228 627020
rect 289820 626832 289872 626884
rect 292672 626832 292724 626884
rect 425060 626832 425112 626884
rect 427912 626832 427964 626884
rect 540980 626832 541032 626884
rect 548616 626832 548668 626884
rect 4068 623772 4120 623824
rect 4988 623772 5040 623824
rect 429476 618196 429528 618248
rect 429660 618196 429712 618248
rect 559196 618196 559248 618248
rect 559380 618196 559432 618248
rect 299572 611328 299624 611380
rect 299756 611328 299808 611380
rect 3424 609968 3476 610020
rect 28264 609968 28316 610020
rect 429292 608608 429344 608660
rect 429660 608608 429712 608660
rect 559104 608540 559156 608592
rect 559472 608540 559524 608592
rect 429200 608472 429252 608524
rect 429292 608472 429344 608524
rect 560300 603440 560352 603492
rect 565176 603440 565228 603492
rect 289820 603304 289872 603356
rect 292672 603304 292724 603356
rect 425060 603304 425112 603356
rect 429936 603304 429988 603356
rect 540980 603304 541032 603356
rect 548616 603304 548668 603356
rect 299664 599020 299716 599072
rect 299848 599020 299900 599072
rect 429200 598952 429252 599004
rect 429384 598952 429436 599004
rect 299664 598884 299716 598936
rect 299848 598884 299900 598936
rect 429200 598816 429252 598868
rect 429384 598816 429436 598868
rect 559196 597524 559248 597576
rect 559380 597524 559432 597576
rect 3240 594804 3292 594856
rect 17316 594804 17368 594856
rect 59728 592016 59780 592068
rect 580172 592016 580224 592068
rect 299664 589296 299716 589348
rect 299940 589296 299992 589348
rect 429200 589296 429252 589348
rect 429476 589296 429528 589348
rect 559196 589296 559248 589348
rect 559380 589296 559432 589348
rect 299940 582428 299992 582480
rect 559380 582428 559432 582480
rect 299848 582292 299900 582344
rect 559288 582292 559340 582344
rect 58348 579640 58400 579692
rect 580172 579640 580224 579692
rect 429384 579572 429436 579624
rect 429568 579572 429620 579624
rect 429384 569916 429436 569968
rect 429660 569916 429712 569968
rect 429476 563728 429528 563780
rect 429660 563728 429712 563780
rect 299572 563116 299624 563168
rect 559012 563116 559064 563168
rect 299572 562980 299624 563032
rect 559012 562980 559064 563032
rect 429292 560192 429344 560244
rect 429476 560192 429528 560244
rect 58256 556180 58308 556232
rect 580172 556180 580224 556232
rect 263784 554004 263836 554056
rect 378508 554004 378560 554056
rect 507860 554004 507912 554056
rect 513380 554004 513432 554056
rect 133696 553392 133748 553444
rect 139584 553392 139636 553444
rect 259184 553392 259236 553444
rect 263784 553392 263836 553444
rect 299572 553460 299624 553512
rect 378508 553392 378560 553444
rect 382924 553392 382976 553444
rect 389364 553392 389416 553444
rect 507860 553392 507912 553444
rect 558920 553392 558972 553444
rect 299480 553324 299532 553376
rect 559012 553324 559064 553376
rect 3148 552032 3200 552084
rect 32404 552032 32456 552084
rect 429292 550604 429344 550656
rect 429568 550604 429620 550656
rect 558920 550604 558972 550656
rect 559012 550604 559064 550656
rect 139400 550264 139452 550316
rect 266452 550264 266504 550316
rect 302240 550264 302292 550316
rect 389180 550264 389232 550316
rect 516416 550264 516468 550316
rect 270408 549244 270460 549296
rect 302240 549244 302292 549296
rect 299480 549176 299532 549228
rect 299572 549176 299624 549228
rect 150348 546456 150400 546508
rect 187700 546456 187752 546508
rect 399484 546456 399536 546508
rect 437480 546456 437532 546508
rect 147588 545096 147640 545148
rect 187700 545096 187752 545148
rect 304448 545096 304500 545148
rect 307668 545096 307720 545148
rect 398104 545096 398156 545148
rect 437480 545096 437532 545148
rect 144828 543736 144880 543788
rect 187700 543736 187752 543788
rect 299572 543736 299624 543788
rect 395344 543736 395396 543788
rect 437480 543736 437532 543788
rect 558920 543736 558972 543788
rect 299572 543600 299624 543652
rect 559012 543600 559064 543652
rect 143448 542376 143500 542428
rect 187700 542376 187752 542428
rect 304356 542376 304408 542428
rect 307208 542376 307260 542428
rect 393964 542376 394016 542428
rect 437480 542376 437532 542428
rect 140688 539656 140740 539708
rect 187792 539656 187844 539708
rect 392584 539656 392636 539708
rect 437572 539656 437624 539708
rect 139308 539588 139360 539640
rect 187700 539588 187752 539640
rect 304264 539588 304316 539640
rect 307668 539588 307720 539640
rect 391204 539588 391256 539640
rect 437480 539588 437532 539640
rect 388444 536800 388496 536852
rect 437480 536800 437532 536852
rect 559012 534012 559064 534064
rect 559196 534012 559248 534064
rect 299572 531292 299624 531344
rect 299664 531292 299716 531344
rect 429200 531292 429252 531344
rect 429476 531292 429528 531344
rect 429476 524424 429528 524476
rect 559196 524424 559248 524476
rect 429568 524356 429620 524408
rect 559288 524356 559340 524408
rect 299480 521636 299532 521688
rect 299756 521636 299808 521688
rect 429384 511980 429436 512032
rect 429660 511980 429712 512032
rect 559104 511980 559156 512032
rect 559380 511980 559432 512032
rect 299480 502324 299532 502376
rect 299756 502324 299808 502376
rect 429476 502324 429528 502376
rect 429660 502324 429712 502376
rect 559196 502324 559248 502376
rect 559380 502324 559432 502376
rect 299480 492600 299532 492652
rect 299664 492600 299716 492652
rect 559104 492600 559156 492652
rect 559196 492600 559248 492652
rect 429476 485800 429528 485852
rect 429568 485732 429620 485784
rect 559104 485732 559156 485784
rect 559196 485732 559248 485784
rect 269120 484372 269172 484424
rect 302884 484372 302936 484424
rect 429568 482944 429620 482996
rect 429660 482944 429712 482996
rect 2964 480224 3016 480276
rect 20076 480224 20128 480276
rect 402244 480224 402296 480276
rect 437480 480224 437532 480276
rect 302976 477504 303028 477556
rect 307116 477504 307168 477556
rect 429660 476076 429712 476128
rect 559012 476076 559064 476128
rect 559196 476076 559248 476128
rect 429568 476008 429620 476060
rect 559104 473288 559156 473340
rect 559196 473288 559248 473340
rect 299664 466420 299716 466472
rect 559196 466420 559248 466472
rect 299756 466352 299808 466404
rect 559104 466352 559156 466404
rect 299756 463632 299808 463684
rect 299848 463632 299900 463684
rect 188896 460164 188948 460216
rect 302976 460164 303028 460216
rect 59820 459484 59872 459536
rect 188896 459484 188948 459536
rect 302976 459484 303028 459536
rect 438124 459484 438176 459536
rect 302884 459416 302936 459468
rect 389180 459416 389232 459468
rect 77300 458124 77352 458176
rect 86316 458124 86368 458176
rect 86868 458124 86920 458176
rect 99380 458124 99432 458176
rect 105360 458124 105412 458176
rect 122748 458124 122800 458176
rect 127072 458124 127124 458176
rect 142068 458124 142120 458176
rect 146944 458124 146996 458176
rect 161388 458124 161440 458176
rect 190460 458124 190512 458176
rect 200028 458124 200080 458176
rect 209780 458124 209832 458176
rect 215300 458124 215352 458176
rect 217232 458124 217284 458176
rect 219348 458124 219400 458176
rect 226340 458124 226392 458176
rect 335360 458124 335412 458176
rect 344744 458124 344796 458176
rect 353300 458124 353352 458176
rect 354036 458124 354088 458176
rect 484400 458124 484452 458176
rect 79968 458056 80020 458108
rect 89076 458056 89128 458108
rect 91100 458056 91152 458108
rect 100576 458056 100628 458108
rect 107660 458056 107712 458108
rect 223580 458056 223632 458108
rect 223672 458056 223724 458108
rect 231860 458056 231912 458108
rect 329104 458056 329156 458108
rect 338028 458056 338080 458108
rect 344376 458056 344428 458108
rect 351920 458056 351972 458108
rect 352748 458056 352800 458108
rect 483020 458056 483072 458108
rect 75828 457988 75880 458040
rect 84200 457988 84252 458040
rect 93584 457988 93636 458040
rect 102784 457988 102836 458040
rect 106280 457988 106332 458040
rect 220820 457988 220872 458040
rect 224316 457988 224368 458040
rect 233240 457988 233292 458040
rect 343548 457988 343600 458040
rect 351828 457988 351880 458040
rect 353944 457988 353996 458040
rect 483204 457988 483256 458040
rect 86868 457920 86920 457972
rect 95792 457920 95844 457972
rect 99380 457920 99432 457972
rect 108764 457920 108816 457972
rect 122748 457920 122800 457972
rect 127072 457920 127124 457972
rect 142068 457920 142120 457972
rect 146944 457920 146996 457972
rect 161388 457920 161440 457972
rect 190460 457920 190512 457972
rect 200028 457920 200080 457972
rect 224960 457920 225012 457972
rect 225880 457920 225932 457972
rect 234620 457920 234672 457972
rect 336556 457920 336608 457972
rect 345940 457920 345992 457972
rect 353668 457920 353720 457972
rect 471796 457920 471848 457972
rect 480444 457920 480496 457972
rect 81348 457852 81400 457904
rect 90180 457852 90232 457904
rect 99472 457852 99524 457904
rect 208216 457852 208268 457904
rect 216680 457852 216732 457904
rect 217140 457852 217192 457904
rect 217232 457852 217284 457904
rect 224316 457852 224368 457904
rect 331312 457852 331364 457904
rect 331864 457852 331916 457904
rect 341248 457852 341300 457904
rect 350540 457852 350592 457904
rect 350632 457852 350684 457904
rect 356060 457852 356112 457904
rect 460204 457852 460256 457904
rect 468760 457852 468812 457904
rect 478328 457852 478380 457904
rect 487160 457852 487212 457904
rect 78588 457784 78640 457836
rect 87880 457784 87932 457836
rect 97172 457784 97224 457836
rect 97908 457784 97960 457836
rect 213092 457784 213144 457836
rect 222568 457784 222620 457836
rect 231860 457784 231912 457836
rect 339040 457784 339092 457836
rect 340880 457784 340932 457836
rect 464988 457784 465040 457836
rect 89076 457716 89128 457768
rect 98552 457716 98604 457768
rect 107660 457716 107712 457768
rect 214012 457716 214064 457768
rect 223672 457716 223724 457768
rect 226432 457716 226484 457768
rect 227168 457716 227220 457768
rect 236000 457716 236052 457768
rect 332600 457716 332652 457768
rect 333152 457716 333204 457768
rect 342536 457716 342588 457768
rect 343548 457716 343600 457768
rect 349252 457716 349304 457768
rect 73068 457648 73120 457700
rect 81900 457648 81952 457700
rect 91100 457648 91152 457700
rect 97908 457648 97960 457700
rect 106280 457648 106332 457700
rect 176568 457648 176620 457700
rect 201500 457648 201552 457700
rect 207756 457648 207808 457700
rect 209688 457648 209740 457700
rect 218888 457648 218940 457700
rect 228364 457648 228416 457700
rect 237380 457648 237432 457700
rect 338028 457648 338080 457700
rect 346860 457648 346912 457700
rect 349712 457716 349764 457768
rect 453488 457716 453540 457768
rect 463056 457716 463108 457768
rect 471336 457716 471388 457768
rect 471520 457784 471572 457836
rect 475476 457784 475528 457836
rect 484400 457784 484452 457836
rect 473452 457716 473504 457768
rect 480260 457716 480312 457768
rect 74172 457580 74224 457632
rect 82820 457580 82872 457632
rect 92480 457580 92532 457632
rect 101864 457580 101916 457632
rect 175188 457580 175240 457632
rect 200212 457580 200264 457632
rect 209136 457580 209188 457632
rect 210516 457580 210568 457632
rect 220176 457580 220228 457632
rect 229560 457580 229612 457632
rect 238760 457580 238812 457632
rect 339868 457580 339920 457632
rect 349252 457580 349304 457632
rect 350632 457580 350684 457632
rect 357440 457648 357492 457700
rect 359464 457648 359516 457700
rect 458180 457648 458232 457700
rect 460388 457648 460440 457700
rect 469956 457648 470008 457700
rect 479432 457648 479484 457700
rect 488540 457648 488592 457700
rect 358820 457580 358872 457632
rect 453304 457580 453356 457632
rect 461768 457580 461820 457632
rect 471796 457580 471848 457632
rect 77208 457512 77260 457564
rect 85488 457512 85540 457564
rect 94780 457512 94832 457564
rect 104256 457512 104308 457564
rect 172428 457512 172480 457564
rect 198740 457512 198792 457564
rect 212448 457512 212500 457564
rect 221372 457512 221424 457564
rect 230480 457512 230532 457564
rect 334072 457512 334124 457564
rect 344376 457512 344428 457564
rect 353668 457512 353720 457564
rect 355048 457512 355100 457564
rect 358084 457512 358136 457564
rect 456800 457512 456852 457564
rect 465172 457512 465224 457564
rect 471244 457512 471296 457564
rect 471336 457512 471388 457564
rect 472256 457580 472308 457632
rect 481640 457580 481692 457632
rect 476304 457512 476356 457564
rect 476948 457512 477000 457564
rect 485780 457512 485832 457564
rect 60740 457444 60792 457496
rect 63684 457444 63736 457496
rect 193864 457444 193916 457496
rect 313740 457444 313792 457496
rect 443000 457444 443052 457496
rect 443644 457444 443696 457496
rect 459560 457444 459612 457496
rect 465724 457444 465776 457496
rect 487160 457444 487212 457496
rect 171048 457376 171100 457428
rect 197360 457376 197412 457428
rect 209044 457376 209096 457428
rect 133788 457308 133840 457360
rect 195980 457308 196032 457360
rect 202144 457308 202196 457360
rect 212448 457308 212500 457360
rect 217140 457376 217192 457428
rect 224960 457376 225012 457428
rect 309784 457376 309836 457428
rect 331220 457376 331272 457428
rect 340880 457376 340932 457428
rect 348240 457376 348292 457428
rect 349712 457376 349764 457428
rect 355324 457376 355376 457428
rect 454040 457376 454092 457428
rect 454684 457376 454736 457428
rect 464988 457376 465040 457428
rect 467104 457376 467156 457428
rect 488540 457376 488592 457428
rect 217600 457308 217652 457360
rect 226432 457308 226484 457360
rect 322204 457308 322256 457360
rect 331312 457308 331364 457360
rect 342904 457308 342956 457360
rect 452660 457308 452712 457360
rect 464344 457308 464396 457360
rect 485780 457308 485832 457360
rect 100576 457240 100628 457292
rect 209780 457240 209832 457292
rect 209872 457240 209924 457292
rect 219348 457240 219400 457292
rect 312544 457240 312596 457292
rect 329840 457240 329892 457292
rect 349804 457240 349856 457292
rect 477500 457240 477552 457292
rect 480260 457240 480312 457292
rect 483112 457240 483164 457292
rect 101864 457172 101916 457224
rect 212540 457172 212592 457224
rect 327908 457172 327960 457224
rect 336556 457172 336608 457224
rect 351184 457172 351236 457224
rect 478880 457172 478932 457224
rect 63408 457104 63460 457156
rect 73160 457104 73212 457156
rect 102784 457104 102836 457156
rect 213920 457104 213972 457156
rect 215208 457104 215260 457156
rect 246304 457104 246356 457156
rect 315304 457104 315356 457156
rect 328460 457104 328512 457156
rect 329288 457104 329340 457156
rect 339040 457104 339092 457156
rect 352564 457104 352616 457156
rect 480536 457104 480588 457156
rect 70308 457036 70360 457088
rect 77300 457036 77352 457088
rect 104256 457036 104308 457088
rect 216680 457036 216732 457088
rect 323584 457036 323636 457088
rect 332600 457036 332652 457088
rect 352656 457036 352708 457088
rect 481640 457036 481692 457088
rect 68928 456968 68980 457020
rect 75920 456968 75972 457020
rect 105360 456968 105412 457020
rect 219440 456968 219492 457020
rect 308404 456968 308456 457020
rect 317420 456968 317472 457020
rect 347044 456968 347096 457020
rect 476120 456968 476172 457020
rect 66168 456900 66220 456952
rect 74724 456900 74776 456952
rect 206836 456900 206888 456952
rect 215300 456900 215352 456952
rect 324964 456900 325016 456952
rect 334072 456900 334124 456952
rect 459376 456900 459428 456952
rect 468024 456900 468076 456952
rect 476304 456900 476356 456952
rect 73068 456832 73120 456884
rect 78772 456832 78824 456884
rect 205456 456832 205508 456884
rect 214012 456832 214064 456884
rect 216588 456832 216640 456884
rect 244924 456832 244976 456884
rect 326344 456832 326396 456884
rect 335452 456832 335504 456884
rect 356704 456832 356756 456884
rect 455420 456832 455472 456884
rect 456708 456832 456760 456884
rect 465172 456832 465224 456884
rect 62028 456764 62080 456816
rect 71780 456764 71832 456816
rect 76564 456764 76616 456816
rect 78680 456764 78732 456816
rect 203524 456764 203576 456816
rect 213092 456764 213144 456816
rect 217968 456764 218020 456816
rect 242164 456764 242216 456816
rect 299848 456764 299900 456816
rect 316684 456764 316736 456816
rect 324320 456764 324372 456816
rect 330484 456764 330536 456816
rect 339868 456764 339920 456816
rect 458088 456764 458140 456816
rect 466644 456832 466696 456884
rect 471152 456832 471204 456884
rect 471244 456832 471296 456884
rect 474832 456832 474884 456884
rect 483020 456832 483072 456884
rect 559012 456764 559064 456816
rect 559196 456764 559248 456816
rect 299756 456696 299808 456748
rect 57612 451256 57664 451308
rect 580172 451256 580224 451308
rect 429476 447176 429528 447228
rect 559196 447176 559248 447228
rect 429476 447040 429528 447092
rect 559196 447040 559248 447092
rect 299664 444388 299716 444440
rect 299848 444388 299900 444440
rect 327632 444388 327684 444440
rect 327724 444388 327776 444440
rect 429384 444388 429436 444440
rect 429476 444388 429528 444440
rect 559104 444388 559156 444440
rect 559196 444388 559248 444440
rect 242348 443232 242400 443284
rect 245108 443232 245160 443284
rect 61108 442892 61160 442944
rect 62028 442892 62080 442944
rect 67824 442892 67876 442944
rect 68928 442892 68980 442944
rect 74632 442892 74684 442944
rect 76564 442892 76616 442944
rect 76932 442892 76984 442944
rect 80060 442892 80112 442944
rect 81440 442892 81492 442944
rect 82820 442892 82872 442944
rect 86868 442892 86920 442944
rect 87972 442892 88024 442944
rect 88248 442892 88300 442944
rect 90456 442892 90508 442944
rect 92388 442892 92440 442944
rect 97264 442892 97316 442944
rect 97908 442892 97960 442944
rect 108580 442892 108632 442944
rect 110328 442892 110380 442944
rect 131304 442892 131356 442944
rect 138020 442892 138072 442944
rect 139308 442892 139360 442944
rect 139400 442892 139452 442944
rect 188344 442892 188396 442944
rect 206008 442892 206060 442944
rect 207756 442892 207808 442944
rect 208216 442892 208268 442944
rect 209136 442892 209188 442944
rect 224868 442892 224920 442944
rect 269396 442892 269448 442944
rect 67548 442824 67600 442876
rect 142528 442824 142580 442876
rect 142620 442824 142672 442876
rect 143448 442824 143500 442876
rect 149336 442824 149388 442876
rect 150348 442824 150400 442876
rect 226248 442824 226300 442876
rect 271696 442824 271748 442876
rect 57060 442756 57112 442808
rect 153936 442756 153988 442808
rect 201500 442756 201552 442808
rect 207664 442756 207716 442808
rect 226156 442756 226208 442808
rect 273904 442756 273956 442808
rect 57152 442688 57204 442740
rect 156144 442688 156196 442740
rect 227628 442688 227680 442740
rect 276204 442688 276256 442740
rect 56784 442620 56836 442672
rect 158444 442620 158496 442672
rect 199200 442620 199252 442672
rect 206284 442620 206336 442672
rect 229008 442620 229060 442672
rect 278412 442620 278464 442672
rect 57336 442552 57388 442604
rect 160652 442552 160704 442604
rect 187884 442552 187936 442604
rect 188988 442552 189040 442604
rect 202788 442552 202840 442604
rect 228640 442552 228692 442604
rect 230388 442552 230440 442604
rect 280712 442552 280764 442604
rect 68836 442484 68888 442536
rect 178776 442484 178828 442536
rect 204168 442484 204220 442536
rect 230848 442484 230900 442536
rect 231768 442484 231820 442536
rect 283012 442484 283064 442536
rect 70124 442416 70176 442468
rect 181076 442416 181128 442468
rect 205548 442416 205600 442468
rect 232780 442416 232832 442468
rect 233056 442416 233108 442468
rect 285220 442416 285272 442468
rect 70216 442348 70268 442400
rect 183376 442348 183428 442400
rect 194692 442348 194744 442400
rect 203524 442348 203576 442400
rect 206928 442348 206980 442400
rect 235448 442348 235500 442400
rect 235908 442348 235960 442400
rect 292028 442348 292080 442400
rect 71688 442280 71740 442332
rect 185584 442280 185636 442332
rect 196900 442280 196952 442332
rect 204904 442280 204956 442332
rect 208308 442280 208360 442332
rect 237656 442280 237708 442332
rect 238668 442280 238720 442332
rect 296536 442280 296588 442332
rect 56968 442212 57020 442264
rect 190092 442212 190144 442264
rect 192392 442212 192444 442264
rect 202144 442212 202196 442264
rect 209688 442212 209740 442264
rect 239956 442212 240008 442264
rect 242072 442212 242124 442264
rect 246212 442212 246264 442264
rect 246304 442212 246356 442264
rect 251272 442212 251324 442264
rect 251364 442212 251416 442264
rect 298836 442212 298888 442264
rect 79140 442144 79192 442196
rect 81348 442144 81400 442196
rect 89628 442144 89680 442196
rect 92756 442144 92808 442196
rect 96528 442144 96580 442196
rect 106372 442144 106424 442196
rect 108948 442144 109000 442196
rect 129004 442144 129056 442196
rect 135812 442144 135864 442196
rect 139400 442144 139452 442196
rect 142528 442144 142580 442196
rect 151636 442144 151688 442196
rect 174268 442144 174320 442196
rect 175188 442144 175240 442196
rect 223488 442144 223540 442196
rect 267096 442144 267148 442196
rect 95148 442076 95200 442128
rect 104072 442076 104124 442128
rect 106188 442076 106240 442128
rect 124496 442076 124548 442128
rect 220728 442076 220780 442128
rect 262588 442076 262640 442128
rect 93676 442008 93728 442060
rect 101864 442008 101916 442060
rect 107568 442008 107620 442060
rect 126704 442008 126756 442060
rect 222108 442008 222160 442060
rect 264888 442008 264940 442060
rect 93768 441940 93820 441992
rect 99564 441940 99616 441992
rect 104808 441940 104860 441992
rect 122196 441940 122248 441992
rect 169760 441940 169812 441992
rect 171048 441940 171100 441992
rect 217876 441940 217928 441992
rect 258080 441940 258132 441992
rect 101956 441872 102008 441924
rect 117688 441872 117740 441924
rect 203708 441872 203760 441924
rect 209044 441872 209096 441924
rect 219348 441872 219400 441924
rect 260288 441872 260340 441924
rect 103428 441804 103480 441856
rect 119896 441804 119948 441856
rect 213828 441804 213880 441856
rect 91008 441736 91060 441788
rect 95056 441736 95108 441788
rect 100668 441736 100720 441788
rect 113180 441736 113232 441788
rect 211068 441736 211120 441788
rect 244464 441736 244516 441788
rect 244924 441804 244976 441856
rect 253572 441804 253624 441856
rect 248604 441736 248656 441788
rect 248696 441736 248748 441788
rect 251364 441736 251416 441788
rect 102048 441668 102100 441720
rect 115388 441668 115440 441720
rect 212448 441668 212500 441720
rect 242072 441668 242124 441720
rect 99288 441600 99340 441652
rect 110880 441600 110932 441652
rect 210976 441600 211028 441652
rect 242256 441600 242308 441652
rect 245108 441600 245160 441652
rect 255780 441600 255832 441652
rect 56968 439832 57020 439884
rect 136364 439832 136416 439884
rect 56784 439764 56836 439816
rect 136456 439764 136508 439816
rect 56876 439696 56928 439748
rect 299664 439696 299716 439748
rect 57060 439628 57112 439680
rect 429384 439628 429436 439680
rect 57980 439560 58032 439612
rect 580356 439560 580408 439612
rect 58072 439492 58124 439544
rect 580724 439492 580776 439544
rect 58164 438948 58216 439000
rect 580080 438948 580132 439000
rect 48964 438880 49016 438932
rect 56600 438880 56652 438932
rect 57520 438880 57572 438932
rect 580632 438880 580684 438932
rect 57244 438268 57296 438320
rect 580540 438268 580592 438320
rect 57336 438200 57388 438252
rect 580816 438200 580868 438252
rect 56692 438132 56744 438184
rect 580264 438132 580316 438184
rect 60004 437996 60056 438048
rect 580356 437996 580408 438048
rect 57428 437928 57480 437980
rect 580448 437928 580500 437980
rect 302792 437384 302844 437436
rect 467104 437384 467156 437436
rect 51724 436092 51776 436144
rect 56600 436092 56652 436144
rect 15844 434732 15896 434784
rect 56692 434732 56744 434784
rect 302792 434664 302844 434716
rect 323492 434664 323544 434716
rect 327540 434664 327592 434716
rect 327632 434664 327684 434716
rect 327724 434664 327776 434716
rect 465724 434664 465776 434716
rect 323492 434460 323544 434512
rect 327724 434460 327776 434512
rect 302792 433236 302844 433288
rect 464344 433236 464396 433288
rect 39304 431944 39356 431996
rect 56692 431944 56744 431996
rect 302792 430516 302844 430568
rect 354036 430516 354088 430568
rect 46204 429156 46256 429208
rect 57152 429156 57204 429208
rect 302792 429088 302844 429140
rect 353944 429088 353996 429140
rect 10324 427796 10376 427848
rect 57152 427796 57204 427848
rect 302792 426368 302844 426420
rect 352748 426368 352800 426420
rect 17224 425076 17276 425128
rect 57152 425076 57204 425128
rect 43444 423648 43496 423700
rect 57152 423648 57204 423700
rect 327540 423648 327592 423700
rect 327632 423648 327684 423700
rect 302792 423580 302844 423632
rect 352656 423580 352708 423632
rect 302792 422220 302844 422272
rect 352564 422220 352616 422272
rect 4896 420928 4948 420980
rect 57152 420928 57204 420980
rect 19984 419500 20036 419552
rect 57152 419500 57204 419552
rect 302792 419432 302844 419484
rect 351184 419432 351236 419484
rect 302792 418072 302844 418124
rect 349804 418072 349856 418124
rect 33784 416780 33836 416832
rect 57152 416780 57204 416832
rect 5080 415420 5132 415472
rect 57152 415420 57204 415472
rect 302792 415352 302844 415404
rect 347044 415352 347096 415404
rect 327540 413924 327592 413976
rect 327724 413924 327776 413976
rect 53104 412632 53156 412684
rect 57152 412632 57204 412684
rect 302792 412564 302844 412616
rect 476212 412564 476264 412616
rect 31024 411272 31076 411324
rect 57152 411272 57204 411324
rect 302792 411204 302844 411256
rect 474740 411204 474792 411256
rect 3516 408484 3568 408536
rect 57152 408484 57204 408536
rect 302792 408416 302844 408468
rect 473360 408416 473412 408468
rect 37924 407124 37976 407176
rect 57152 407124 57204 407176
rect 302792 407056 302844 407108
rect 471980 407056 472032 407108
rect 5172 404336 5224 404388
rect 57152 404336 57204 404388
rect 327540 404336 327592 404388
rect 327724 404336 327776 404388
rect 302700 404268 302752 404320
rect 470600 404268 470652 404320
rect 302792 401548 302844 401600
rect 469220 401548 469272 401600
rect 35164 400188 35216 400240
rect 56692 400188 56744 400240
rect 302792 400120 302844 400172
rect 467932 400120 467984 400172
rect 5264 398828 5316 398880
rect 56692 398828 56744 398880
rect 302792 397400 302844 397452
rect 467840 397400 467892 397452
rect 302516 395972 302568 396024
rect 466460 395972 466512 396024
rect 2780 394748 2832 394800
rect 5356 394748 5408 394800
rect 4068 394680 4120 394732
rect 56508 394680 56560 394732
rect 327540 394612 327592 394664
rect 327632 394612 327684 394664
rect 302700 393252 302752 393304
rect 465080 393252 465132 393304
rect 3884 391960 3936 392012
rect 56600 391960 56652 392012
rect 302792 390464 302844 390516
rect 463700 390464 463752 390516
rect 3240 389172 3292 389224
rect 56600 389172 56652 389224
rect 302792 389104 302844 389156
rect 462320 389104 462372 389156
rect 302516 386316 302568 386368
rect 461032 386316 461084 386368
rect 3056 385024 3108 385076
rect 56600 385024 56652 385076
rect 327632 385024 327684 385076
rect 327816 385024 327868 385076
rect 302516 384956 302568 385008
rect 460940 384956 460992 385008
rect 22100 384888 22152 384940
rect 38660 384888 38712 384940
rect 42892 384888 42944 384940
rect 5356 384820 5408 384872
rect 19340 384820 19392 384872
rect 56600 384752 56652 384804
rect 3332 382168 3384 382220
rect 56600 382168 56652 382220
rect 302792 382168 302844 382220
rect 443644 382168 443696 382220
rect 302608 380808 302660 380860
rect 359464 380808 359516 380860
rect 3332 380740 3384 380792
rect 56600 380740 56652 380792
rect 3148 380604 3200 380656
rect 56600 380604 56652 380656
rect 3976 378088 4028 378140
rect 56600 378088 56652 378140
rect 302792 378088 302844 378140
rect 358084 378088 358136 378140
rect 327632 376728 327684 376780
rect 327816 376728 327868 376780
rect 3792 376660 3844 376712
rect 56600 376660 56652 376712
rect 302792 375300 302844 375352
rect 356704 375300 356756 375352
rect 20076 373940 20128 373992
rect 56600 373940 56652 373992
rect 302792 373940 302844 373992
rect 355324 373940 355376 373992
rect 3700 372512 3752 372564
rect 56600 372512 56652 372564
rect 302332 371152 302384 371204
rect 342904 371152 342956 371204
rect 32404 369792 32456 369844
rect 56600 369792 56652 369844
rect 302608 369792 302660 369844
rect 452752 369792 452804 369844
rect 3608 368432 3660 368484
rect 56600 368432 56652 368484
rect 302792 367004 302844 367056
rect 330484 367004 330536 367056
rect 3424 365644 3476 365696
rect 56600 365644 56652 365696
rect 28264 364284 28316 364336
rect 56600 364284 56652 364336
rect 302516 364284 302568 364336
rect 329288 364284 329340 364336
rect 302424 362856 302476 362908
rect 329104 362856 329156 362908
rect 17316 361496 17368 361548
rect 56600 361496 56652 361548
rect 4988 360136 5040 360188
rect 56600 360136 56652 360188
rect 302332 360136 302384 360188
rect 328092 360136 328144 360188
rect 302516 358708 302568 358760
rect 326344 358708 326396 358760
rect 21364 357348 21416 357400
rect 56600 357348 56652 357400
rect 14464 355988 14516 356040
rect 56600 355988 56652 356040
rect 302792 355988 302844 356040
rect 324964 355988 325016 356040
rect 4804 353200 4856 353252
rect 56600 353200 56652 353252
rect 302792 353200 302844 353252
rect 323584 353200 323636 353252
rect 24768 351840 24820 351892
rect 56600 351840 56652 351892
rect 302424 351840 302476 351892
rect 322204 351840 322256 351892
rect 13084 349052 13136 349104
rect 56600 349052 56652 349104
rect 302700 349052 302752 349104
rect 460388 349052 460440 349104
rect 302516 347692 302568 347744
rect 460204 347692 460256 347744
rect 42064 346332 42116 346384
rect 56600 346332 56652 346384
rect 302792 344972 302844 345024
rect 458824 344972 458876 345024
rect 302792 342184 302844 342236
rect 457444 342184 457496 342236
rect 302424 340824 302476 340876
rect 456064 340824 456116 340876
rect 302700 338036 302752 338088
rect 454684 338036 454736 338088
rect 302516 336676 302568 336728
rect 453488 336676 453540 336728
rect 302792 333888 302844 333940
rect 453304 333888 453356 333940
rect 302516 331100 302568 331152
rect 305828 331100 305880 331152
rect 302332 329400 302384 329452
rect 304448 329400 304500 329452
rect 302516 326884 302568 326936
rect 305736 326884 305788 326936
rect 302332 324436 302384 324488
rect 304356 324436 304408 324488
rect 302332 322668 302384 322720
rect 305644 322668 305696 322720
rect 302332 320084 302384 320136
rect 304264 320084 304316 320136
rect 57796 319472 57848 319524
rect 60004 319472 60056 319524
rect 302700 318316 302752 318368
rect 307024 318316 307076 318368
rect 302792 315936 302844 315988
rect 316040 315936 316092 315988
rect 302792 314576 302844 314628
rect 399484 314576 399536 314628
rect 302700 311788 302752 311840
rect 398104 311788 398156 311840
rect 302792 309068 302844 309120
rect 395344 309068 395396 309120
rect 302792 307708 302844 307760
rect 393964 307708 394016 307760
rect 302792 304920 302844 304972
rect 392584 304920 392636 304972
rect 302792 303560 302844 303612
rect 391204 303560 391256 303612
rect 302700 300772 302752 300824
rect 388444 300772 388496 300824
rect 302792 298052 302844 298104
rect 445760 298052 445812 298104
rect 302608 295876 302660 295928
rect 305920 295876 305972 295928
rect 3056 295264 3108 295316
rect 56692 295264 56744 295316
rect 302792 293904 302844 293956
rect 402244 293904 402296 293956
rect 302516 292476 302568 292528
rect 320272 292476 320324 292528
rect 302700 289756 302752 289808
rect 320180 289756 320232 289808
rect 302792 286968 302844 287020
rect 318800 286968 318852 287020
rect 302700 285268 302752 285320
rect 308404 285268 308456 285320
rect 302516 282820 302568 282872
rect 450544 282820 450596 282872
rect 302516 281460 302568 281512
rect 449164 281460 449216 281512
rect 3424 280100 3476 280152
rect 35164 280100 35216 280152
rect 302332 278672 302384 278724
rect 447784 278672 447836 278724
rect 302608 277312 302660 277364
rect 446404 277312 446456 277364
rect 302792 274592 302844 274644
rect 358820 274592 358872 274644
rect 302516 271804 302568 271856
rect 357440 271804 357492 271856
rect 302516 270444 302568 270496
rect 356060 270444 356112 270496
rect 302332 267656 302384 267708
rect 354680 267656 354732 267708
rect 302608 266296 302660 266348
rect 353300 266296 353352 266348
rect 2780 266228 2832 266280
rect 5264 266228 5316 266280
rect 302792 263508 302844 263560
rect 352012 263508 352064 263560
rect 302516 260788 302568 260840
rect 351920 260788 351972 260840
rect 302424 259360 302476 259412
rect 350540 259360 350592 259412
rect 302332 256640 302384 256692
rect 349160 256640 349212 256692
rect 302516 255212 302568 255264
rect 347780 255212 347832 255264
rect 3424 252492 3476 252544
rect 57152 252492 57204 252544
rect 302792 252492 302844 252544
rect 346400 252492 346452 252544
rect 302792 249704 302844 249756
rect 345020 249704 345072 249756
rect 302424 248344 302476 248396
rect 343732 248344 343784 248396
rect 302700 245556 302752 245608
rect 343640 245556 343692 245608
rect 302516 244196 302568 244248
rect 342260 244196 342312 244248
rect 302792 241408 302844 241460
rect 340880 241408 340932 241460
rect 302792 238688 302844 238740
rect 339500 238688 339552 238740
rect 3424 237328 3476 237380
rect 37924 237328 37976 237380
rect 302424 237328 302476 237380
rect 338120 237328 338172 237380
rect 302700 234540 302752 234592
rect 336832 234540 336884 234592
rect 302516 233180 302568 233232
rect 336740 233180 336792 233232
rect 302792 230392 302844 230444
rect 335360 230392 335412 230444
rect 302792 227672 302844 227724
rect 333980 227672 334032 227724
rect 302792 226244 302844 226296
rect 332600 226244 332652 226296
rect 302700 223524 302752 223576
rect 309784 223524 309836 223576
rect 2780 223048 2832 223100
rect 5172 223048 5224 223100
rect 302792 222096 302844 222148
rect 329932 222096 329984 222148
rect 302792 219376 302844 219428
rect 312544 219376 312596 219428
rect 302792 216588 302844 216640
rect 315304 216588 315356 216640
rect 302792 215228 302844 215280
rect 327080 215228 327132 215280
rect 302608 212440 302660 212492
rect 325700 212440 325752 212492
rect 302792 211080 302844 211132
rect 316684 211080 316736 211132
rect 302792 208292 302844 208344
rect 322940 208292 322992 208344
rect 302792 205572 302844 205624
rect 321560 205572 321612 205624
rect 56968 205504 57020 205556
rect 579896 205368 579948 205420
rect 580172 205368 580224 205420
rect 57152 205164 57204 205216
rect 57152 201560 57204 201612
rect 57152 201424 57204 201476
rect 57520 201560 57572 201612
rect 57520 201424 57572 201476
rect 57796 201424 57848 201476
rect 57980 201356 58032 201408
rect 57060 200812 57112 200864
rect 580816 200812 580868 200864
rect 56968 200744 57020 200796
rect 579988 200744 580040 200796
rect 57704 200676 57756 200728
rect 580540 200676 580592 200728
rect 57152 200608 57204 200660
rect 580172 200608 580224 200660
rect 57520 200540 57572 200592
rect 580080 200540 580132 200592
rect 57980 200472 58032 200524
rect 579896 200472 579948 200524
rect 59820 200404 59872 200456
rect 580356 200404 580408 200456
rect 57244 200064 57296 200116
rect 580724 200064 580776 200116
rect 57612 199996 57664 200048
rect 580908 199996 580960 200048
rect 56876 199928 56928 199980
rect 580632 199928 580684 199980
rect 57888 199860 57940 199912
rect 580448 199860 580500 199912
rect 71688 198636 71740 198688
rect 186320 198636 186372 198688
rect 79968 198568 80020 198620
rect 201132 198568 201184 198620
rect 78588 198500 78640 198552
rect 199016 198500 199068 198552
rect 32404 198432 32456 198484
rect 69480 198432 69532 198484
rect 85488 198432 85540 198484
rect 211804 198432 211856 198484
rect 10968 198364 11020 198416
rect 77944 198364 77996 198416
rect 86868 198364 86920 198416
rect 213920 198364 213972 198416
rect 12348 198296 12400 198348
rect 80060 198296 80112 198348
rect 92388 198296 92440 198348
rect 224500 198296 224552 198348
rect 15108 198228 15160 198280
rect 86500 198228 86552 198280
rect 93768 198228 93820 198280
rect 226616 198228 226668 198280
rect 16488 198160 16540 198212
rect 88616 198160 88668 198212
rect 99196 198160 99248 198212
rect 237288 198160 237340 198212
rect 20628 198092 20680 198144
rect 94964 198092 95016 198144
rect 100668 198092 100720 198144
rect 239404 198092 239456 198144
rect 21916 198024 21968 198076
rect 97080 198024 97132 198076
rect 107568 198024 107620 198076
rect 249984 198024 250036 198076
rect 26148 197956 26200 198008
rect 105544 197956 105596 198008
rect 107476 197956 107528 198008
rect 252100 197956 252152 198008
rect 72976 197888 73028 197940
rect 188436 197888 188488 197940
rect 64788 197820 64840 197872
rect 175648 197820 175700 197872
rect 57888 197752 57940 197804
rect 162952 197752 163004 197804
rect 55128 197684 55180 197736
rect 156512 197684 156564 197736
rect 50988 197616 51040 197668
rect 150164 197616 150216 197668
rect 48136 197548 48188 197600
rect 143816 197548 143868 197600
rect 42708 197480 42760 197532
rect 135352 197480 135404 197532
rect 39948 197412 40000 197464
rect 130292 197412 130344 197464
rect 130384 197412 130436 197464
rect 148048 197412 148100 197464
rect 127624 197344 127676 197396
rect 160836 197344 160888 197396
rect 3148 194488 3200 194540
rect 53104 194488 53156 194540
rect 92204 183540 92256 183592
rect 92388 183540 92440 183592
rect 57336 182112 57388 182164
rect 580172 182112 580224 182164
rect 3240 180752 3292 180804
rect 31024 180752 31076 180804
rect 57428 171028 57480 171080
rect 580172 171028 580224 171080
rect 2780 165452 2832 165504
rect 5080 165452 5132 165504
rect 56784 158652 56836 158704
rect 579804 158652 579856 158704
rect 92204 154504 92256 154556
rect 92388 154504 92440 154556
rect 3148 151716 3200 151768
rect 19984 151716 20036 151768
rect 3240 136552 3292 136604
rect 33784 136552 33836 136604
rect 56600 135192 56652 135244
rect 580172 135192 580224 135244
rect 92112 135124 92164 135176
rect 92388 135124 92440 135176
rect 56692 124108 56744 124160
rect 580172 124108 580224 124160
rect 2780 122340 2832 122392
rect 4896 122340 4948 122392
rect 92204 115880 92256 115932
rect 92388 115880 92440 115932
rect 89628 110780 89680 110832
rect 96528 110780 96580 110832
rect 147588 110644 147640 110696
rect 154488 110644 154540 110696
rect 116032 110508 116084 110560
rect 118792 110508 118844 110560
rect 3240 108944 3292 108996
rect 17224 108944 17276 108996
rect 92204 106292 92256 106344
rect 92388 106292 92440 106344
rect 92388 96568 92440 96620
rect 92572 96568 92624 96620
rect 3424 93780 3476 93832
rect 43444 93780 43496 93832
rect 89628 87252 89680 87304
rect 96528 87252 96580 87304
rect 145564 87116 145616 87168
rect 154488 87116 154540 87168
rect 92388 86980 92440 87032
rect 92572 86980 92624 87032
rect 116032 86980 116084 87032
rect 120816 86980 120868 87032
rect 3424 79976 3476 80028
rect 10324 79976 10376 80028
rect 89628 76236 89680 76288
rect 96528 76236 96580 76288
rect 147588 76100 147640 76152
rect 154488 76100 154540 76152
rect 116032 75964 116084 76016
rect 118792 75964 118844 76016
rect 3332 64812 3384 64864
rect 39304 64812 39356 64864
rect 88892 63860 88944 63912
rect 96528 63860 96580 63912
rect 147588 63724 147640 63776
rect 154488 63724 154540 63776
rect 116032 63588 116084 63640
rect 118792 63588 118844 63640
rect 92204 57876 92256 57928
rect 92388 57876 92440 57928
rect 3424 51008 3476 51060
rect 46204 51008 46256 51060
rect 92204 48288 92256 48340
rect 92388 48288 92440 48340
rect 88892 40332 88944 40384
rect 96528 40332 96580 40384
rect 147588 40196 147640 40248
rect 154488 40196 154540 40248
rect 116032 40060 116084 40112
rect 118792 40060 118844 40112
rect 92204 38564 92256 38616
rect 92388 38564 92440 38616
rect 3424 35844 3476 35896
rect 15844 35844 15896 35896
rect 89628 29316 89680 29368
rect 96528 29316 96580 29368
rect 116032 29044 116084 29096
rect 120816 29044 120868 29096
rect 145012 29044 145064 29096
rect 154488 29044 154540 29096
rect 92204 28976 92256 29028
rect 92388 28976 92440 29028
rect 3148 22040 3200 22092
rect 48964 22040 49016 22092
rect 92204 19252 92256 19304
rect 92388 19252 92440 19304
rect 57796 17892 57848 17944
rect 579804 17892 579856 17944
rect 92204 9664 92256 9716
rect 92388 9664 92440 9716
rect 3424 8236 3476 8288
rect 51724 8236 51776 8288
rect 52828 6672 52880 6724
rect 153200 6672 153252 6724
rect 60004 6604 60056 6656
rect 167000 6604 167052 6656
rect 63592 6536 63644 6588
rect 172520 6536 172572 6588
rect 101588 6468 101640 6520
rect 241520 6468 241572 6520
rect 108764 6400 108816 6452
rect 253940 6400 253992 6452
rect 112352 6332 112404 6384
rect 259460 6332 259512 6384
rect 116124 6264 116176 6316
rect 266360 6264 266412 6316
rect 119436 6196 119488 6248
rect 273260 6196 273312 6248
rect 123024 6128 123076 6180
rect 278780 6128 278832 6180
rect 65524 5448 65576 5500
rect 80060 5516 80112 5568
rect 103980 5516 104032 5568
rect 109408 5516 109460 5568
rect 76656 5448 76708 5500
rect 195980 5448 196032 5500
rect 12440 5380 12492 5432
rect 81440 5380 81492 5432
rect 83832 5380 83884 5432
rect 208400 5380 208452 5432
rect 80060 5312 80112 5364
rect 17224 5244 17276 5296
rect 89720 5244 89772 5296
rect 91192 5312 91244 5364
rect 222200 5312 222252 5364
rect 103980 5244 104032 5296
rect 104256 5244 104308 5296
rect 22008 5176 22060 5228
rect 98000 5176 98052 5228
rect 98828 5176 98880 5228
rect 106464 5244 106516 5296
rect 234620 5244 234672 5296
rect 107660 5176 107712 5228
rect 126612 5176 126664 5228
rect 285680 5176 285732 5228
rect 26700 5108 26752 5160
rect 104072 5108 104124 5160
rect 106280 5108 106332 5160
rect 109408 5108 109460 5160
rect 118608 5108 118660 5160
rect 127808 5108 127860 5160
rect 287060 5108 287112 5160
rect 49332 5040 49384 5092
rect 118516 5040 118568 5092
rect 118792 5040 118844 5092
rect 130384 5040 130436 5092
rect 30288 4972 30340 5024
rect 113180 4972 113232 5024
rect 114744 4972 114796 5024
rect 115848 4972 115900 5024
rect 118884 4972 118936 5024
rect 127624 4972 127676 5024
rect 130200 4972 130252 5024
rect 291200 5040 291252 5092
rect 33876 4904 33928 4956
rect 120080 4904 120132 4956
rect 129004 4904 129056 4956
rect 289820 4972 289872 5024
rect 131396 4904 131448 4956
rect 293960 4904 294012 4956
rect 37372 4836 37424 4888
rect 125600 4836 125652 4888
rect 134892 4836 134944 4888
rect 298100 4836 298152 4888
rect 40960 4768 41012 4820
rect 132500 4768 132552 4820
rect 132592 4768 132644 4820
rect 296720 4768 296772 4820
rect 56416 4700 56468 4752
rect 65524 4700 65576 4752
rect 73068 4700 73120 4752
rect 190460 4700 190512 4752
rect 69480 4632 69532 4684
rect 183560 4632 183612 4684
rect 65984 4564 66036 4616
rect 176660 4564 176712 4616
rect 62396 4496 62448 4548
rect 171140 4496 171192 4548
rect 58808 4428 58860 4480
rect 164240 4428 164292 4480
rect 55220 4360 55272 4412
rect 158720 4360 158772 4412
rect 51632 4292 51684 4344
rect 151820 4292 151872 4344
rect 48228 4224 48280 4276
rect 144920 4224 144972 4276
rect 44548 4156 44600 4208
rect 139400 4156 139452 4208
rect 8852 4088 8904 4140
rect 65616 4088 65668 4140
rect 13636 4020 13688 4072
rect 84200 4088 84252 4140
rect 84936 4088 84988 4140
rect 85488 4088 85540 4140
rect 86132 4088 86184 4140
rect 86868 4088 86920 4140
rect 86960 4088 87012 4140
rect 207020 4088 207072 4140
rect 18328 3952 18380 4004
rect 92480 4020 92532 4072
rect 93308 4020 93360 4072
rect 93768 4020 93820 4072
rect 82636 3952 82688 4004
rect 86960 3952 87012 4004
rect 88524 3952 88576 4004
rect 218060 4020 218112 4072
rect 95700 3952 95752 4004
rect 230480 3952 230532 4004
rect 24308 3816 24360 3868
rect 102140 3884 102192 3936
rect 102784 3884 102836 3936
rect 106280 3884 106332 3936
rect 106372 3884 106424 3936
rect 107568 3884 107620 3936
rect 115664 3884 115716 3936
rect 242900 3884 242952 3936
rect 23112 3748 23164 3800
rect 100760 3816 100812 3868
rect 103980 3816 104032 3868
rect 27896 3748 27948 3800
rect 109040 3748 109092 3800
rect 109776 3748 109828 3800
rect 114652 3748 114704 3800
rect 245660 3816 245712 3868
rect 115848 3748 115900 3800
rect 255320 3748 255372 3800
rect 29092 3680 29144 3732
rect 111800 3680 111852 3732
rect 113548 3680 113600 3732
rect 262220 3680 262272 3732
rect 31484 3612 31536 3664
rect 32680 3544 32732 3596
rect 109776 3544 109828 3596
rect 118240 3612 118292 3664
rect 270500 3612 270552 3664
rect 115940 3544 115992 3596
rect 120632 3544 120684 3596
rect 274640 3544 274692 3596
rect 10048 3476 10100 3528
rect 10968 3476 11020 3528
rect 11244 3476 11296 3528
rect 12348 3476 12400 3528
rect 16028 3476 16080 3528
rect 16488 3476 16540 3528
rect 19524 3476 19576 3528
rect 20628 3476 20680 3528
rect 20720 3476 20772 3528
rect 21916 3476 21968 3528
rect 25504 3476 25556 3528
rect 26148 3476 26200 3528
rect 34980 3476 35032 3528
rect 121460 3476 121512 3528
rect 121828 3476 121880 3528
rect 277400 3476 277452 3528
rect 5264 3408 5316 3460
rect 32404 3408 32456 3460
rect 42156 3408 42208 3460
rect 42708 3408 42760 3460
rect 42800 3408 42852 3460
rect 124128 3408 124180 3460
rect 124220 3408 124272 3460
rect 281540 3408 281592 3460
rect 7656 3340 7708 3392
rect 65156 3340 65208 3392
rect 6460 3272 6512 3324
rect 70492 3340 70544 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 71872 3340 71924 3392
rect 72976 3340 73028 3392
rect 77852 3340 77904 3392
rect 78588 3340 78640 3392
rect 79048 3340 79100 3392
rect 79968 3340 80020 3392
rect 81440 3340 81492 3392
rect 204260 3340 204312 3392
rect 65616 3272 65668 3324
rect 74540 3272 74592 3324
rect 75460 3272 75512 3324
rect 194600 3272 194652 3324
rect 4068 3204 4120 3256
rect 2872 3136 2924 3188
rect 64972 3136 65024 3188
rect 65156 3204 65208 3256
rect 73160 3204 73212 3256
rect 74264 3204 74316 3256
rect 191840 3204 191892 3256
rect 66260 3136 66312 3188
rect 68284 3136 68336 3188
rect 180800 3136 180852 3188
rect 572 3068 624 3120
rect 60740 3068 60792 3120
rect 1676 3000 1728 3052
rect 62212 3068 62264 3120
rect 67180 3068 67232 3120
rect 179420 3068 179472 3120
rect 61200 3000 61252 3052
rect 168380 3000 168432 3052
rect 36176 2932 36228 2984
rect 42800 2932 42852 2984
rect 43352 2932 43404 2984
rect 46940 2932 46992 2984
rect 48136 2932 48188 2984
rect 50528 2932 50580 2984
rect 50988 2932 51040 2984
rect 54024 2932 54076 2984
rect 55036 2932 55088 2984
rect 55128 2932 55180 2984
rect 140780 2932 140832 2984
rect 136640 2864 136692 2916
rect 38568 2796 38620 2848
rect 128452 2796 128504 2848
rect 45744 2728 45796 2780
rect 55128 2728 55180 2780
rect 109960 1912 110012 1964
rect 115848 1912 115900 1964
rect 92112 552 92164 604
rect 92480 552 92532 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700398 8156 703520
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 13084 700392 13136 700398
rect 13084 700334 13136 700340
rect 4802 682272 4858 682281
rect 4802 682207 4858 682216
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 4066 624880 4122 624889
rect 4066 624815 4122 624824
rect 4080 623830 4108 624815
rect 4068 623824 4120 623830
rect 4068 623766 4120 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 2962 481128 3018 481137
rect 2962 481063 3018 481072
rect 2976 480282 3004 481063
rect 2964 480276 3016 480282
rect 2964 480218 3016 480224
rect 3330 438016 3386 438025
rect 3330 437951 3386 437960
rect 3146 423736 3202 423745
rect 3146 423671 3202 423680
rect 2778 395040 2834 395049
rect 2778 394975 2834 394984
rect 2792 394806 2820 394975
rect 2780 394800 2832 394806
rect 2780 394742 2832 394748
rect 3056 385076 3108 385082
rect 3056 385018 3108 385024
rect 3068 366217 3096 385018
rect 3160 380662 3188 423671
rect 3240 389224 3292 389230
rect 3240 389166 3292 389172
rect 3148 380656 3200 380662
rect 3148 380598 3200 380604
rect 3054 366208 3110 366217
rect 3054 366143 3110 366152
rect 3252 337521 3280 389166
rect 3344 382226 3372 437951
rect 3332 382220 3384 382226
rect 3332 382162 3384 382168
rect 3332 380792 3384 380798
rect 3332 380734 3384 380740
rect 3344 380633 3372 380734
rect 3330 380624 3386 380633
rect 3330 380559 3386 380568
rect 3436 365702 3464 567287
rect 3606 538656 3662 538665
rect 3606 538591 3662 538600
rect 3516 408536 3568 408542
rect 3516 408478 3568 408484
rect 3424 365696 3476 365702
rect 3424 365638 3476 365644
rect 3238 337512 3294 337521
rect 3238 337447 3294 337456
rect 3056 295316 3108 295322
rect 3056 295258 3108 295264
rect 3068 294409 3096 295258
rect 3054 294400 3110 294409
rect 3054 294335 3110 294344
rect 3424 280152 3476 280158
rect 3422 280120 3424 280129
rect 3476 280120 3478 280129
rect 3422 280055 3478 280064
rect 2780 266280 2832 266286
rect 2780 266222 2832 266228
rect 2792 265713 2820 266222
rect 2778 265704 2834 265713
rect 2778 265639 2834 265648
rect 3424 252544 3476 252550
rect 3424 252486 3476 252492
rect 3436 251297 3464 252486
rect 3422 251288 3478 251297
rect 3422 251223 3478 251232
rect 3424 237380 3476 237386
rect 3424 237322 3476 237328
rect 3436 237017 3464 237322
rect 3422 237008 3478 237017
rect 3422 236943 3478 236952
rect 2780 223100 2832 223106
rect 2780 223042 2832 223048
rect 2792 222601 2820 223042
rect 2778 222592 2834 222601
rect 2778 222527 2834 222536
rect 3528 208185 3556 408478
rect 3620 368490 3648 538591
rect 3698 509960 3754 509969
rect 3698 509895 3754 509904
rect 3712 372570 3740 509895
rect 3790 495544 3846 495553
rect 3790 495479 3846 495488
rect 3804 376718 3832 495479
rect 3974 452432 4030 452441
rect 3974 452367 4030 452376
rect 3884 392012 3936 392018
rect 3884 391954 3936 391960
rect 3792 376712 3844 376718
rect 3792 376654 3844 376660
rect 3700 372564 3752 372570
rect 3700 372506 3752 372512
rect 3608 368484 3660 368490
rect 3608 368426 3660 368432
rect 3896 308825 3924 391954
rect 3988 378146 4016 452367
rect 4068 394732 4120 394738
rect 4068 394674 4120 394680
rect 3976 378140 4028 378146
rect 3976 378082 4028 378088
rect 4080 323105 4108 394674
rect 4816 353258 4844 682207
rect 4988 623824 5040 623830
rect 4988 623766 5040 623772
rect 4896 420980 4948 420986
rect 4896 420922 4948 420928
rect 4804 353252 4856 353258
rect 4804 353194 4856 353200
rect 4066 323096 4122 323105
rect 4066 323031 4122 323040
rect 3882 308816 3938 308825
rect 3882 308751 3938 308760
rect 3514 208176 3570 208185
rect 3514 208111 3570 208120
rect 3148 194540 3200 194546
rect 3148 194482 3200 194488
rect 3160 193905 3188 194482
rect 3146 193896 3202 193905
rect 3146 193831 3202 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 2780 165504 2832 165510
rect 2780 165446 2832 165452
rect 2792 165073 2820 165446
rect 2778 165064 2834 165073
rect 2778 164999 2834 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3240 136604 3292 136610
rect 3240 136546 3292 136552
rect 3252 136377 3280 136546
rect 3238 136368 3294 136377
rect 3238 136303 3294 136312
rect 4908 122398 4936 420922
rect 5000 360194 5028 623766
rect 10324 427848 10376 427854
rect 10324 427790 10376 427796
rect 5080 415472 5132 415478
rect 5080 415414 5132 415420
rect 4988 360188 5040 360194
rect 4988 360130 5040 360136
rect 5092 165510 5120 415414
rect 5172 404388 5224 404394
rect 5172 404330 5224 404336
rect 5184 223106 5212 404330
rect 5264 398880 5316 398886
rect 5264 398822 5316 398828
rect 5276 266286 5304 398822
rect 5356 394800 5408 394806
rect 5356 394742 5408 394748
rect 5368 384878 5396 394742
rect 5356 384872 5408 384878
rect 5356 384814 5408 384820
rect 5264 266280 5316 266286
rect 5264 266222 5316 266228
rect 5172 223100 5224 223106
rect 5172 223042 5224 223048
rect 5080 165504 5132 165510
rect 5080 165446 5132 165452
rect 2780 122392 2832 122398
rect 2780 122334 2832 122340
rect 4896 122392 4948 122398
rect 4896 122334 4948 122340
rect 2792 122097 2820 122334
rect 2778 122088 2834 122097
rect 2778 122023 2834 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 10336 80034 10364 427790
rect 13096 349110 13124 700334
rect 24320 699718 24348 703520
rect 40512 699990 40540 703520
rect 57704 701004 57756 701010
rect 57704 700946 57756 700952
rect 40500 699984 40552 699990
rect 40500 699926 40552 699932
rect 42064 699984 42116 699990
rect 42064 699926 42116 699932
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 21364 667956 21416 667962
rect 21364 667898 21416 667904
rect 14464 652792 14516 652798
rect 14464 652734 14516 652740
rect 14476 356046 14504 652734
rect 17316 594856 17368 594862
rect 17316 594798 17368 594804
rect 15844 434784 15896 434790
rect 15844 434726 15896 434732
rect 14464 356040 14516 356046
rect 14464 355982 14516 355988
rect 13084 349104 13136 349110
rect 13084 349046 13136 349052
rect 10968 198416 11020 198422
rect 10968 198358 11020 198364
rect 3424 80028 3476 80034
rect 3424 79970 3476 79976
rect 10324 80028 10376 80034
rect 10324 79970 10376 79976
rect 3436 78985 3464 79970
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 4068 3256 4120 3262
rect 4068 3198 4120 3204
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 572 3120 624 3126
rect 572 3062 624 3068
rect 584 480 612 3062
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1688 480 1716 2994
rect 2884 480 2912 3130
rect 4080 480 4108 3198
rect 5276 480 5304 3402
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 6460 3324 6512 3330
rect 6460 3266 6512 3272
rect 6472 480 6500 3266
rect 7668 480 7696 3334
rect 8864 480 8892 4082
rect 10980 3534 11008 198358
rect 12348 198348 12400 198354
rect 12348 198290 12400 198296
rect 12360 3534 12388 198290
rect 15108 198280 15160 198286
rect 15108 198222 15160 198228
rect 12440 5432 12492 5438
rect 12440 5374 12492 5380
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 10060 480 10088 3470
rect 11256 480 11284 3470
rect 12452 480 12480 5374
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13648 480 13676 4014
rect 15120 3482 15148 198222
rect 15856 35902 15884 434726
rect 17224 425128 17276 425134
rect 17224 425070 17276 425076
rect 16488 198212 16540 198218
rect 16488 198154 16540 198160
rect 15844 35896 15896 35902
rect 15844 35838 15896 35844
rect 16500 3534 16528 198154
rect 17236 109002 17264 425070
rect 17328 361554 17356 594798
rect 20076 480276 20128 480282
rect 20076 480218 20128 480224
rect 19984 419552 20036 419558
rect 19984 419494 20036 419500
rect 19340 384872 19392 384878
rect 19338 384840 19340 384849
rect 19392 384840 19394 384849
rect 19338 384775 19394 384784
rect 17316 361548 17368 361554
rect 17316 361490 17368 361496
rect 19996 151774 20024 419494
rect 20088 373998 20116 480218
rect 20076 373992 20128 373998
rect 20076 373934 20128 373940
rect 21376 357406 21404 667898
rect 22100 384940 22152 384946
rect 22100 384882 22152 384888
rect 22112 384849 22140 384882
rect 22098 384840 22154 384849
rect 22098 384775 22154 384784
rect 21364 357400 21416 357406
rect 21364 357342 21416 357348
rect 24780 351898 24808 699654
rect 28264 610020 28316 610026
rect 28264 609962 28316 609968
rect 28276 364342 28304 609962
rect 32404 552084 32456 552090
rect 32404 552026 32456 552032
rect 31024 411324 31076 411330
rect 31024 411266 31076 411272
rect 28264 364336 28316 364342
rect 28264 364278 28316 364284
rect 24768 351892 24820 351898
rect 24768 351834 24820 351840
rect 20628 198144 20680 198150
rect 20628 198086 20680 198092
rect 19984 151768 20036 151774
rect 19984 151710 20036 151716
rect 17224 108996 17276 109002
rect 17224 108938 17276 108944
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 14844 3454 15148 3482
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 14844 480 14872 3454
rect 16040 480 16068 3470
rect 17236 480 17264 5238
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 18340 480 18368 3946
rect 20640 3534 20668 198086
rect 21916 198076 21968 198082
rect 21916 198018 21968 198024
rect 21928 3534 21956 198018
rect 26148 198008 26200 198014
rect 26148 197950 26200 197956
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 19536 480 19564 3470
rect 20732 480 20760 3470
rect 22020 2666 22048 5170
rect 24308 3868 24360 3874
rect 24308 3810 24360 3816
rect 23112 3800 23164 3806
rect 23112 3742 23164 3748
rect 21928 2638 22048 2666
rect 21928 480 21956 2638
rect 23124 480 23152 3742
rect 24320 480 24348 3810
rect 26160 3534 26188 197950
rect 31036 180810 31064 411266
rect 32416 369850 32444 552026
rect 39304 431996 39356 432002
rect 39304 431938 39356 431944
rect 33784 416832 33836 416838
rect 33784 416774 33836 416780
rect 32404 369844 32456 369850
rect 32404 369786 32456 369792
rect 32404 198484 32456 198490
rect 32404 198426 32456 198432
rect 31024 180804 31076 180810
rect 31024 180746 31076 180752
rect 26700 5160 26752 5166
rect 26700 5102 26752 5108
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 25516 480 25544 3470
rect 26712 480 26740 5102
rect 30288 5024 30340 5030
rect 30288 4966 30340 4972
rect 27896 3800 27948 3806
rect 27896 3742 27948 3748
rect 27908 480 27936 3742
rect 29092 3732 29144 3738
rect 29092 3674 29144 3680
rect 29104 480 29132 3674
rect 30300 480 30328 4966
rect 31484 3664 31536 3670
rect 31484 3606 31536 3612
rect 31496 480 31524 3606
rect 32416 3466 32444 198426
rect 33796 136610 33824 416774
rect 37924 407176 37976 407182
rect 37924 407118 37976 407124
rect 35164 400240 35216 400246
rect 35164 400182 35216 400188
rect 35176 280158 35204 400182
rect 35164 280152 35216 280158
rect 35164 280094 35216 280100
rect 37936 237386 37964 407118
rect 38658 384976 38714 384985
rect 38658 384911 38660 384920
rect 38712 384911 38714 384920
rect 38660 384882 38712 384888
rect 37924 237380 37976 237386
rect 37924 237322 37976 237328
rect 33784 136604 33836 136610
rect 33784 136546 33836 136552
rect 39316 64870 39344 431938
rect 42076 346390 42104 699926
rect 57518 546544 57574 546553
rect 57518 546479 57574 546488
rect 57426 545184 57482 545193
rect 57426 545119 57482 545128
rect 56874 543824 56930 543833
rect 56874 543759 56930 543768
rect 56782 540424 56838 540433
rect 56782 540359 56838 540368
rect 56796 442678 56824 540359
rect 56784 442672 56836 442678
rect 56784 442614 56836 442620
rect 56888 442513 56916 543759
rect 57334 542464 57390 542473
rect 57334 542399 57390 542408
rect 57150 539608 57206 539617
rect 57150 539543 57206 539552
rect 57058 537568 57114 537577
rect 57058 537503 57114 537512
rect 56966 480312 57022 480321
rect 56966 480247 57022 480256
rect 56874 442504 56930 442513
rect 56874 442439 56930 442448
rect 56980 442270 57008 480247
rect 57072 442814 57100 537503
rect 57060 442808 57112 442814
rect 57060 442750 57112 442756
rect 57164 442746 57192 539543
rect 57152 442740 57204 442746
rect 57152 442682 57204 442688
rect 57348 442610 57376 542399
rect 57336 442604 57388 442610
rect 57336 442546 57388 442552
rect 57440 442377 57468 545119
rect 57426 442368 57482 442377
rect 57426 442303 57482 442312
rect 56968 442264 57020 442270
rect 57532 442241 57560 546479
rect 57612 451308 57664 451314
rect 57612 451250 57664 451256
rect 56968 442206 57020 442212
rect 57518 442232 57574 442241
rect 57518 442167 57574 442176
rect 56968 439884 57020 439890
rect 56968 439826 57020 439832
rect 56784 439816 56836 439822
rect 56784 439758 56836 439764
rect 56598 438968 56654 438977
rect 48964 438932 49016 438938
rect 56598 438903 56600 438912
rect 48964 438874 49016 438880
rect 56652 438903 56654 438912
rect 56600 438874 56652 438880
rect 46204 429208 46256 429214
rect 46204 429150 46256 429156
rect 43444 423700 43496 423706
rect 43444 423642 43496 423648
rect 42890 384976 42946 384985
rect 42890 384911 42892 384920
rect 42944 384911 42946 384920
rect 42892 384882 42944 384888
rect 42064 346384 42116 346390
rect 42064 346326 42116 346332
rect 42708 197532 42760 197538
rect 42708 197474 42760 197480
rect 39948 197464 40000 197470
rect 39948 197406 40000 197412
rect 39304 64864 39356 64870
rect 39304 64806 39356 64812
rect 33876 4956 33928 4962
rect 33876 4898 33928 4904
rect 32680 3596 32732 3602
rect 32680 3538 32732 3544
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 32692 480 32720 3538
rect 33888 480 33916 4898
rect 37372 4888 37424 4894
rect 37372 4830 37424 4836
rect 34980 3528 35032 3534
rect 34980 3470 35032 3476
rect 34992 480 35020 3470
rect 36176 2984 36228 2990
rect 36176 2926 36228 2932
rect 36188 480 36216 2926
rect 37384 480 37412 4830
rect 39960 3482 39988 197406
rect 40960 4820 41012 4826
rect 40960 4762 41012 4768
rect 39776 3454 39988 3482
rect 38568 2848 38620 2854
rect 38568 2790 38620 2796
rect 38580 480 38608 2790
rect 39776 480 39804 3454
rect 40972 480 41000 4762
rect 42720 3466 42748 197474
rect 43456 93838 43484 423642
rect 43444 93832 43496 93838
rect 43444 93774 43496 93780
rect 46216 51066 46244 429150
rect 48136 197600 48188 197606
rect 48136 197542 48188 197548
rect 46204 51060 46256 51066
rect 46204 51002 46256 51008
rect 44548 4208 44600 4214
rect 44548 4150 44600 4156
rect 42156 3460 42208 3466
rect 42156 3402 42208 3408
rect 42708 3460 42760 3466
rect 42708 3402 42760 3408
rect 42800 3460 42852 3466
rect 42800 3402 42852 3408
rect 42168 480 42196 3402
rect 42812 2990 42840 3402
rect 42800 2984 42852 2990
rect 42800 2926 42852 2932
rect 43352 2984 43404 2990
rect 43352 2926 43404 2932
rect 43364 480 43392 2926
rect 44560 480 44588 4150
rect 48148 2990 48176 197542
rect 48976 22098 49004 438874
rect 56692 438184 56744 438190
rect 56692 438126 56744 438132
rect 51724 436144 51776 436150
rect 56600 436144 56652 436150
rect 51724 436086 51776 436092
rect 56598 436112 56600 436121
rect 56652 436112 56654 436121
rect 50988 197668 51040 197674
rect 50988 197610 51040 197616
rect 48964 22092 49016 22098
rect 48964 22034 49016 22040
rect 49332 5092 49384 5098
rect 49332 5034 49384 5040
rect 48228 4276 48280 4282
rect 48228 4218 48280 4224
rect 46940 2984 46992 2990
rect 46940 2926 46992 2932
rect 48136 2984 48188 2990
rect 48136 2926 48188 2932
rect 45744 2780 45796 2786
rect 45744 2722 45796 2728
rect 45756 480 45784 2722
rect 46952 480 46980 2926
rect 48240 2122 48268 4218
rect 48148 2094 48268 2122
rect 48148 480 48176 2094
rect 49344 480 49372 5034
rect 51000 2990 51028 197610
rect 51736 8294 51764 436086
rect 56598 436047 56654 436056
rect 56704 435962 56732 438126
rect 56612 435934 56732 435962
rect 53104 412684 53156 412690
rect 53104 412626 53156 412632
rect 53116 194546 53144 412626
rect 56506 394768 56562 394777
rect 56506 394703 56508 394712
rect 56560 394703 56562 394712
rect 56508 394674 56560 394680
rect 56612 392714 56640 435934
rect 56692 434784 56744 434790
rect 56690 434752 56692 434761
rect 56744 434752 56746 434761
rect 56690 434687 56746 434696
rect 56690 432032 56746 432041
rect 56690 431967 56692 431976
rect 56744 431967 56746 431976
rect 56692 431938 56744 431944
rect 56690 401024 56746 401033
rect 56690 400959 56746 400968
rect 56704 400246 56732 400959
rect 56692 400240 56744 400246
rect 56692 400182 56744 400188
rect 56690 398984 56746 398993
rect 56690 398919 56746 398928
rect 56704 398886 56732 398919
rect 56692 398880 56744 398886
rect 56692 398822 56744 398828
rect 56690 396808 56746 396817
rect 56690 396743 56746 396752
rect 56520 392686 56640 392714
rect 56520 391898 56548 392686
rect 56598 392592 56654 392601
rect 56598 392527 56654 392536
rect 56612 392018 56640 392527
rect 56600 392012 56652 392018
rect 56600 391954 56652 391960
rect 56520 391870 56640 391898
rect 56612 390674 56640 391870
rect 56520 390646 56640 390674
rect 56520 389042 56548 390646
rect 56598 390552 56654 390561
rect 56598 390487 56654 390496
rect 56612 389230 56640 390487
rect 56600 389224 56652 389230
rect 56600 389166 56652 389172
rect 56520 389014 56640 389042
rect 56612 387841 56640 389014
rect 56598 387832 56654 387841
rect 56598 387767 56654 387776
rect 56598 387696 56654 387705
rect 56598 387631 56654 387640
rect 56612 386458 56640 387631
rect 56520 386430 56640 386458
rect 56520 384010 56548 386430
rect 56598 386336 56654 386345
rect 56598 386271 56654 386280
rect 56612 385082 56640 386271
rect 56600 385076 56652 385082
rect 56600 385018 56652 385024
rect 56600 384804 56652 384810
rect 56600 384746 56652 384752
rect 56612 384169 56640 384746
rect 56598 384160 56654 384169
rect 56598 384095 56654 384104
rect 56520 383982 56640 384010
rect 56612 382378 56640 383982
rect 56520 382350 56640 382378
rect 56520 381970 56548 382350
rect 56600 382220 56652 382226
rect 56600 382162 56652 382168
rect 56612 382129 56640 382162
rect 56598 382120 56654 382129
rect 56598 382055 56654 382064
rect 56520 381942 56640 381970
rect 56612 380798 56640 381942
rect 56600 380792 56652 380798
rect 56600 380734 56652 380740
rect 56600 380656 56652 380662
rect 56600 380598 56652 380604
rect 56612 380089 56640 380598
rect 56598 380080 56654 380089
rect 56598 380015 56654 380024
rect 56600 378140 56652 378146
rect 56600 378082 56652 378088
rect 56612 377913 56640 378082
rect 56598 377904 56654 377913
rect 56598 377839 56654 377848
rect 56600 376712 56652 376718
rect 56600 376654 56652 376660
rect 56612 375873 56640 376654
rect 56598 375864 56654 375873
rect 56598 375799 56654 375808
rect 56600 373992 56652 373998
rect 56600 373934 56652 373940
rect 56612 373697 56640 373934
rect 56598 373688 56654 373697
rect 56598 373623 56654 373632
rect 56600 372564 56652 372570
rect 56600 372506 56652 372512
rect 56612 371657 56640 372506
rect 56598 371648 56654 371657
rect 56598 371583 56654 371592
rect 56600 369844 56652 369850
rect 56600 369786 56652 369792
rect 56612 369481 56640 369786
rect 56598 369472 56654 369481
rect 56598 369407 56654 369416
rect 56600 368484 56652 368490
rect 56600 368426 56652 368432
rect 56612 367441 56640 368426
rect 56598 367432 56654 367441
rect 56598 367367 56654 367376
rect 56600 365696 56652 365702
rect 56600 365638 56652 365644
rect 56612 365265 56640 365638
rect 56598 365256 56654 365265
rect 56598 365191 56654 365200
rect 56600 364336 56652 364342
rect 56600 364278 56652 364284
rect 56612 363225 56640 364278
rect 56598 363216 56654 363225
rect 56598 363151 56654 363160
rect 56600 361548 56652 361554
rect 56600 361490 56652 361496
rect 56612 361049 56640 361490
rect 56598 361040 56654 361049
rect 56598 360975 56654 360984
rect 56600 360188 56652 360194
rect 56600 360130 56652 360136
rect 56612 359009 56640 360130
rect 56598 359000 56654 359009
rect 56598 358935 56654 358944
rect 56600 357400 56652 357406
rect 56600 357342 56652 357348
rect 56612 356833 56640 357342
rect 56598 356824 56654 356833
rect 56598 356759 56654 356768
rect 56600 356040 56652 356046
rect 56600 355982 56652 355988
rect 56612 354793 56640 355982
rect 56598 354784 56654 354793
rect 56598 354719 56654 354728
rect 56600 353252 56652 353258
rect 56600 353194 56652 353200
rect 56612 352617 56640 353194
rect 56598 352608 56654 352617
rect 56598 352543 56654 352552
rect 56600 351892 56652 351898
rect 56600 351834 56652 351840
rect 56612 350577 56640 351834
rect 56598 350568 56654 350577
rect 56598 350503 56654 350512
rect 56600 349104 56652 349110
rect 56600 349046 56652 349052
rect 56612 348401 56640 349046
rect 56598 348392 56654 348401
rect 56598 348327 56654 348336
rect 56600 346384 56652 346390
rect 56598 346352 56600 346361
rect 56652 346352 56654 346361
rect 56598 346287 56654 346296
rect 56704 295322 56732 396743
rect 56796 327321 56824 439758
rect 56876 439748 56928 439754
rect 56876 439690 56928 439696
rect 56782 327312 56838 327321
rect 56782 327247 56838 327256
rect 56888 321065 56916 439690
rect 56874 321056 56930 321065
rect 56874 320991 56930 321000
rect 56980 314809 57008 439826
rect 57060 439680 57112 439686
rect 57060 439622 57112 439628
rect 56966 314800 57022 314809
rect 56966 314735 57022 314744
rect 57072 308417 57100 439622
rect 57520 438932 57572 438938
rect 57520 438874 57572 438880
rect 57244 438320 57296 438326
rect 57244 438262 57296 438268
rect 57150 430536 57206 430545
rect 57150 430471 57206 430480
rect 57164 429214 57192 430471
rect 57152 429208 57204 429214
rect 57152 429150 57204 429156
rect 57150 428496 57206 428505
rect 57150 428431 57206 428440
rect 57164 427854 57192 428431
rect 57152 427848 57204 427854
rect 57152 427790 57204 427796
rect 57150 426320 57206 426329
rect 57150 426255 57206 426264
rect 57164 425134 57192 426255
rect 57152 425128 57204 425134
rect 57152 425070 57204 425076
rect 57150 424280 57206 424289
rect 57150 424215 57206 424224
rect 57164 423706 57192 424215
rect 57152 423700 57204 423706
rect 57152 423642 57204 423648
rect 57150 422104 57206 422113
rect 57150 422039 57206 422048
rect 57164 420986 57192 422039
rect 57152 420980 57204 420986
rect 57152 420922 57204 420928
rect 57150 420064 57206 420073
rect 57150 419999 57206 420008
rect 57164 419558 57192 419999
rect 57152 419552 57204 419558
rect 57152 419494 57204 419500
rect 57150 417888 57206 417897
rect 57150 417823 57206 417832
rect 57164 416838 57192 417823
rect 57152 416832 57204 416838
rect 57152 416774 57204 416780
rect 57150 415848 57206 415857
rect 57150 415783 57206 415792
rect 57164 415478 57192 415783
rect 57152 415472 57204 415478
rect 57152 415414 57204 415420
rect 57150 413672 57206 413681
rect 57150 413607 57206 413616
rect 57164 412690 57192 413607
rect 57152 412684 57204 412690
rect 57152 412626 57204 412632
rect 57150 411632 57206 411641
rect 57150 411567 57206 411576
rect 57164 411330 57192 411567
rect 57152 411324 57204 411330
rect 57152 411266 57204 411272
rect 57150 409456 57206 409465
rect 57150 409391 57206 409400
rect 57164 408542 57192 409391
rect 57152 408536 57204 408542
rect 57152 408478 57204 408484
rect 57150 407416 57206 407425
rect 57150 407351 57206 407360
rect 57164 407182 57192 407351
rect 57152 407176 57204 407182
rect 57152 407118 57204 407124
rect 57150 405240 57206 405249
rect 57150 405175 57206 405184
rect 57164 404394 57192 405175
rect 57152 404388 57204 404394
rect 57152 404330 57204 404336
rect 57150 403200 57206 403209
rect 57150 403135 57206 403144
rect 57058 308408 57114 308417
rect 57058 308343 57114 308352
rect 56692 295316 56744 295322
rect 56692 295258 56744 295264
rect 57164 252550 57192 403135
rect 57256 268433 57284 438262
rect 57336 438252 57388 438258
rect 57336 438194 57388 438200
rect 57242 268424 57298 268433
rect 57242 268359 57298 268368
rect 57348 260001 57376 438194
rect 57428 437980 57480 437986
rect 57428 437922 57480 437928
rect 57334 259992 57390 260001
rect 57334 259927 57390 259936
rect 57440 253745 57468 437922
rect 57426 253736 57482 253745
rect 57426 253671 57482 253680
rect 57152 252544 57204 252550
rect 57152 252486 57204 252492
rect 57532 251569 57560 438874
rect 57624 262041 57652 451250
rect 57716 333713 57744 700946
rect 58808 700936 58860 700942
rect 58808 700878 58860 700884
rect 57796 700868 57848 700874
rect 57796 700810 57848 700816
rect 57702 333704 57758 333713
rect 57702 333639 57758 333648
rect 57808 331537 57836 700810
rect 57888 700528 57940 700534
rect 57888 700470 57940 700476
rect 57794 331528 57850 331537
rect 57794 331463 57850 331472
rect 57796 319524 57848 319530
rect 57796 319466 57848 319472
rect 57610 262032 57666 262041
rect 57610 261967 57666 261976
rect 57808 255785 57836 319466
rect 57900 319025 57928 700470
rect 58440 700256 58492 700262
rect 58440 700198 58492 700204
rect 58164 696992 58216 696998
rect 58164 696934 58216 696940
rect 57980 439612 58032 439618
rect 57980 439554 58032 439560
rect 57886 319016 57942 319025
rect 57886 318951 57942 318960
rect 57992 270473 58020 439554
rect 58072 439544 58124 439550
rect 58072 439486 58124 439492
rect 57978 270464 58034 270473
rect 57978 270399 58034 270408
rect 58084 264217 58112 439486
rect 58176 439385 58204 696934
rect 58348 579692 58400 579698
rect 58348 579634 58400 579640
rect 58256 556232 58308 556238
rect 58256 556174 58308 556180
rect 58162 439376 58218 439385
rect 58162 439311 58218 439320
rect 58164 439000 58216 439006
rect 58164 438942 58216 438948
rect 58070 264208 58126 264217
rect 58070 264143 58126 264152
rect 58176 257961 58204 438942
rect 58268 272649 58296 556174
rect 58360 276865 58388 579634
rect 58452 344185 58480 700198
rect 58624 700188 58676 700194
rect 58624 700130 58676 700136
rect 58532 700052 58584 700058
rect 58532 699994 58584 700000
rect 58438 344176 58494 344185
rect 58438 344111 58494 344120
rect 58544 342145 58572 699994
rect 58530 342136 58586 342145
rect 58530 342071 58586 342080
rect 58636 337929 58664 700130
rect 58716 700120 58768 700126
rect 58716 700062 58768 700068
rect 58622 337920 58678 337929
rect 58622 337855 58678 337864
rect 58728 335753 58756 700062
rect 58714 335744 58770 335753
rect 58714 335679 58770 335688
rect 58820 329497 58848 700878
rect 58900 700800 58952 700806
rect 58900 700742 58952 700748
rect 58806 329488 58862 329497
rect 58806 329423 58862 329432
rect 58912 323105 58940 700742
rect 59452 700732 59504 700738
rect 59452 700674 59504 700680
rect 58992 700596 59044 700602
rect 58992 700538 59044 700544
rect 58898 323096 58954 323105
rect 58898 323031 58954 323040
rect 59004 316849 59032 700538
rect 59176 700460 59228 700466
rect 59176 700402 59228 700408
rect 59084 700392 59136 700398
rect 59084 700334 59136 700340
rect 58990 316840 59046 316849
rect 58990 316775 59046 316784
rect 59096 312633 59124 700334
rect 59082 312624 59138 312633
rect 59082 312559 59138 312568
rect 59188 310593 59216 700402
rect 59268 700324 59320 700330
rect 59268 700266 59320 700272
rect 59174 310584 59230 310593
rect 59174 310519 59230 310528
rect 59280 304201 59308 700266
rect 59360 685908 59412 685914
rect 59360 685850 59412 685856
rect 59266 304192 59322 304201
rect 59266 304127 59322 304136
rect 59372 293729 59400 685850
rect 59464 325281 59492 700674
rect 59544 700664 59596 700670
rect 59544 700606 59596 700612
rect 59556 339969 59584 700606
rect 72988 700058 73016 703520
rect 89180 700262 89208 703520
rect 105464 700670 105492 703520
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 136364 700664 136416 700670
rect 136364 700606 136416 700612
rect 89168 700256 89220 700262
rect 89168 700198 89220 700204
rect 72976 700052 73028 700058
rect 72976 699994 73028 700000
rect 59636 638988 59688 638994
rect 59636 638930 59688 638936
rect 59542 339960 59598 339969
rect 59542 339895 59598 339904
rect 59450 325272 59506 325281
rect 59450 325207 59506 325216
rect 59358 293720 59414 293729
rect 59358 293655 59414 293664
rect 59648 287337 59676 638930
rect 59726 603392 59782 603401
rect 59726 603327 59782 603336
rect 59740 596329 59768 603327
rect 59726 596320 59782 596329
rect 59726 596255 59782 596264
rect 59728 592068 59780 592074
rect 59728 592010 59780 592016
rect 59634 287328 59690 287337
rect 59634 287263 59690 287272
rect 59740 281081 59768 592010
rect 59818 579592 59874 579601
rect 59818 579527 59874 579536
rect 59832 570217 59860 579527
rect 59818 570208 59874 570217
rect 59818 570143 59874 570152
rect 133694 553480 133750 553489
rect 133694 553415 133696 553424
rect 133748 553415 133750 553424
rect 133696 553386 133748 553392
rect 59818 478583 59874 478592
rect 59818 478518 59874 478527
rect 59832 459542 59860 478518
rect 59820 459536 59872 459542
rect 59820 459478 59872 459484
rect 77298 459504 77354 459513
rect 77298 459439 77354 459448
rect 77312 458182 77340 459439
rect 105372 458182 105400 458213
rect 77300 458176 77352 458182
rect 74170 458144 74226 458153
rect 74170 458079 74226 458088
rect 75826 458144 75882 458153
rect 86316 458176 86368 458182
rect 77300 458118 77352 458124
rect 79966 458144 80022 458153
rect 75826 458079 75882 458088
rect 79966 458079 79968 458088
rect 73066 457736 73122 457745
rect 73066 457671 73068 457680
rect 73120 457671 73122 457680
rect 73068 457642 73120 457648
rect 74184 457638 74212 458079
rect 75840 458046 75868 458079
rect 80020 458079 80022 458088
rect 81898 458144 81954 458153
rect 81898 458079 81954 458088
rect 82818 458144 82874 458153
rect 82818 458079 82874 458088
rect 84198 458144 84254 458153
rect 84198 458079 84254 458088
rect 85486 458144 85542 458153
rect 85486 458079 85542 458088
rect 86314 458144 86316 458153
rect 86868 458176 86920 458182
rect 86368 458144 86370 458153
rect 99380 458176 99432 458182
rect 86868 458118 86920 458124
rect 87878 458144 87934 458153
rect 86314 458079 86370 458088
rect 79968 458050 80020 458056
rect 75828 458040 75880 458046
rect 75828 457982 75880 457988
rect 81346 458008 81402 458017
rect 81346 457943 81402 457952
rect 81360 457910 81388 457943
rect 81348 457904 81400 457910
rect 78586 457872 78642 457881
rect 81348 457846 81400 457852
rect 78586 457807 78588 457816
rect 78640 457807 78642 457816
rect 78588 457778 78640 457784
rect 81912 457706 81940 458079
rect 81900 457700 81952 457706
rect 81900 457642 81952 457648
rect 82832 457638 82860 458079
rect 84212 458046 84240 458079
rect 84200 458040 84252 458046
rect 84200 457982 84252 457988
rect 74172 457632 74224 457638
rect 63682 457600 63738 457609
rect 82820 457632 82872 457638
rect 74172 457574 74224 457580
rect 77206 457600 77262 457609
rect 63682 457535 63738 457544
rect 82820 457574 82872 457580
rect 85500 457570 85528 458079
rect 86880 457978 86908 458118
rect 87878 458079 87934 458088
rect 89074 458144 89130 458153
rect 89074 458079 89076 458088
rect 86868 457972 86920 457978
rect 86868 457914 86920 457920
rect 87892 457842 87920 458079
rect 89128 458079 89130 458088
rect 90178 458144 90234 458153
rect 90178 458079 90234 458088
rect 91098 458144 91154 458153
rect 91098 458079 91100 458088
rect 89076 458050 89128 458056
rect 87880 457836 87932 457842
rect 87880 457778 87932 457784
rect 89088 457774 89116 458050
rect 90192 457910 90220 458079
rect 91152 458079 91154 458088
rect 92478 458144 92534 458153
rect 92478 458079 92534 458088
rect 93582 458144 93638 458153
rect 93582 458079 93638 458088
rect 94778 458144 94834 458153
rect 94778 458079 94834 458088
rect 95790 458144 95846 458153
rect 95790 458079 95846 458088
rect 97170 458144 97226 458153
rect 97170 458079 97226 458088
rect 98550 458144 98606 458153
rect 105360 458176 105412 458182
rect 99380 458118 99432 458124
rect 99470 458144 99526 458153
rect 98550 458079 98606 458088
rect 91100 458050 91152 458056
rect 90180 457904 90232 457910
rect 90180 457846 90232 457852
rect 89076 457768 89128 457774
rect 89076 457710 89128 457716
rect 91112 457706 91140 458050
rect 91100 457700 91152 457706
rect 91100 457642 91152 457648
rect 92492 457638 92520 458079
rect 93596 458046 93624 458079
rect 93584 458040 93636 458046
rect 93584 457982 93636 457988
rect 92480 457632 92532 457638
rect 92480 457574 92532 457580
rect 94792 457570 94820 458079
rect 95804 457978 95832 458079
rect 95792 457972 95844 457978
rect 95792 457914 95844 457920
rect 97184 457842 97212 458079
rect 97172 457836 97224 457842
rect 97172 457778 97224 457784
rect 97908 457836 97960 457842
rect 97908 457778 97960 457784
rect 97920 457706 97948 457778
rect 98564 457774 98592 458079
rect 99392 457978 99420 458118
rect 100666 458144 100722 458153
rect 99470 458079 99526 458088
rect 100576 458108 100628 458114
rect 99380 457972 99432 457978
rect 99380 457914 99432 457920
rect 99484 457910 99512 458079
rect 100666 458079 100722 458088
rect 101954 458144 102010 458153
rect 101954 458079 102010 458088
rect 102782 458144 102838 458153
rect 102782 458079 102838 458088
rect 103426 458144 103482 458153
rect 103426 458079 103482 458088
rect 104254 458144 104310 458153
rect 104254 458079 104310 458088
rect 104806 458144 104862 458153
rect 104806 458079 104862 458088
rect 105358 458144 105360 458153
rect 122748 458176 122800 458182
rect 105412 458144 105414 458153
rect 105358 458079 105414 458088
rect 106186 458144 106242 458153
rect 106186 458079 106242 458088
rect 107566 458144 107622 458153
rect 108762 458144 108818 458153
rect 107566 458079 107622 458088
rect 107660 458108 107712 458114
rect 100576 458050 100628 458056
rect 100588 458017 100616 458050
rect 100574 458008 100630 458017
rect 100574 457943 100630 457952
rect 99472 457904 99524 457910
rect 99472 457846 99524 457852
rect 98552 457768 98604 457774
rect 98552 457710 98604 457716
rect 97908 457700 97960 457706
rect 97908 457642 97960 457648
rect 77206 457535 77208 457544
rect 63696 457502 63724 457535
rect 77260 457535 77262 457544
rect 85488 457564 85540 457570
rect 77208 457506 77260 457512
rect 85488 457506 85540 457512
rect 94780 457564 94832 457570
rect 94780 457506 94832 457512
rect 60740 457496 60792 457502
rect 60740 457438 60792 457444
rect 63684 457496 63736 457502
rect 63684 457438 63736 457444
rect 73158 457464 73214 457473
rect 60004 438048 60056 438054
rect 60004 437990 60056 437996
rect 60016 319530 60044 437990
rect 60004 319524 60056 319530
rect 60004 319466 60056 319472
rect 59726 281072 59782 281081
rect 59726 281007 59782 281016
rect 58346 276856 58402 276865
rect 58346 276791 58402 276800
rect 58254 272640 58310 272649
rect 58254 272575 58310 272584
rect 58162 257952 58218 257961
rect 58162 257887 58218 257896
rect 57794 255776 57850 255785
rect 57794 255711 57850 255720
rect 57518 251560 57574 251569
rect 57518 251495 57574 251504
rect 57886 245304 57942 245313
rect 57886 245239 57942 245248
rect 56874 243128 56930 243137
rect 56874 243063 56930 243072
rect 56782 220008 56838 220017
rect 56782 219943 56838 219952
rect 56690 217832 56746 217841
rect 56690 217767 56746 217776
rect 56598 215792 56654 215801
rect 56598 215727 56654 215736
rect 55128 197736 55180 197742
rect 55128 197678 55180 197684
rect 53104 194540 53156 194546
rect 53104 194482 53156 194488
rect 51724 8288 51776 8294
rect 51724 8230 51776 8236
rect 52828 6724 52880 6730
rect 52828 6666 52880 6672
rect 51632 4344 51684 4350
rect 51632 4286 51684 4292
rect 50528 2984 50580 2990
rect 50528 2926 50580 2932
rect 50988 2984 51040 2990
rect 50988 2926 51040 2932
rect 50540 480 50568 2926
rect 51644 480 51672 4286
rect 52840 480 52868 6666
rect 55140 3074 55168 197678
rect 56612 135250 56640 215727
rect 56600 135244 56652 135250
rect 56600 135186 56652 135192
rect 56704 124166 56732 217767
rect 56796 158710 56824 219943
rect 56888 199986 56916 243063
rect 57702 241088 57758 241097
rect 57702 241023 57758 241032
rect 57242 238912 57298 238921
rect 57242 238847 57298 238856
rect 57150 234696 57206 234705
rect 57150 234631 57206 234640
rect 56966 232656 57022 232665
rect 56966 232591 57022 232600
rect 56980 205562 57008 232591
rect 57058 230480 57114 230489
rect 57058 230415 57114 230424
rect 56968 205556 57020 205562
rect 56968 205498 57020 205504
rect 57072 205442 57100 230415
rect 56980 205414 57100 205442
rect 56980 200802 57008 205414
rect 57164 205306 57192 234631
rect 57072 205278 57192 205306
rect 57072 200870 57100 205278
rect 57152 205216 57204 205222
rect 57152 205158 57204 205164
rect 57164 201618 57192 205158
rect 57152 201612 57204 201618
rect 57152 201554 57204 201560
rect 57152 201476 57204 201482
rect 57152 201418 57204 201424
rect 57060 200864 57112 200870
rect 57060 200806 57112 200812
rect 56968 200796 57020 200802
rect 56968 200738 57020 200744
rect 57164 200666 57192 201418
rect 57152 200660 57204 200666
rect 57152 200602 57204 200608
rect 57256 200122 57284 238847
rect 57610 236872 57666 236881
rect 57610 236807 57666 236816
rect 57518 226264 57574 226273
rect 57518 226199 57574 226208
rect 57426 224224 57482 224233
rect 57426 224159 57482 224168
rect 57334 222048 57390 222057
rect 57334 221983 57390 221992
rect 57244 200116 57296 200122
rect 57244 200058 57296 200064
rect 56876 199980 56928 199986
rect 56876 199922 56928 199928
rect 57348 182170 57376 221983
rect 57336 182164 57388 182170
rect 57336 182106 57388 182112
rect 57440 171086 57468 224159
rect 57532 201618 57560 226199
rect 57520 201612 57572 201618
rect 57520 201554 57572 201560
rect 57520 201476 57572 201482
rect 57520 201418 57572 201424
rect 57532 200598 57560 201418
rect 57520 200592 57572 200598
rect 57520 200534 57572 200540
rect 57624 200054 57652 236807
rect 57716 200734 57744 241023
rect 57794 228440 57850 228449
rect 57794 228375 57850 228384
rect 57808 201482 57836 228375
rect 57796 201476 57848 201482
rect 57796 201418 57848 201424
rect 57794 201104 57850 201113
rect 57794 201039 57850 201048
rect 57704 200728 57756 200734
rect 57704 200670 57756 200676
rect 57612 200048 57664 200054
rect 57612 199990 57664 199996
rect 57428 171080 57480 171086
rect 57428 171022 57480 171028
rect 56784 158704 56836 158710
rect 56784 158646 56836 158652
rect 56692 124160 56744 124166
rect 56692 124102 56744 124108
rect 57808 17950 57836 201039
rect 57900 199918 57928 245239
rect 59818 205048 59874 205057
rect 59818 204983 59874 204992
rect 57980 201408 58032 201414
rect 57980 201350 58032 201356
rect 57992 200530 58020 201350
rect 57980 200524 58032 200530
rect 57980 200466 58032 200472
rect 59832 200462 59860 204983
rect 60752 200682 60780 457438
rect 73158 457399 73214 457408
rect 75918 457464 75974 457473
rect 75918 457399 75974 457408
rect 71778 457192 71834 457201
rect 63408 457156 63460 457162
rect 73172 457162 73200 457399
rect 71778 457127 71834 457136
rect 73160 457156 73212 457162
rect 63408 457098 63460 457104
rect 62028 456816 62080 456822
rect 62028 456758 62080 456764
rect 62040 442950 62068 456758
rect 61108 442944 61160 442950
rect 61108 442886 61160 442892
rect 62028 442944 62080 442950
rect 62028 442886 62080 442892
rect 61120 439892 61148 442886
rect 63420 439906 63448 457098
rect 70308 457088 70360 457094
rect 70214 457056 70270 457065
rect 68928 457020 68980 457026
rect 70308 457030 70360 457036
rect 70214 456991 70270 457000
rect 68928 456962 68980 456968
rect 66168 456952 66220 456958
rect 66168 456894 66220 456900
rect 67546 456920 67602 456929
rect 63342 439878 63448 439906
rect 66180 439770 66208 456894
rect 67546 456855 67602 456864
rect 68834 456920 68890 456929
rect 68834 456855 68890 456864
rect 67560 442882 67588 456855
rect 67824 442944 67876 442950
rect 67824 442886 67876 442892
rect 67548 442876 67600 442882
rect 67548 442818 67600 442824
rect 67836 439892 67864 442886
rect 68848 442542 68876 456855
rect 68940 442950 68968 456962
rect 70122 456920 70178 456929
rect 70122 456855 70178 456864
rect 68928 442944 68980 442950
rect 68928 442886 68980 442892
rect 68836 442536 68888 442542
rect 68836 442478 68888 442484
rect 70136 442474 70164 456855
rect 70124 442468 70176 442474
rect 70124 442410 70176 442416
rect 70228 442406 70256 456991
rect 70216 442400 70268 442406
rect 70216 442342 70268 442348
rect 70320 439906 70348 457030
rect 71686 456920 71742 456929
rect 71686 456855 71742 456864
rect 71700 442338 71728 456855
rect 71792 456822 71820 457127
rect 73160 457098 73212 457104
rect 74722 457056 74778 457065
rect 75932 457026 75960 457399
rect 100588 457298 100616 457943
rect 100576 457292 100628 457298
rect 100576 457234 100628 457240
rect 77298 457192 77354 457201
rect 77298 457127 77354 457136
rect 95146 457192 95202 457201
rect 95146 457127 95202 457136
rect 99286 457192 99342 457201
rect 99286 457127 99342 457136
rect 77312 457094 77340 457127
rect 77300 457088 77352 457094
rect 77300 457030 77352 457036
rect 78770 457056 78826 457065
rect 74722 456991 74778 457000
rect 75920 457020 75972 457026
rect 74736 456958 74764 456991
rect 78770 456991 78826 457000
rect 93766 457056 93822 457065
rect 93766 456991 93822 457000
rect 75920 456962 75972 456968
rect 74724 456952 74776 456958
rect 74724 456894 74776 456900
rect 78678 456920 78734 456929
rect 73068 456884 73120 456890
rect 78784 456890 78812 456991
rect 80058 456920 80114 456929
rect 78678 456855 78734 456864
rect 78772 456884 78824 456890
rect 73068 456826 73120 456832
rect 71780 456816 71832 456822
rect 71780 456758 71832 456764
rect 71688 442332 71740 442338
rect 71688 442274 71740 442280
rect 70150 439878 70348 439906
rect 73080 439770 73108 456826
rect 78692 456822 78720 456855
rect 80058 456855 80114 456864
rect 81438 456920 81494 456929
rect 81438 456855 81494 456864
rect 82818 456920 82874 456929
rect 82818 456855 82874 456864
rect 84198 456920 84254 456929
rect 84198 456855 84254 456864
rect 86222 456920 86278 456929
rect 86222 456855 86278 456864
rect 86866 456920 86922 456929
rect 86866 456855 86922 456864
rect 88246 456920 88302 456929
rect 88246 456855 88302 456864
rect 89626 456920 89682 456929
rect 89626 456855 89682 456864
rect 91006 456920 91062 456929
rect 91006 456855 91062 456864
rect 92386 456920 92442 456929
rect 92386 456855 92442 456864
rect 93674 456920 93730 456929
rect 93674 456855 93730 456864
rect 78772 456826 78824 456832
rect 76564 456816 76616 456822
rect 76564 456758 76616 456764
rect 78680 456816 78732 456822
rect 78680 456758 78732 456764
rect 76576 442950 76604 456758
rect 80072 442950 80100 456855
rect 81452 443034 81480 456855
rect 81360 443006 81480 443034
rect 74632 442944 74684 442950
rect 74632 442886 74684 442892
rect 76564 442944 76616 442950
rect 76564 442886 76616 442892
rect 76932 442944 76984 442950
rect 76932 442886 76984 442892
rect 80060 442944 80112 442950
rect 80060 442886 80112 442892
rect 74644 439892 74672 442886
rect 76944 439892 76972 442886
rect 81360 442202 81388 443006
rect 82832 442950 82860 456855
rect 81440 442944 81492 442950
rect 81440 442886 81492 442892
rect 82820 442944 82872 442950
rect 82820 442886 82872 442892
rect 79140 442196 79192 442202
rect 79140 442138 79192 442144
rect 81348 442196 81400 442202
rect 81348 442138 81400 442144
rect 79152 439892 79180 442138
rect 81452 439892 81480 442886
rect 84212 441674 84240 456855
rect 84120 441646 84240 441674
rect 84120 439906 84148 441646
rect 86236 439906 86264 456855
rect 86880 442950 86908 456855
rect 88260 442950 88288 456855
rect 86868 442944 86920 442950
rect 86868 442886 86920 442892
rect 87972 442944 88024 442950
rect 87972 442886 88024 442892
rect 88248 442944 88300 442950
rect 88248 442886 88300 442892
rect 83766 439878 84148 439906
rect 85974 439878 86264 439906
rect 87984 439906 88012 442886
rect 89640 442202 89668 456855
rect 90456 442944 90508 442950
rect 90456 442886 90508 442892
rect 89628 442196 89680 442202
rect 89628 442138 89680 442144
rect 87984 439878 88274 439906
rect 90468 439892 90496 442886
rect 91020 441794 91048 456855
rect 92400 442950 92428 456855
rect 92388 442944 92440 442950
rect 92388 442886 92440 442892
rect 92756 442196 92808 442202
rect 92756 442138 92808 442144
rect 91008 441788 91060 441794
rect 91008 441730 91060 441736
rect 92768 439892 92796 442138
rect 93688 442066 93716 456855
rect 93676 442060 93728 442066
rect 93676 442002 93728 442008
rect 93780 441998 93808 456991
rect 95160 442134 95188 457127
rect 96526 456920 96582 456929
rect 96526 456855 96582 456864
rect 97906 456920 97962 456929
rect 97906 456855 97962 456864
rect 96540 442202 96568 456855
rect 97920 442950 97948 456855
rect 97264 442944 97316 442950
rect 97264 442886 97316 442892
rect 97908 442944 97960 442950
rect 97908 442886 97960 442892
rect 96528 442196 96580 442202
rect 96528 442138 96580 442144
rect 95148 442128 95200 442134
rect 95148 442070 95200 442076
rect 93768 441992 93820 441998
rect 93768 441934 93820 441940
rect 95056 441788 95108 441794
rect 95056 441730 95108 441736
rect 95068 439892 95096 441730
rect 97276 439892 97304 442886
rect 99300 441658 99328 457127
rect 99564 441992 99616 441998
rect 99564 441934 99616 441940
rect 99288 441652 99340 441658
rect 99288 441594 99340 441600
rect 99576 439892 99604 441934
rect 100680 441794 100708 458079
rect 101862 457872 101918 457881
rect 101862 457807 101918 457816
rect 101876 457638 101904 457807
rect 101864 457632 101916 457638
rect 101864 457574 101916 457580
rect 101876 457230 101904 457574
rect 101864 457224 101916 457230
rect 101864 457166 101916 457172
rect 101864 442060 101916 442066
rect 101864 442002 101916 442008
rect 100668 441788 100720 441794
rect 100668 441730 100720 441736
rect 101876 439892 101904 442002
rect 101968 441930 101996 458079
rect 102796 458046 102824 458079
rect 102784 458040 102836 458046
rect 102046 458008 102102 458017
rect 102784 457982 102836 457988
rect 102046 457943 102102 457952
rect 101956 441924 102008 441930
rect 101956 441866 102008 441872
rect 102060 441726 102088 457943
rect 102796 457162 102824 457982
rect 102784 457156 102836 457162
rect 102784 457098 102836 457104
rect 103440 441862 103468 458079
rect 104268 457570 104296 458079
rect 104256 457564 104308 457570
rect 104256 457506 104308 457512
rect 104268 457094 104296 457506
rect 104256 457088 104308 457094
rect 104256 457030 104308 457036
rect 104072 442128 104124 442134
rect 104072 442070 104124 442076
rect 103428 441856 103480 441862
rect 103428 441798 103480 441804
rect 102048 441720 102100 441726
rect 102048 441662 102100 441668
rect 104084 439892 104112 442070
rect 104820 441998 104848 458079
rect 105372 457026 105400 458079
rect 105360 457020 105412 457026
rect 105360 456962 105412 456968
rect 106200 442134 106228 458079
rect 106280 458040 106332 458046
rect 106278 458008 106280 458017
rect 106332 458008 106334 458017
rect 106278 457943 106334 457952
rect 106292 457706 106320 457943
rect 106280 457700 106332 457706
rect 106280 457642 106332 457648
rect 106372 442196 106424 442202
rect 106372 442138 106424 442144
rect 106188 442128 106240 442134
rect 106188 442070 106240 442076
rect 104808 441992 104860 441998
rect 104808 441934 104860 441940
rect 106384 439892 106412 442138
rect 107580 442066 107608 458079
rect 108762 458079 108818 458088
rect 110326 458144 110382 458153
rect 122748 458118 122800 458124
rect 127072 458176 127124 458182
rect 127072 458118 127124 458124
rect 110326 458079 110382 458088
rect 107660 458050 107712 458056
rect 107672 458017 107700 458050
rect 107658 458008 107714 458017
rect 108776 457978 108804 458079
rect 108946 458008 109002 458017
rect 107658 457943 107714 457952
rect 108764 457972 108816 457978
rect 107672 457774 107700 457943
rect 108946 457943 109002 457952
rect 108764 457914 108816 457920
rect 107660 457768 107712 457774
rect 107660 457710 107712 457716
rect 108580 442944 108632 442950
rect 108580 442886 108632 442892
rect 107568 442060 107620 442066
rect 107568 442002 107620 442008
rect 108592 439892 108620 442886
rect 108960 442202 108988 457943
rect 110340 442950 110368 458079
rect 122760 457978 122788 458118
rect 127084 457978 127112 458118
rect 122748 457972 122800 457978
rect 122748 457914 122800 457920
rect 127072 457972 127124 457978
rect 127072 457914 127124 457920
rect 133788 457360 133840 457366
rect 133788 457302 133840 457308
rect 110328 442944 110380 442950
rect 110328 442886 110380 442892
rect 131304 442944 131356 442950
rect 131304 442886 131356 442892
rect 108948 442196 109000 442202
rect 108948 442138 109000 442144
rect 129004 442196 129056 442202
rect 129004 442138 129056 442144
rect 124496 442128 124548 442134
rect 124496 442070 124548 442076
rect 122196 441992 122248 441998
rect 122196 441934 122248 441940
rect 117688 441924 117740 441930
rect 117688 441866 117740 441872
rect 113180 441788 113232 441794
rect 113180 441730 113232 441736
rect 110880 441652 110932 441658
rect 110880 441594 110932 441600
rect 110892 439892 110920 441594
rect 113192 439892 113220 441730
rect 115388 441720 115440 441726
rect 115388 441662 115440 441668
rect 115400 439892 115428 441662
rect 117700 439892 117728 441866
rect 119896 441856 119948 441862
rect 119896 441798 119948 441804
rect 119908 439892 119936 441798
rect 122208 439892 122236 441934
rect 124508 439892 124536 442070
rect 126704 442060 126756 442066
rect 126704 442002 126756 442008
rect 126716 439892 126744 442002
rect 129016 439892 129044 442138
rect 131316 439892 131344 442886
rect 133800 439906 133828 457302
rect 135812 442196 135864 442202
rect 135812 442138 135864 442144
rect 133538 439878 133828 439906
rect 135824 439892 135852 442138
rect 136376 439890 136404 700606
rect 136456 700256 136508 700262
rect 136456 700198 136508 700204
rect 136364 439884 136416 439890
rect 136364 439826 136416 439832
rect 136468 439822 136496 700198
rect 137848 700126 137876 703520
rect 154132 700194 154160 703520
rect 170324 701010 170352 703520
rect 170312 701004 170364 701010
rect 170312 700946 170364 700952
rect 202800 700942 202828 703520
rect 202788 700936 202840 700942
rect 202788 700878 202840 700884
rect 218992 700874 219020 703520
rect 218980 700868 219032 700874
rect 218980 700810 219032 700816
rect 235184 700262 235212 703520
rect 267660 700806 267688 703520
rect 267648 700800 267700 700806
rect 267648 700742 267700 700748
rect 283852 700738 283880 703520
rect 283840 700732 283892 700738
rect 283840 700674 283892 700680
rect 235172 700256 235224 700262
rect 235172 700198 235224 700204
rect 154120 700188 154172 700194
rect 154120 700130 154172 700136
rect 137836 700120 137888 700126
rect 137836 700062 137888 700068
rect 300136 688634 300164 703520
rect 332520 700602 332548 703520
rect 332508 700596 332560 700602
rect 332508 700538 332560 700544
rect 348804 700534 348832 703520
rect 364996 700670 365024 703520
rect 364984 700664 365036 700670
rect 364984 700606 365036 700612
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 397472 700466 397500 703520
rect 397460 700460 397512 700466
rect 397460 700402 397512 700408
rect 413664 700398 413692 703520
rect 429856 703474 429884 703520
rect 429856 703446 429976 703474
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 429948 692850 429976 703446
rect 462332 700330 462360 703520
rect 478524 700777 478552 703520
rect 478510 700768 478566 700777
rect 478510 700703 478566 700712
rect 494808 700641 494836 703520
rect 494794 700632 494850 700641
rect 494794 700567 494850 700576
rect 527192 700505 527220 703520
rect 527178 700496 527234 700505
rect 527178 700431 527234 700440
rect 543476 700369 543504 703520
rect 543462 700360 543518 700369
rect 462320 700324 462372 700330
rect 543462 700295 543518 700304
rect 462320 700266 462372 700272
rect 429200 692844 429252 692850
rect 429200 692786 429252 692792
rect 429936 692844 429988 692850
rect 429936 692786 429988 692792
rect 299664 688628 299716 688634
rect 299664 688570 299716 688576
rect 300124 688628 300176 688634
rect 300124 688570 300176 688576
rect 299676 685930 299704 688570
rect 299584 685902 299704 685930
rect 299584 684486 299612 685902
rect 299572 684480 299624 684486
rect 299572 684422 299624 684428
rect 299664 684480 299716 684486
rect 299664 684422 299716 684428
rect 299676 679046 299704 684422
rect 299664 679040 299716 679046
rect 299664 678982 299716 678988
rect 299664 678904 299716 678910
rect 299664 678846 299716 678852
rect 289818 673840 289874 673849
rect 289818 673775 289820 673784
rect 289872 673775 289874 673784
rect 292672 673804 292724 673810
rect 289820 673746 289872 673752
rect 292672 673746 292724 673752
rect 292684 673577 292712 673746
rect 292670 673568 292726 673577
rect 292670 673503 292726 673512
rect 299676 666602 299704 678846
rect 429212 673470 429240 692786
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 559104 684480 559156 684486
rect 559104 684422 559156 684428
rect 559116 679046 559144 684422
rect 559104 679040 559156 679046
rect 559104 678982 559156 678988
rect 559104 678904 559156 678910
rect 559104 678846 559156 678852
rect 553306 673976 553362 673985
rect 553490 673976 553546 673985
rect 553362 673934 553490 673962
rect 553306 673911 553362 673920
rect 553490 673911 553546 673920
rect 540978 673840 541034 673849
rect 540978 673775 540980 673784
rect 541032 673775 541034 673784
rect 548616 673804 548668 673810
rect 540980 673746 541032 673752
rect 548616 673746 548668 673752
rect 548628 673577 548656 673746
rect 548614 673568 548670 673577
rect 548614 673503 548670 673512
rect 429200 673464 429252 673470
rect 429200 673406 429252 673412
rect 429476 673464 429528 673470
rect 429476 673406 429528 673412
rect 299664 666596 299716 666602
rect 299664 666538 299716 666544
rect 299940 666596 299992 666602
rect 299940 666538 299992 666544
rect 299952 661774 299980 666538
rect 299664 661768 299716 661774
rect 299664 661710 299716 661716
rect 299940 661768 299992 661774
rect 299940 661710 299992 661716
rect 299676 656946 299704 661710
rect 299664 656940 299716 656946
rect 299664 656882 299716 656888
rect 299756 656940 299808 656946
rect 299756 656882 299808 656888
rect 299768 647290 299796 656882
rect 425058 650312 425114 650321
rect 425058 650247 425060 650256
rect 425112 650247 425114 650256
rect 425060 650218 425112 650224
rect 429488 647290 429516 673406
rect 559116 666602 559144 678846
rect 560298 673976 560354 673985
rect 560298 673911 560300 673920
rect 560352 673911 560354 673920
rect 565176 673940 565228 673946
rect 560300 673882 560352 673888
rect 565176 673882 565228 673888
rect 565188 673849 565216 673882
rect 565174 673840 565230 673849
rect 572718 673840 572774 673849
rect 565174 673775 565230 673784
rect 572640 673798 572718 673826
rect 572640 673713 572668 673798
rect 572718 673775 572774 673784
rect 572626 673704 572682 673713
rect 572626 673639 572682 673648
rect 559104 666596 559156 666602
rect 559104 666538 559156 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 559392 661774 559420 666538
rect 559104 661768 559156 661774
rect 559104 661710 559156 661716
rect 559380 661768 559432 661774
rect 559380 661710 559432 661716
rect 559116 656946 559144 661710
rect 559104 656940 559156 656946
rect 559104 656882 559156 656888
rect 559196 656940 559248 656946
rect 559196 656882 559248 656888
rect 553306 650448 553362 650457
rect 553490 650448 553546 650457
rect 553362 650406 553490 650434
rect 553306 650383 553362 650392
rect 553490 650383 553546 650392
rect 540978 650312 541034 650321
rect 434536 650276 434588 650282
rect 540978 650247 540980 650256
rect 434536 650218 434588 650224
rect 541032 650247 541034 650256
rect 548616 650276 548668 650282
rect 540980 650218 541032 650224
rect 548616 650218 548668 650224
rect 434548 650185 434576 650218
rect 434534 650176 434590 650185
rect 434534 650111 434590 650120
rect 548628 650049 548656 650218
rect 548614 650040 548670 650049
rect 548614 649975 548670 649984
rect 559208 647290 559236 656882
rect 560298 650448 560354 650457
rect 560298 650383 560300 650392
rect 560352 650383 560354 650392
rect 565176 650412 565228 650418
rect 560300 650354 560352 650360
rect 565176 650354 565228 650360
rect 565188 650321 565216 650354
rect 565174 650312 565230 650321
rect 572718 650312 572774 650321
rect 565174 650247 565230 650256
rect 572640 650270 572718 650298
rect 572640 650185 572668 650270
rect 572718 650247 572774 650256
rect 572626 650176 572682 650185
rect 572626 650111 572682 650120
rect 299664 647284 299716 647290
rect 299664 647226 299716 647232
rect 299756 647284 299808 647290
rect 299756 647226 299808 647232
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 299676 640422 299704 647226
rect 429396 640422 429424 647226
rect 559116 640422 559144 647226
rect 299664 640416 299716 640422
rect 299664 640358 299716 640364
rect 299756 640416 299808 640422
rect 299756 640358 299808 640364
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 299768 630698 299796 640358
rect 429488 630698 429516 640358
rect 559208 630698 559236 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299756 630692 299808 630698
rect 299756 630634 299808 630640
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 299584 630578 299612 630634
rect 429304 630578 429332 630634
rect 559024 630578 559052 630634
rect 299584 630550 299704 630578
rect 429304 630550 429424 630578
rect 559024 630550 559144 630578
rect 289818 626920 289874 626929
rect 289818 626855 289820 626864
rect 289872 626855 289874 626864
rect 292672 626884 292724 626890
rect 289820 626826 289872 626832
rect 292672 626826 292724 626832
rect 292684 626657 292712 626826
rect 292670 626648 292726 626657
rect 292670 626583 292726 626592
rect 299676 621058 299704 630550
rect 425058 626920 425114 626929
rect 425058 626855 425060 626864
rect 425112 626855 425114 626864
rect 427912 626884 427964 626890
rect 425060 626826 425112 626832
rect 427912 626826 427964 626832
rect 427924 626657 427952 626826
rect 427910 626648 427966 626657
rect 427910 626583 427966 626592
rect 429396 621058 429424 630550
rect 553306 627056 553362 627065
rect 553490 627056 553546 627065
rect 553362 627014 553490 627042
rect 553306 626991 553362 627000
rect 553490 626991 553546 627000
rect 540978 626920 541034 626929
rect 540978 626855 540980 626864
rect 541032 626855 541034 626864
rect 548616 626884 548668 626890
rect 540980 626826 541032 626832
rect 548616 626826 548668 626832
rect 548628 626657 548656 626826
rect 548614 626648 548670 626657
rect 548614 626583 548670 626592
rect 559116 621058 559144 630550
rect 560298 627056 560354 627065
rect 560298 626991 560300 627000
rect 560352 626991 560354 627000
rect 565176 627020 565228 627026
rect 560300 626962 560352 626968
rect 565176 626962 565228 626968
rect 565188 626929 565216 626962
rect 565174 626920 565230 626929
rect 572718 626920 572774 626929
rect 565174 626855 565230 626864
rect 572640 626878 572718 626906
rect 572640 626793 572668 626878
rect 572718 626855 572774 626864
rect 572626 626784 572682 626793
rect 572626 626719 572682 626728
rect 299676 621030 299796 621058
rect 429396 621030 429516 621058
rect 559116 621030 559236 621058
rect 299768 611386 299796 621030
rect 429488 618254 429516 621030
rect 559208 618254 559236 621030
rect 429476 618248 429528 618254
rect 429476 618190 429528 618196
rect 429660 618248 429712 618254
rect 429660 618190 429712 618196
rect 559196 618248 559248 618254
rect 559196 618190 559248 618196
rect 559380 618248 559432 618254
rect 559380 618190 559432 618196
rect 299572 611380 299624 611386
rect 299572 611322 299624 611328
rect 299756 611380 299808 611386
rect 299756 611322 299808 611328
rect 299584 611266 299612 611322
rect 299584 611238 299704 611266
rect 289818 603392 289874 603401
rect 289818 603327 289820 603336
rect 289872 603327 289874 603336
rect 292672 603356 292724 603362
rect 289820 603298 289872 603304
rect 292672 603298 292724 603304
rect 292684 603129 292712 603298
rect 292670 603120 292726 603129
rect 292670 603055 292726 603064
rect 299676 599078 299704 611238
rect 429672 608666 429700 618190
rect 559392 608705 559420 618190
rect 559102 608696 559158 608705
rect 429292 608660 429344 608666
rect 429292 608602 429344 608608
rect 429660 608660 429712 608666
rect 559102 608631 559158 608640
rect 559378 608696 559434 608705
rect 559378 608631 559434 608640
rect 429660 608602 429712 608608
rect 429304 608530 429332 608602
rect 559116 608598 559144 608631
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 559472 608592 559524 608598
rect 559472 608534 559524 608540
rect 429200 608524 429252 608530
rect 429200 608466 429252 608472
rect 429292 608524 429344 608530
rect 429292 608466 429344 608472
rect 425058 603392 425114 603401
rect 425058 603327 425060 603336
rect 425112 603327 425114 603336
rect 425060 603298 425112 603304
rect 299664 599072 299716 599078
rect 299664 599014 299716 599020
rect 299848 599072 299900 599078
rect 299848 599014 299900 599020
rect 299860 598942 299888 599014
rect 429212 599010 429240 608466
rect 559484 607186 559512 608534
rect 559392 607158 559512 607186
rect 553398 603528 553454 603537
rect 553398 603463 553454 603472
rect 441526 603392 441582 603401
rect 429936 603356 429988 603362
rect 441526 603327 441582 603336
rect 540978 603392 541034 603401
rect 540978 603327 540980 603336
rect 429936 603298 429988 603304
rect 429948 603265 429976 603298
rect 429934 603256 429990 603265
rect 429934 603191 429990 603200
rect 441540 602993 441568 603327
rect 541032 603327 541034 603336
rect 548616 603356 548668 603362
rect 540980 603298 541032 603304
rect 548616 603298 548668 603304
rect 548628 603129 548656 603298
rect 548614 603120 548670 603129
rect 548614 603055 548670 603064
rect 553306 603120 553362 603129
rect 553412 603106 553440 603463
rect 553362 603078 553440 603106
rect 553306 603055 553362 603064
rect 441526 602984 441582 602993
rect 441526 602919 441582 602928
rect 429200 599004 429252 599010
rect 429200 598946 429252 598952
rect 429384 599004 429436 599010
rect 429384 598946 429436 598952
rect 299664 598936 299716 598942
rect 299664 598878 299716 598884
rect 299848 598936 299900 598942
rect 299848 598878 299900 598884
rect 299676 589354 299704 598878
rect 429396 598874 429424 598946
rect 429200 598868 429252 598874
rect 429200 598810 429252 598816
rect 429384 598868 429436 598874
rect 429384 598810 429436 598816
rect 429212 589354 429240 598810
rect 559392 597582 559420 607158
rect 560298 603528 560354 603537
rect 560298 603463 560300 603472
rect 560352 603463 560354 603472
rect 565176 603492 565228 603498
rect 560300 603434 560352 603440
rect 565176 603434 565228 603440
rect 565188 603401 565216 603434
rect 565174 603392 565230 603401
rect 572718 603392 572774 603401
rect 565174 603327 565230 603336
rect 572640 603350 572718 603378
rect 572640 603265 572668 603350
rect 572718 603327 572774 603336
rect 572626 603256 572682 603265
rect 572626 603191 572682 603200
rect 559196 597576 559248 597582
rect 559196 597518 559248 597524
rect 559380 597576 559432 597582
rect 559380 597518 559432 597524
rect 559208 589354 559236 597518
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 299664 589348 299716 589354
rect 299664 589290 299716 589296
rect 299940 589348 299992 589354
rect 299940 589290 299992 589296
rect 429200 589348 429252 589354
rect 429200 589290 429252 589296
rect 429476 589348 429528 589354
rect 429476 589290 429528 589296
rect 559196 589348 559248 589354
rect 559196 589290 559248 589296
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 299952 582486 299980 589290
rect 299940 582480 299992 582486
rect 299940 582422 299992 582428
rect 429488 582434 429516 589290
rect 559392 582486 559420 589290
rect 559380 582480 559432 582486
rect 429488 582406 429608 582434
rect 559380 582422 559432 582428
rect 299848 582344 299900 582350
rect 299848 582286 299900 582292
rect 299860 572642 299888 582286
rect 429580 579630 429608 582406
rect 559288 582344 559340 582350
rect 559288 582286 559340 582292
rect 429384 579624 429436 579630
rect 429384 579566 429436 579572
rect 429568 579624 429620 579630
rect 429568 579566 429620 579572
rect 299676 572614 299888 572642
rect 299676 569922 299704 572614
rect 429396 569974 429424 579566
rect 559300 572642 559328 582286
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 559116 572614 559328 572642
rect 299584 569894 299704 569922
rect 429384 569968 429436 569974
rect 429384 569910 429436 569916
rect 429660 569968 429712 569974
rect 559116 569922 559144 572614
rect 429660 569910 429712 569916
rect 299584 563174 299612 569894
rect 429672 563786 429700 569910
rect 559024 569894 559144 569922
rect 429476 563780 429528 563786
rect 429476 563722 429528 563728
rect 429660 563780 429712 563786
rect 429660 563722 429712 563728
rect 299572 563168 299624 563174
rect 299572 563110 299624 563116
rect 299572 563032 299624 563038
rect 299572 562974 299624 562980
rect 263784 554056 263836 554062
rect 263784 553998 263836 554004
rect 263796 553489 263824 553998
rect 299584 553518 299612 562974
rect 429488 560250 429516 563722
rect 559024 563174 559052 569894
rect 559012 563168 559064 563174
rect 559012 563110 559064 563116
rect 559012 563032 559064 563038
rect 559012 562974 559064 562980
rect 559024 560266 559052 562974
rect 429292 560244 429344 560250
rect 429292 560186 429344 560192
rect 429476 560244 429528 560250
rect 429476 560186 429528 560192
rect 558932 560238 559052 560266
rect 378508 554056 378560 554062
rect 378508 553998 378560 554004
rect 299572 553512 299624 553518
rect 259182 553480 259238 553489
rect 139584 553444 139636 553450
rect 259182 553415 259184 553424
rect 139584 553386 139636 553392
rect 259236 553415 259238 553424
rect 263782 553480 263838 553489
rect 378520 553489 378548 553998
rect 299572 553454 299624 553460
rect 378506 553480 378562 553489
rect 263782 553415 263784 553424
rect 259184 553386 259236 553392
rect 263836 553415 263838 553424
rect 378506 553415 378508 553424
rect 263784 553386 263836 553392
rect 378560 553415 378562 553424
rect 382922 553480 382978 553489
rect 382922 553415 382924 553424
rect 378508 553386 378560 553392
rect 382976 553415 382978 553424
rect 389364 553444 389416 553450
rect 382924 553386 382976 553392
rect 389364 553386 389416 553392
rect 139400 550316 139452 550322
rect 139400 550258 139452 550264
rect 139412 549953 139440 550258
rect 139398 549944 139454 549953
rect 139398 549879 139454 549888
rect 139596 549794 139624 553386
rect 263796 553355 263824 553386
rect 299480 553376 299532 553382
rect 378520 553355 378548 553386
rect 299480 553318 299532 553324
rect 266452 550316 266504 550322
rect 266452 550258 266504 550264
rect 266464 549953 266492 550258
rect 266450 549944 266506 549953
rect 266450 549879 266506 549888
rect 139412 549766 139624 549794
rect 139308 539640 139360 539646
rect 139308 539582 139360 539588
rect 139320 442950 139348 539582
rect 139412 489569 139440 549766
rect 270406 549400 270462 549409
rect 270406 549335 270462 549344
rect 270420 549302 270448 549335
rect 270408 549296 270460 549302
rect 270408 549238 270460 549244
rect 299492 549234 299520 553318
rect 302240 550316 302292 550322
rect 302240 550258 302292 550264
rect 389180 550316 389232 550322
rect 389180 550258 389232 550264
rect 302252 549302 302280 550258
rect 389192 549953 389220 550258
rect 389178 549944 389234 549953
rect 389178 549879 389234 549888
rect 302240 549296 302292 549302
rect 302240 549238 302292 549244
rect 299480 549228 299532 549234
rect 299480 549170 299532 549176
rect 299572 549228 299624 549234
rect 299572 549170 299624 549176
rect 187698 546544 187754 546553
rect 150348 546508 150400 546514
rect 187698 546479 187700 546488
rect 150348 546450 150400 546456
rect 187752 546479 187754 546488
rect 187700 546450 187752 546456
rect 147588 545148 147640 545154
rect 147588 545090 147640 545096
rect 144828 543788 144880 543794
rect 144828 543730 144880 543736
rect 143448 542428 143500 542434
rect 143448 542370 143500 542376
rect 140688 539708 140740 539714
rect 140688 539650 140740 539656
rect 139398 489560 139454 489569
rect 139398 489495 139454 489504
rect 138020 442944 138072 442950
rect 138020 442886 138072 442892
rect 139308 442944 139360 442950
rect 139308 442886 139360 442892
rect 139400 442944 139452 442950
rect 139400 442886 139452 442892
rect 138032 439892 138060 442886
rect 139412 442202 139440 442886
rect 139400 442196 139452 442202
rect 139400 442138 139452 442144
rect 140700 439906 140728 539650
rect 142068 458176 142120 458182
rect 142068 458118 142120 458124
rect 142080 457978 142108 458118
rect 142068 457972 142120 457978
rect 142068 457914 142120 457920
rect 143460 442882 143488 542370
rect 142528 442876 142580 442882
rect 142528 442818 142580 442824
rect 142620 442876 142672 442882
rect 142620 442818 142672 442824
rect 143448 442876 143500 442882
rect 143448 442818 143500 442824
rect 142540 442202 142568 442818
rect 142528 442196 142580 442202
rect 142528 442138 142580 442144
rect 140346 439878 140728 439906
rect 142632 439892 142660 442818
rect 144840 439892 144868 543730
rect 146944 458176 146996 458182
rect 146944 458118 146996 458124
rect 146956 457978 146984 458118
rect 146944 457972 146996 457978
rect 146944 457914 146996 457920
rect 147600 439906 147628 545090
rect 150360 442882 150388 546450
rect 187698 545184 187754 545193
rect 187698 545119 187700 545128
rect 187752 545119 187754 545128
rect 187700 545090 187752 545096
rect 187698 543824 187754 543833
rect 299584 543794 299612 549170
rect 187698 543759 187700 543768
rect 187752 543759 187754 543768
rect 299572 543788 299624 543794
rect 187700 543730 187752 543736
rect 299572 543730 299624 543736
rect 299572 543652 299624 543658
rect 299572 543594 299624 543600
rect 187698 542600 187754 542609
rect 187698 542535 187754 542544
rect 187712 542434 187740 542535
rect 187700 542428 187752 542434
rect 187700 542370 187752 542376
rect 187790 540424 187846 540433
rect 187790 540359 187846 540368
rect 187698 539880 187754 539889
rect 187698 539815 187754 539824
rect 187712 539646 187740 539815
rect 187804 539714 187832 540359
rect 187792 539708 187844 539714
rect 187792 539650 187844 539656
rect 187700 539640 187752 539646
rect 187700 539582 187752 539588
rect 188342 537568 188398 537577
rect 188342 537503 188398 537512
rect 161388 458176 161440 458182
rect 161388 458118 161440 458124
rect 161400 457978 161428 458118
rect 161388 457972 161440 457978
rect 161388 457914 161440 457920
rect 176568 457700 176620 457706
rect 176568 457642 176620 457648
rect 175188 457632 175240 457638
rect 175188 457574 175240 457580
rect 172428 457564 172480 457570
rect 172428 457506 172480 457512
rect 171048 457428 171100 457434
rect 171048 457370 171100 457376
rect 149336 442876 149388 442882
rect 149336 442818 149388 442824
rect 150348 442876 150400 442882
rect 150348 442818 150400 442824
rect 147154 439878 147628 439906
rect 149348 439892 149376 442818
rect 153936 442808 153988 442814
rect 153936 442750 153988 442756
rect 151636 442196 151688 442202
rect 151636 442138 151688 442144
rect 151648 439892 151676 442138
rect 153948 439892 153976 442750
rect 156144 442740 156196 442746
rect 156144 442682 156196 442688
rect 156156 439892 156184 442682
rect 158444 442672 158496 442678
rect 158444 442614 158496 442620
rect 158456 439892 158484 442614
rect 160652 442604 160704 442610
rect 160652 442546 160704 442552
rect 160664 439892 160692 442546
rect 162950 442504 163006 442513
rect 162950 442439 163006 442448
rect 162964 439892 162992 442439
rect 165250 442368 165306 442377
rect 165250 442303 165306 442312
rect 165264 439892 165292 442303
rect 167458 442232 167514 442241
rect 167458 442167 167514 442176
rect 167472 439892 167500 442167
rect 171060 441998 171088 457370
rect 169760 441992 169812 441998
rect 169760 441934 169812 441940
rect 171048 441992 171100 441998
rect 171048 441934 171100 441940
rect 169772 439892 169800 441934
rect 172440 439906 172468 457506
rect 175200 442202 175228 457574
rect 174268 442196 174320 442202
rect 174268 442138 174320 442144
rect 175188 442196 175240 442202
rect 175188 442138 175240 442144
rect 172086 439878 172468 439906
rect 174280 439892 174308 442138
rect 176580 439892 176608 457642
rect 188356 442950 188384 537503
rect 299584 531350 299612 543594
rect 299572 531344 299624 531350
rect 299478 531312 299534 531321
rect 299664 531344 299716 531350
rect 299572 531286 299624 531292
rect 299662 531312 299664 531321
rect 299716 531312 299718 531321
rect 299478 531247 299534 531256
rect 299662 531247 299718 531256
rect 299492 521694 299520 531247
rect 299480 521688 299532 521694
rect 299480 521630 299532 521636
rect 299756 521688 299808 521694
rect 299756 521630 299808 521636
rect 299768 514706 299796 521630
rect 299676 514678 299796 514706
rect 299676 512009 299704 514678
rect 299478 512000 299534 512009
rect 299478 511935 299534 511944
rect 299662 512000 299718 512009
rect 299662 511935 299718 511944
rect 299492 502382 299520 511935
rect 299480 502376 299532 502382
rect 299480 502318 299532 502324
rect 299756 502376 299808 502382
rect 299756 502318 299808 502324
rect 299768 495394 299796 502318
rect 299676 495366 299796 495394
rect 299676 492658 299704 495366
rect 299480 492652 299532 492658
rect 299480 492594 299532 492600
rect 299664 492652 299716 492658
rect 299664 492594 299716 492600
rect 269118 484528 269174 484537
rect 269118 484463 269174 484472
rect 269132 484430 269160 484463
rect 269120 484424 269172 484430
rect 269120 484366 269172 484372
rect 299492 483041 299520 492594
rect 299478 483032 299534 483041
rect 299478 482967 299534 482976
rect 299754 483032 299810 483041
rect 299754 482967 299810 482976
rect 188986 480312 189042 480321
rect 188986 480247 189042 480256
rect 188894 478000 188950 478009
rect 188894 477935 188950 477944
rect 188908 460222 188936 477935
rect 188896 460216 188948 460222
rect 188896 460158 188948 460164
rect 188908 459542 188936 460158
rect 188896 459536 188948 459542
rect 188896 459478 188948 459484
rect 188344 442944 188396 442950
rect 188344 442886 188396 442892
rect 189000 442610 189028 480247
rect 299768 476082 299796 482967
rect 299676 476054 299796 476082
rect 299676 466478 299704 476054
rect 299664 466472 299716 466478
rect 299664 466414 299716 466420
rect 299756 466404 299808 466410
rect 299756 466346 299808 466352
rect 299768 463690 299796 466346
rect 299756 463684 299808 463690
rect 299756 463626 299808 463632
rect 299848 463684 299900 463690
rect 299848 463626 299900 463632
rect 215312 458182 215340 458213
rect 190460 458176 190512 458182
rect 200028 458176 200080 458182
rect 190460 458118 190512 458124
rect 193862 458144 193918 458153
rect 190472 457978 190500 458118
rect 209780 458176 209832 458182
rect 200028 458118 200080 458124
rect 200210 458144 200266 458153
rect 193862 458079 193918 458088
rect 190460 457972 190512 457978
rect 190460 457914 190512 457920
rect 193876 457502 193904 458079
rect 197358 458008 197414 458017
rect 197358 457943 197414 457952
rect 198738 458008 198794 458017
rect 200040 457978 200068 458118
rect 215300 458176 215352 458182
rect 210514 458144 210570 458153
rect 209832 458124 209912 458130
rect 209780 458118 209912 458124
rect 209792 458102 209912 458118
rect 200210 458079 200266 458088
rect 198738 457943 198794 457952
rect 200028 457972 200080 457978
rect 195978 457600 196034 457609
rect 195978 457535 196034 457544
rect 193864 457496 193916 457502
rect 193864 457438 193916 457444
rect 195992 457366 196020 457535
rect 197372 457434 197400 457943
rect 198752 457570 198780 457943
rect 200028 457914 200080 457920
rect 200224 457638 200252 458079
rect 207662 458008 207718 458017
rect 207662 457943 207718 457952
rect 208214 458008 208270 458017
rect 208214 457943 208270 457952
rect 201498 457736 201554 457745
rect 201498 457671 201500 457680
rect 201552 457671 201554 457680
rect 201500 457642 201552 457648
rect 200212 457632 200264 457638
rect 200212 457574 200264 457580
rect 198740 457564 198792 457570
rect 198740 457506 198792 457512
rect 197360 457428 197412 457434
rect 197360 457370 197412 457376
rect 195980 457360 196032 457366
rect 195980 457302 196032 457308
rect 202144 457360 202196 457366
rect 202144 457302 202196 457308
rect 206282 457328 206338 457337
rect 202156 457201 202184 457302
rect 206282 457263 206338 457272
rect 206834 457328 206890 457337
rect 206834 457263 206890 457272
rect 202142 457192 202198 457201
rect 202142 457127 202198 457136
rect 202786 457192 202842 457201
rect 202786 457127 202842 457136
rect 201500 442808 201552 442814
rect 201500 442750 201552 442756
rect 199200 442672 199252 442678
rect 199200 442614 199252 442620
rect 187884 442604 187936 442610
rect 187884 442546 187936 442552
rect 188988 442604 189040 442610
rect 188988 442546 189040 442552
rect 178776 442536 178828 442542
rect 178776 442478 178828 442484
rect 178788 439892 178816 442478
rect 181076 442468 181128 442474
rect 181076 442410 181128 442416
rect 181088 439892 181116 442410
rect 183376 442400 183428 442406
rect 183376 442342 183428 442348
rect 183388 439892 183416 442342
rect 185584 442332 185636 442338
rect 185584 442274 185636 442280
rect 185596 439892 185624 442274
rect 187896 439892 187924 442546
rect 194692 442400 194744 442406
rect 194692 442342 194744 442348
rect 190092 442264 190144 442270
rect 190092 442206 190144 442212
rect 192392 442264 192444 442270
rect 192392 442206 192444 442212
rect 190104 439892 190132 442206
rect 192404 439892 192432 442206
rect 194704 439892 194732 442342
rect 196900 442332 196952 442338
rect 196900 442274 196952 442280
rect 196912 439892 196940 442274
rect 199212 439892 199240 442614
rect 201512 439892 201540 442750
rect 202156 442270 202184 457127
rect 202800 442610 202828 457127
rect 204902 457056 204958 457065
rect 204902 456991 204958 457000
rect 205454 457056 205510 457065
rect 205454 456991 205510 457000
rect 203522 456920 203578 456929
rect 203522 456855 203578 456864
rect 204166 456920 204222 456929
rect 204166 456855 204222 456864
rect 203536 456822 203564 456855
rect 203524 456816 203576 456822
rect 203524 456758 203576 456764
rect 202788 442604 202840 442610
rect 202788 442546 202840 442552
rect 203536 442406 203564 456758
rect 204180 442542 204208 456855
rect 204168 442536 204220 442542
rect 204168 442478 204220 442484
rect 203524 442400 203576 442406
rect 203524 442342 203576 442348
rect 204916 442338 204944 456991
rect 205468 456890 205496 456991
rect 205546 456920 205602 456929
rect 205456 456884 205508 456890
rect 205546 456855 205602 456864
rect 205456 456826 205508 456832
rect 205560 442474 205588 456855
rect 206008 442944 206060 442950
rect 206008 442886 206060 442892
rect 205548 442468 205600 442474
rect 205548 442410 205600 442416
rect 204904 442332 204956 442338
rect 204904 442274 204956 442280
rect 202144 442264 202196 442270
rect 202144 442206 202196 442212
rect 203708 441924 203760 441930
rect 203708 441866 203760 441872
rect 203720 439892 203748 441866
rect 206020 439892 206048 442886
rect 206296 442678 206324 457263
rect 206848 456958 206876 457263
rect 206926 457192 206982 457201
rect 206926 457127 206982 457136
rect 206836 456952 206888 456958
rect 206836 456894 206888 456900
rect 206284 442672 206336 442678
rect 206284 442614 206336 442620
rect 206940 442406 206968 457127
rect 207676 442814 207704 457943
rect 208228 457910 208256 457943
rect 208216 457904 208268 457910
rect 208216 457846 208268 457852
rect 209686 457736 209742 457745
rect 207756 457700 207808 457706
rect 209686 457671 209688 457680
rect 207756 457642 207808 457648
rect 209740 457671 209742 457680
rect 209688 457642 209740 457648
rect 207768 442950 207796 457642
rect 209136 457632 209188 457638
rect 209136 457574 209188 457580
rect 209042 457464 209098 457473
rect 209042 457399 209044 457408
rect 209096 457399 209098 457408
rect 209044 457370 209096 457376
rect 208306 456920 208362 456929
rect 208306 456855 208362 456864
rect 207756 442944 207808 442950
rect 207756 442886 207808 442892
rect 208216 442944 208268 442950
rect 208216 442886 208268 442892
rect 207664 442808 207716 442814
rect 207664 442750 207716 442756
rect 206928 442400 206980 442406
rect 206928 442342 206980 442348
rect 208228 439892 208256 442886
rect 208320 442338 208348 456855
rect 208308 442332 208360 442338
rect 208308 442274 208360 442280
rect 209056 441930 209084 457370
rect 209148 442950 209176 457574
rect 209884 457298 209912 458102
rect 210514 458079 210570 458088
rect 212446 458144 212502 458153
rect 212446 458079 212502 458088
rect 213090 458144 213146 458153
rect 213090 458079 213146 458088
rect 214010 458144 214066 458153
rect 214010 458079 214066 458088
rect 215298 458144 215300 458153
rect 217232 458176 217284 458182
rect 215352 458144 215354 458153
rect 215298 458079 215354 458088
rect 216678 458144 216734 458153
rect 219348 458176 219400 458182
rect 217232 458118 217284 458124
rect 217598 458144 217654 458153
rect 216678 458079 216734 458088
rect 210528 457638 210556 458079
rect 210516 457632 210568 457638
rect 210516 457574 210568 457580
rect 212460 457570 212488 458079
rect 213104 457842 213132 458079
rect 213092 457836 213144 457842
rect 213092 457778 213144 457784
rect 212448 457564 212500 457570
rect 212448 457506 212500 457512
rect 212460 457366 212488 457506
rect 212448 457360 212500 457366
rect 212448 457302 212500 457308
rect 209780 457292 209832 457298
rect 209780 457234 209832 457240
rect 209872 457292 209924 457298
rect 209872 457234 209924 457240
rect 209686 456920 209742 456929
rect 209686 456855 209742 456864
rect 209136 442944 209188 442950
rect 209136 442886 209188 442892
rect 209700 442270 209728 456855
rect 209688 442264 209740 442270
rect 209688 442206 209740 442212
rect 209044 441924 209096 441930
rect 209044 441866 209096 441872
rect 209792 440450 209820 457234
rect 212540 457224 212592 457230
rect 210974 457192 211030 457201
rect 212540 457166 212592 457172
rect 210974 457127 211030 457136
rect 210988 441658 211016 457127
rect 211066 456920 211122 456929
rect 211066 456855 211122 456864
rect 212446 456920 212502 456929
rect 212446 456855 212502 456864
rect 211080 441794 211108 456855
rect 211068 441788 211120 441794
rect 211068 441730 211120 441736
rect 212460 441726 212488 456855
rect 212448 441720 212500 441726
rect 212448 441662 212500 441668
rect 210976 441652 211028 441658
rect 210976 441594 211028 441600
rect 209792 440422 210188 440450
rect 210160 439906 210188 440422
rect 212552 439906 212580 457166
rect 213104 456822 213132 457778
rect 214024 457774 214052 458079
rect 214012 457768 214064 457774
rect 214012 457710 214064 457716
rect 213920 457156 213972 457162
rect 213920 457098 213972 457104
rect 213826 456920 213882 456929
rect 213826 456855 213882 456864
rect 213092 456816 213144 456822
rect 213092 456758 213144 456764
rect 213840 441862 213868 456855
rect 213828 441856 213880 441862
rect 213828 441798 213880 441804
rect 213932 440450 213960 457098
rect 214024 456890 214052 457710
rect 215206 457192 215262 457201
rect 215206 457127 215208 457136
rect 215260 457127 215262 457136
rect 215208 457098 215260 457104
rect 215312 456958 215340 458079
rect 216692 457910 216720 458079
rect 217244 457910 217272 458118
rect 217598 458079 217654 458088
rect 218886 458144 218942 458153
rect 226340 458176 226392 458182
rect 219348 458118 219400 458124
rect 220174 458144 220230 458153
rect 218886 458079 218942 458088
rect 216680 457904 216732 457910
rect 216680 457846 216732 457852
rect 217140 457904 217192 457910
rect 217140 457846 217192 457852
rect 217232 457904 217284 457910
rect 217232 457846 217284 457852
rect 216586 457464 216642 457473
rect 217152 457434 217180 457846
rect 216586 457399 216642 457408
rect 217140 457428 217192 457434
rect 215300 456952 215352 456958
rect 215300 456894 215352 456900
rect 216600 456890 216628 457399
rect 217140 457370 217192 457376
rect 217612 457366 217640 458079
rect 218900 457706 218928 458079
rect 218888 457700 218940 457706
rect 218888 457642 218940 457648
rect 217600 457360 217652 457366
rect 217600 457302 217652 457308
rect 219360 457298 219388 458118
rect 220174 458079 220230 458088
rect 221370 458144 221426 458153
rect 221370 458079 221426 458088
rect 222566 458144 222622 458153
rect 223670 458144 223726 458153
rect 222566 458079 222622 458088
rect 223580 458108 223632 458114
rect 220188 457638 220216 458079
rect 220820 458040 220872 458046
rect 220820 457982 220872 457988
rect 220176 457632 220228 457638
rect 220176 457574 220228 457580
rect 219348 457292 219400 457298
rect 219348 457234 219400 457240
rect 217966 457192 218022 457201
rect 217966 457127 218022 457136
rect 220726 457192 220782 457201
rect 220726 457127 220782 457136
rect 216680 457088 216732 457094
rect 216680 457030 216732 457036
rect 214012 456884 214064 456890
rect 214012 456826 214064 456832
rect 216588 456884 216640 456890
rect 216588 456826 216640 456832
rect 216692 440450 216720 457030
rect 217874 456920 217930 456929
rect 217874 456855 217930 456864
rect 217888 441998 217916 456855
rect 217980 456822 218008 457127
rect 219440 457020 219492 457026
rect 219440 456962 219492 456968
rect 219346 456920 219402 456929
rect 219346 456855 219402 456864
rect 217968 456816 218020 456822
rect 217968 456758 218020 456764
rect 217876 441992 217928 441998
rect 217876 441934 217928 441940
rect 219360 441930 219388 456855
rect 219348 441924 219400 441930
rect 219348 441866 219400 441872
rect 213932 440422 214788 440450
rect 216692 440422 216996 440450
rect 214760 439906 214788 440422
rect 216968 439906 216996 440422
rect 219452 439906 219480 456962
rect 220740 442134 220768 457127
rect 220728 442128 220780 442134
rect 220728 442070 220780 442076
rect 220832 440450 220860 457982
rect 221384 457570 221412 458079
rect 222580 457842 222608 458079
rect 223670 458079 223672 458088
rect 223580 458050 223632 458056
rect 223724 458079 223726 458088
rect 224314 458144 224370 458153
rect 224314 458079 224370 458088
rect 225878 458144 225934 458153
rect 226340 458118 226392 458124
rect 227166 458144 227222 458153
rect 225878 458079 225934 458088
rect 223672 458050 223724 458056
rect 222568 457836 222620 457842
rect 222568 457778 222620 457784
rect 221372 457564 221424 457570
rect 221372 457506 221424 457512
rect 222106 456920 222162 456929
rect 222106 456855 222162 456864
rect 223486 456920 223542 456929
rect 223486 456855 223542 456864
rect 222120 442066 222148 456855
rect 223500 442202 223528 456855
rect 223488 442196 223540 442202
rect 223488 442138 223540 442144
rect 222108 442060 222160 442066
rect 222108 442002 222160 442008
rect 223592 440450 223620 458050
rect 223684 457774 223712 458050
rect 224328 458046 224356 458079
rect 224316 458040 224368 458046
rect 224316 457982 224368 457988
rect 224328 457910 224356 457982
rect 225892 457978 225920 458079
rect 224960 457972 225012 457978
rect 224960 457914 225012 457920
rect 225880 457972 225932 457978
rect 225880 457914 225932 457920
rect 224316 457904 224368 457910
rect 224316 457846 224368 457852
rect 223672 457768 223724 457774
rect 223672 457710 223724 457716
rect 224972 457434 225000 457914
rect 224960 457428 225012 457434
rect 224960 457370 225012 457376
rect 226246 457056 226302 457065
rect 226246 456991 226302 457000
rect 224866 456920 224922 456929
rect 224866 456855 224922 456864
rect 226154 456920 226210 456929
rect 226154 456855 226210 456864
rect 224880 442950 224908 456855
rect 224868 442944 224920 442950
rect 224868 442886 224920 442892
rect 226168 442814 226196 456855
rect 226260 442882 226288 456991
rect 226248 442876 226300 442882
rect 226248 442818 226300 442824
rect 226156 442808 226208 442814
rect 226156 442750 226208 442756
rect 220832 440422 221596 440450
rect 223592 440422 223804 440450
rect 221568 439906 221596 440422
rect 223776 439906 223804 440422
rect 210160 439878 210542 439906
rect 212552 439878 212842 439906
rect 214760 439878 215050 439906
rect 216968 439878 217350 439906
rect 219452 439878 219558 439906
rect 221568 439878 221858 439906
rect 223776 439878 224158 439906
rect 226352 439892 226380 458118
rect 227166 458079 227222 458088
rect 228362 458144 228418 458153
rect 228362 458079 228418 458088
rect 229558 458144 229614 458153
rect 229558 458079 229614 458088
rect 231858 458144 231914 458153
rect 231858 458079 231860 458088
rect 227180 457774 227208 458079
rect 226432 457768 226484 457774
rect 226432 457710 226484 457716
rect 227168 457768 227220 457774
rect 227168 457710 227220 457716
rect 226444 457366 226472 457710
rect 228376 457706 228404 458079
rect 228364 457700 228416 457706
rect 228364 457642 228416 457648
rect 229572 457638 229600 458079
rect 231912 458079 231914 458088
rect 233238 458144 233294 458153
rect 233238 458079 233294 458088
rect 231860 458050 231912 458056
rect 233252 458046 233280 458079
rect 233240 458040 233292 458046
rect 233240 457982 233292 457988
rect 234618 458008 234674 458017
rect 234618 457943 234620 457952
rect 234672 457943 234674 457952
rect 234620 457914 234672 457920
rect 231858 457872 231914 457881
rect 231858 457807 231860 457816
rect 231912 457807 231914 457816
rect 235998 457872 236054 457881
rect 235998 457807 236054 457816
rect 231860 457778 231912 457784
rect 236012 457774 236040 457807
rect 236000 457768 236052 457774
rect 236000 457710 236052 457716
rect 237378 457736 237434 457745
rect 237378 457671 237380 457680
rect 237432 457671 237434 457680
rect 238758 457736 238814 457745
rect 238758 457671 238814 457680
rect 237380 457642 237432 457648
rect 238772 457638 238800 457671
rect 229560 457632 229612 457638
rect 238760 457632 238812 457638
rect 229560 457574 229612 457580
rect 230478 457600 230534 457609
rect 238760 457574 238812 457580
rect 230478 457535 230480 457544
rect 230532 457535 230534 457544
rect 230480 457506 230532 457512
rect 226432 457360 226484 457366
rect 226432 457302 226484 457308
rect 246304 457156 246356 457162
rect 246304 457098 246356 457104
rect 233054 457056 233110 457065
rect 233054 456991 233110 457000
rect 227626 456920 227682 456929
rect 227626 456855 227682 456864
rect 229006 456920 229062 456929
rect 229006 456855 229062 456864
rect 230386 456920 230442 456929
rect 230386 456855 230442 456864
rect 231766 456920 231822 456929
rect 231766 456855 231822 456864
rect 227640 442746 227668 456855
rect 227628 442740 227680 442746
rect 227628 442682 227680 442688
rect 229020 442678 229048 456855
rect 229008 442672 229060 442678
rect 229008 442614 229060 442620
rect 230400 442610 230428 456855
rect 228640 442604 228692 442610
rect 228640 442546 228692 442552
rect 230388 442604 230440 442610
rect 230388 442546 230440 442552
rect 228652 439892 228680 442546
rect 231780 442542 231808 456855
rect 230848 442536 230900 442542
rect 230848 442478 230900 442484
rect 231768 442536 231820 442542
rect 231768 442478 231820 442484
rect 230860 439892 230888 442478
rect 233068 442474 233096 456991
rect 233146 456920 233202 456929
rect 233146 456855 233202 456864
rect 234526 456920 234582 456929
rect 234526 456855 234582 456864
rect 235906 456920 235962 456929
rect 235906 456855 235962 456864
rect 237286 456920 237342 456929
rect 237286 456855 237342 456864
rect 238666 456920 238722 456929
rect 238666 456855 238722 456864
rect 240046 456920 240102 456929
rect 240046 456855 240102 456864
rect 244924 456884 244976 456890
rect 233160 442513 233188 456855
rect 233146 442504 233202 442513
rect 232780 442468 232832 442474
rect 232780 442410 232832 442416
rect 233056 442468 233108 442474
rect 233146 442439 233202 442448
rect 233056 442410 233108 442416
rect 232792 439906 232820 442410
rect 234540 442377 234568 456855
rect 235920 442406 235948 456855
rect 235448 442400 235500 442406
rect 234526 442368 234582 442377
rect 235448 442342 235500 442348
rect 235908 442400 235960 442406
rect 235908 442342 235960 442348
rect 234526 442303 234582 442312
rect 232792 439878 233174 439906
rect 235460 439892 235488 442342
rect 237300 442241 237328 456855
rect 238680 442338 238708 456855
rect 237656 442332 237708 442338
rect 237656 442274 237708 442280
rect 238668 442332 238720 442338
rect 238668 442274 238720 442280
rect 237286 442232 237342 442241
rect 237286 442167 237342 442176
rect 237668 439892 237696 442274
rect 239956 442264 240008 442270
rect 239956 442206 240008 442212
rect 239968 439892 239996 442206
rect 240060 441697 240088 456855
rect 244924 456826 244976 456832
rect 242164 456816 242216 456822
rect 242164 456758 242216 456764
rect 242176 446434 242204 456758
rect 242176 446406 242388 446434
rect 242360 443290 242388 446406
rect 242348 443284 242400 443290
rect 242348 443226 242400 443232
rect 242072 442264 242124 442270
rect 242072 442206 242124 442212
rect 242084 441726 242112 442206
rect 244936 441862 244964 456826
rect 245108 443284 245160 443290
rect 245108 443226 245160 443232
rect 244924 441856 244976 441862
rect 244924 441798 244976 441804
rect 244464 441788 244516 441794
rect 244464 441730 244516 441736
rect 242072 441720 242124 441726
rect 240046 441688 240102 441697
rect 242072 441662 242124 441668
rect 240046 441623 240102 441632
rect 242256 441652 242308 441658
rect 242256 441594 242308 441600
rect 242268 439892 242296 441594
rect 244476 439892 244504 441730
rect 245120 441658 245148 443226
rect 246316 442270 246344 457098
rect 299860 456822 299888 463626
rect 299848 456816 299900 456822
rect 299848 456758 299900 456764
rect 299756 456748 299808 456754
rect 299756 456690 299808 456696
rect 299768 454050 299796 456690
rect 299768 454022 299888 454050
rect 299860 444446 299888 454022
rect 299664 444440 299716 444446
rect 299664 444382 299716 444388
rect 299848 444440 299900 444446
rect 299848 444382 299900 444388
rect 269396 442944 269448 442950
rect 269396 442886 269448 442892
rect 246212 442264 246264 442270
rect 246212 442206 246264 442212
rect 246304 442264 246356 442270
rect 246304 442206 246356 442212
rect 251272 442264 251324 442270
rect 251272 442206 251324 442212
rect 251364 442264 251416 442270
rect 251364 442206 251416 442212
rect 245108 441652 245160 441658
rect 245108 441594 245160 441600
rect 246224 439906 246252 442206
rect 248604 441788 248656 441794
rect 248604 441730 248656 441736
rect 248696 441788 248748 441794
rect 248696 441730 248748 441736
rect 248616 439906 248644 441730
rect 248708 441697 248736 441730
rect 248694 441688 248750 441697
rect 248694 441623 248750 441632
rect 246224 439878 246790 439906
rect 248616 439878 248998 439906
rect 251284 439892 251312 442206
rect 251376 441794 251404 442206
rect 267096 442196 267148 442202
rect 267096 442138 267148 442144
rect 262588 442128 262640 442134
rect 262588 442070 262640 442076
rect 258080 441992 258132 441998
rect 258080 441934 258132 441940
rect 253572 441856 253624 441862
rect 253572 441798 253624 441804
rect 251364 441788 251416 441794
rect 251364 441730 251416 441736
rect 253584 439892 253612 441798
rect 255780 441652 255832 441658
rect 255780 441594 255832 441600
rect 255792 439892 255820 441594
rect 258092 439892 258120 441934
rect 260288 441924 260340 441930
rect 260288 441866 260340 441872
rect 260300 439892 260328 441866
rect 262600 439892 262628 442070
rect 264888 442060 264940 442066
rect 264888 442002 264940 442008
rect 264900 439892 264928 442002
rect 267108 439892 267136 442138
rect 269408 439892 269436 442886
rect 271696 442876 271748 442882
rect 271696 442818 271748 442824
rect 271708 439892 271736 442818
rect 273904 442808 273956 442814
rect 273904 442750 273956 442756
rect 273916 439892 273944 442750
rect 276204 442740 276256 442746
rect 276204 442682 276256 442688
rect 276216 439892 276244 442682
rect 278412 442672 278464 442678
rect 278412 442614 278464 442620
rect 278424 439892 278452 442614
rect 280712 442604 280764 442610
rect 280712 442546 280764 442552
rect 280724 439892 280752 442546
rect 283012 442536 283064 442542
rect 283012 442478 283064 442484
rect 287518 442504 287574 442513
rect 283024 439892 283052 442478
rect 285220 442468 285272 442474
rect 287518 442439 287574 442448
rect 285220 442410 285272 442416
rect 285232 439892 285260 442410
rect 287532 439892 287560 442439
rect 292028 442400 292080 442406
rect 289726 442368 289782 442377
rect 292028 442342 292080 442348
rect 289726 442303 289782 442312
rect 289740 439892 289768 442303
rect 292040 439892 292068 442342
rect 296536 442332 296588 442338
rect 296536 442274 296588 442280
rect 294326 442232 294382 442241
rect 294326 442167 294382 442176
rect 294340 439892 294368 442167
rect 296548 439892 296576 442274
rect 298836 442264 298888 442270
rect 298836 442206 298888 442212
rect 298848 439892 298876 442206
rect 65642 439742 66208 439770
rect 72450 439742 73108 439770
rect 136456 439816 136508 439822
rect 136456 439758 136508 439764
rect 299676 439754 299704 444382
rect 299664 439748 299716 439754
rect 299664 439690 299716 439696
rect 302252 203425 302280 549238
rect 389376 547890 389404 553386
rect 429304 550662 429332 560186
rect 507860 554056 507912 554062
rect 507860 553998 507912 554004
rect 513380 554056 513432 554062
rect 513380 553998 513432 554004
rect 507872 553489 507900 553998
rect 513392 553489 513420 553998
rect 507858 553480 507914 553489
rect 507858 553415 507860 553424
rect 507912 553415 507914 553424
rect 513378 553480 513434 553489
rect 558932 553450 558960 560238
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 513378 553415 513434 553424
rect 558920 553444 558972 553450
rect 507860 553386 507912 553392
rect 558920 553386 558972 553392
rect 507872 553355 507900 553386
rect 559012 553376 559064 553382
rect 559012 553318 559064 553324
rect 518898 550760 518954 550769
rect 518898 550695 518954 550704
rect 429292 550656 429344 550662
rect 429292 550598 429344 550604
rect 429568 550656 429620 550662
rect 429568 550598 429620 550604
rect 389192 547862 389404 547890
rect 305826 546544 305882 546553
rect 305826 546479 305882 546488
rect 304448 545148 304500 545154
rect 304448 545090 304500 545096
rect 304356 542428 304408 542434
rect 304356 542370 304408 542376
rect 304264 539640 304316 539646
rect 304264 539582 304316 539588
rect 302884 484424 302936 484430
rect 302884 484366 302936 484372
rect 302896 459474 302924 484366
rect 302976 477556 303028 477562
rect 302976 477498 303028 477504
rect 302988 460222 303016 477498
rect 302976 460216 303028 460222
rect 302976 460158 303028 460164
rect 302988 459542 303016 460158
rect 302976 459536 303028 459542
rect 302976 459478 303028 459484
rect 302884 459468 302936 459474
rect 302884 459410 302936 459416
rect 302792 437436 302844 437442
rect 302792 437378 302844 437384
rect 302804 436801 302832 437378
rect 302790 436792 302846 436801
rect 302790 436727 302846 436736
rect 302792 434716 302844 434722
rect 302792 434658 302844 434664
rect 302804 434625 302832 434658
rect 302790 434616 302846 434625
rect 302790 434551 302846 434560
rect 302792 433288 302844 433294
rect 302792 433230 302844 433236
rect 302804 432449 302832 433230
rect 302790 432440 302846 432449
rect 302790 432375 302846 432384
rect 302792 430568 302844 430574
rect 302792 430510 302844 430516
rect 302804 430273 302832 430510
rect 302790 430264 302846 430273
rect 302790 430199 302846 430208
rect 302792 429140 302844 429146
rect 302792 429082 302844 429088
rect 302804 427961 302832 429082
rect 302790 427952 302846 427961
rect 302790 427887 302846 427896
rect 302792 426420 302844 426426
rect 302792 426362 302844 426368
rect 302804 425785 302832 426362
rect 302790 425776 302846 425785
rect 302790 425711 302846 425720
rect 302792 423632 302844 423638
rect 302790 423600 302792 423609
rect 302844 423600 302846 423609
rect 302790 423535 302846 423544
rect 302792 422272 302844 422278
rect 302792 422214 302844 422220
rect 302804 421433 302832 422214
rect 302790 421424 302846 421433
rect 302790 421359 302846 421368
rect 302792 419484 302844 419490
rect 302792 419426 302844 419432
rect 302804 419257 302832 419426
rect 302790 419248 302846 419257
rect 302790 419183 302846 419192
rect 302792 418124 302844 418130
rect 302792 418066 302844 418072
rect 302804 416945 302832 418066
rect 302790 416936 302846 416945
rect 302790 416871 302846 416880
rect 302792 415404 302844 415410
rect 302792 415346 302844 415352
rect 302804 414769 302832 415346
rect 302790 414760 302846 414769
rect 302790 414695 302846 414704
rect 302792 412616 302844 412622
rect 302790 412584 302792 412593
rect 302844 412584 302846 412593
rect 302790 412519 302846 412528
rect 302792 411256 302844 411262
rect 302792 411198 302844 411204
rect 302804 410417 302832 411198
rect 302790 410408 302846 410417
rect 302790 410343 302846 410352
rect 302792 408468 302844 408474
rect 302792 408410 302844 408416
rect 302804 408241 302832 408410
rect 302790 408232 302846 408241
rect 302790 408167 302846 408176
rect 302792 407108 302844 407114
rect 302792 407050 302844 407056
rect 302804 405929 302832 407050
rect 302790 405920 302846 405929
rect 302790 405855 302846 405864
rect 302700 404320 302752 404326
rect 302700 404262 302752 404268
rect 302712 403753 302740 404262
rect 302698 403744 302754 403753
rect 302698 403679 302754 403688
rect 302792 401600 302844 401606
rect 302790 401568 302792 401577
rect 302844 401568 302846 401577
rect 302790 401503 302846 401512
rect 302792 400172 302844 400178
rect 302792 400114 302844 400120
rect 302804 399401 302832 400114
rect 302790 399392 302846 399401
rect 302790 399327 302846 399336
rect 302792 397452 302844 397458
rect 302792 397394 302844 397400
rect 302804 397225 302832 397394
rect 302790 397216 302846 397225
rect 302790 397151 302846 397160
rect 302516 396024 302568 396030
rect 302516 395966 302568 395972
rect 302528 394913 302556 395966
rect 302514 394904 302570 394913
rect 302514 394839 302570 394848
rect 302700 393304 302752 393310
rect 302700 393246 302752 393252
rect 302712 392737 302740 393246
rect 302698 392728 302754 392737
rect 302698 392663 302754 392672
rect 302790 390552 302846 390561
rect 302790 390487 302792 390496
rect 302844 390487 302846 390496
rect 302792 390458 302844 390464
rect 302792 389156 302844 389162
rect 302792 389098 302844 389104
rect 302804 388385 302832 389098
rect 302790 388376 302846 388385
rect 302790 388311 302846 388320
rect 302516 386368 302568 386374
rect 302516 386310 302568 386316
rect 302528 386209 302556 386310
rect 302514 386200 302570 386209
rect 302514 386135 302570 386144
rect 302516 385008 302568 385014
rect 302516 384950 302568 384956
rect 302528 383897 302556 384950
rect 302514 383888 302570 383897
rect 302514 383823 302570 383832
rect 302792 382220 302844 382226
rect 302792 382162 302844 382168
rect 302804 381721 302832 382162
rect 302790 381712 302846 381721
rect 302790 381647 302846 381656
rect 302608 380860 302660 380866
rect 302608 380802 302660 380808
rect 302620 379545 302648 380802
rect 302606 379536 302662 379545
rect 302606 379471 302662 379480
rect 302792 378140 302844 378146
rect 302792 378082 302844 378088
rect 302804 377369 302832 378082
rect 302790 377360 302846 377369
rect 302790 377295 302846 377304
rect 302792 375352 302844 375358
rect 302792 375294 302844 375300
rect 302804 375193 302832 375294
rect 302790 375184 302846 375193
rect 302790 375119 302846 375128
rect 302792 373992 302844 373998
rect 302792 373934 302844 373940
rect 302804 373017 302832 373934
rect 302790 373008 302846 373017
rect 302790 372943 302846 372952
rect 302332 371204 302384 371210
rect 302332 371146 302384 371152
rect 302344 370705 302372 371146
rect 302330 370696 302386 370705
rect 302330 370631 302386 370640
rect 302608 369844 302660 369850
rect 302608 369786 302660 369792
rect 302620 368529 302648 369786
rect 302606 368520 302662 368529
rect 302606 368455 302662 368464
rect 302792 367056 302844 367062
rect 302792 366998 302844 367004
rect 302804 366353 302832 366998
rect 302790 366344 302846 366353
rect 302790 366279 302846 366288
rect 302516 364336 302568 364342
rect 302516 364278 302568 364284
rect 302528 364177 302556 364278
rect 302514 364168 302570 364177
rect 302514 364103 302570 364112
rect 302424 362908 302476 362914
rect 302424 362850 302476 362856
rect 302436 362001 302464 362850
rect 302422 361992 302478 362001
rect 302422 361927 302478 361936
rect 302332 360188 302384 360194
rect 302332 360130 302384 360136
rect 302344 359689 302372 360130
rect 302330 359680 302386 359689
rect 302330 359615 302386 359624
rect 302516 358760 302568 358766
rect 302516 358702 302568 358708
rect 302528 357513 302556 358702
rect 302514 357504 302570 357513
rect 302514 357439 302570 357448
rect 302792 356040 302844 356046
rect 302792 355982 302844 355988
rect 302804 355337 302832 355982
rect 302790 355328 302846 355337
rect 302790 355263 302846 355272
rect 302792 353252 302844 353258
rect 302792 353194 302844 353200
rect 302804 353161 302832 353194
rect 302790 353152 302846 353161
rect 302790 353087 302846 353096
rect 302424 351892 302476 351898
rect 302424 351834 302476 351840
rect 302436 350985 302464 351834
rect 302422 350976 302478 350985
rect 302422 350911 302478 350920
rect 302700 349104 302752 349110
rect 302700 349046 302752 349052
rect 302712 348673 302740 349046
rect 302698 348664 302754 348673
rect 302698 348599 302754 348608
rect 302516 347744 302568 347750
rect 302516 347686 302568 347692
rect 302528 346497 302556 347686
rect 302514 346488 302570 346497
rect 302514 346423 302570 346432
rect 302792 345024 302844 345030
rect 302792 344966 302844 344972
rect 302804 344321 302832 344966
rect 302790 344312 302846 344321
rect 302790 344247 302846 344256
rect 302792 342236 302844 342242
rect 302792 342178 302844 342184
rect 302804 342145 302832 342178
rect 302790 342136 302846 342145
rect 302790 342071 302846 342080
rect 302424 340876 302476 340882
rect 302424 340818 302476 340824
rect 302436 339969 302464 340818
rect 302422 339960 302478 339969
rect 302422 339895 302478 339904
rect 302700 338088 302752 338094
rect 302700 338030 302752 338036
rect 302712 337657 302740 338030
rect 302698 337648 302754 337657
rect 302698 337583 302754 337592
rect 302516 336728 302568 336734
rect 302516 336670 302568 336676
rect 302528 335481 302556 336670
rect 302514 335472 302570 335481
rect 302514 335407 302570 335416
rect 302792 333940 302844 333946
rect 302792 333882 302844 333888
rect 302804 333305 302832 333882
rect 302790 333296 302846 333305
rect 302790 333231 302846 333240
rect 302516 331152 302568 331158
rect 302514 331120 302516 331129
rect 302568 331120 302570 331129
rect 302514 331055 302570 331064
rect 302332 329452 302384 329458
rect 302332 329394 302384 329400
rect 302344 328953 302372 329394
rect 302330 328944 302386 328953
rect 302330 328879 302386 328888
rect 302516 326936 302568 326942
rect 302516 326878 302568 326884
rect 302528 326641 302556 326878
rect 302514 326632 302570 326641
rect 302514 326567 302570 326576
rect 302332 324488 302384 324494
rect 302330 324456 302332 324465
rect 302384 324456 302386 324465
rect 302330 324391 302386 324400
rect 302332 322720 302384 322726
rect 302332 322662 302384 322668
rect 302344 322289 302372 322662
rect 302330 322280 302386 322289
rect 302330 322215 302386 322224
rect 302332 320136 302384 320142
rect 302330 320104 302332 320113
rect 302384 320104 302386 320113
rect 302330 320039 302386 320048
rect 302700 318368 302752 318374
rect 302700 318310 302752 318316
rect 302712 317937 302740 318310
rect 302698 317928 302754 317937
rect 302698 317863 302754 317872
rect 302792 315988 302844 315994
rect 302792 315930 302844 315936
rect 302804 315761 302832 315930
rect 302790 315752 302846 315761
rect 302790 315687 302846 315696
rect 302792 314628 302844 314634
rect 302792 314570 302844 314576
rect 302804 313449 302832 314570
rect 302790 313440 302846 313449
rect 302790 313375 302846 313384
rect 302700 311840 302752 311846
rect 302700 311782 302752 311788
rect 302712 311273 302740 311782
rect 302698 311264 302754 311273
rect 302698 311199 302754 311208
rect 302792 309120 302844 309126
rect 302790 309088 302792 309097
rect 302844 309088 302846 309097
rect 302790 309023 302846 309032
rect 302792 307760 302844 307766
rect 302792 307702 302844 307708
rect 302804 306921 302832 307702
rect 302790 306912 302846 306921
rect 302790 306847 302846 306856
rect 302792 304972 302844 304978
rect 302792 304914 302844 304920
rect 302804 304745 302832 304914
rect 302790 304736 302846 304745
rect 302790 304671 302846 304680
rect 302792 303612 302844 303618
rect 302792 303554 302844 303560
rect 302804 302433 302832 303554
rect 302790 302424 302846 302433
rect 302790 302359 302846 302368
rect 302700 300824 302752 300830
rect 302700 300766 302752 300772
rect 302712 300257 302740 300766
rect 302698 300248 302754 300257
rect 302698 300183 302754 300192
rect 302792 298104 302844 298110
rect 302790 298072 302792 298081
rect 302844 298072 302846 298081
rect 302790 298007 302846 298016
rect 302608 295928 302660 295934
rect 302606 295896 302608 295905
rect 302660 295896 302662 295905
rect 302606 295831 302662 295840
rect 302792 293956 302844 293962
rect 302792 293898 302844 293904
rect 302804 293729 302832 293898
rect 302790 293720 302846 293729
rect 302790 293655 302846 293664
rect 302516 292528 302568 292534
rect 302516 292470 302568 292476
rect 302528 291417 302556 292470
rect 302514 291408 302570 291417
rect 302514 291343 302570 291352
rect 302700 289808 302752 289814
rect 302700 289750 302752 289756
rect 302712 289241 302740 289750
rect 302698 289232 302754 289241
rect 302698 289167 302754 289176
rect 302790 287056 302846 287065
rect 302790 286991 302792 287000
rect 302844 286991 302846 287000
rect 302792 286962 302844 286968
rect 302700 285320 302752 285326
rect 302700 285262 302752 285268
rect 302712 284889 302740 285262
rect 302698 284880 302754 284889
rect 302698 284815 302754 284824
rect 302516 282872 302568 282878
rect 302516 282814 302568 282820
rect 302528 282713 302556 282814
rect 302514 282704 302570 282713
rect 302514 282639 302570 282648
rect 302516 281512 302568 281518
rect 302516 281454 302568 281460
rect 302528 280401 302556 281454
rect 302514 280392 302570 280401
rect 302514 280327 302570 280336
rect 302332 278724 302384 278730
rect 302332 278666 302384 278672
rect 302344 278225 302372 278666
rect 302330 278216 302386 278225
rect 302330 278151 302386 278160
rect 302608 277364 302660 277370
rect 302608 277306 302660 277312
rect 302620 276049 302648 277306
rect 302606 276040 302662 276049
rect 302606 275975 302662 275984
rect 302792 274644 302844 274650
rect 302792 274586 302844 274592
rect 302804 273873 302832 274586
rect 302790 273864 302846 273873
rect 302790 273799 302846 273808
rect 302516 271856 302568 271862
rect 302516 271798 302568 271804
rect 302528 271697 302556 271798
rect 302514 271688 302570 271697
rect 302514 271623 302570 271632
rect 302516 270496 302568 270502
rect 302516 270438 302568 270444
rect 302528 269385 302556 270438
rect 302514 269376 302570 269385
rect 302514 269311 302570 269320
rect 302332 267708 302384 267714
rect 302332 267650 302384 267656
rect 302344 267209 302372 267650
rect 302330 267200 302386 267209
rect 302330 267135 302386 267144
rect 302608 266348 302660 266354
rect 302608 266290 302660 266296
rect 302620 265033 302648 266290
rect 302606 265024 302662 265033
rect 302606 264959 302662 264968
rect 302792 263560 302844 263566
rect 302792 263502 302844 263508
rect 302804 262857 302832 263502
rect 302790 262848 302846 262857
rect 302790 262783 302846 262792
rect 302516 260840 302568 260846
rect 302516 260782 302568 260788
rect 302528 260681 302556 260782
rect 302514 260672 302570 260681
rect 302514 260607 302570 260616
rect 302424 259412 302476 259418
rect 302424 259354 302476 259360
rect 302436 258505 302464 259354
rect 302422 258496 302478 258505
rect 302422 258431 302478 258440
rect 302332 256692 302384 256698
rect 302332 256634 302384 256640
rect 302344 256193 302372 256634
rect 302330 256184 302386 256193
rect 302330 256119 302386 256128
rect 302516 255264 302568 255270
rect 302516 255206 302568 255212
rect 302528 254017 302556 255206
rect 302514 254008 302570 254017
rect 302514 253943 302570 253952
rect 302792 252544 302844 252550
rect 302792 252486 302844 252492
rect 302804 251841 302832 252486
rect 302790 251832 302846 251841
rect 302790 251767 302846 251776
rect 302792 249756 302844 249762
rect 302792 249698 302844 249704
rect 302804 249665 302832 249698
rect 302790 249656 302846 249665
rect 302790 249591 302846 249600
rect 302424 248396 302476 248402
rect 302424 248338 302476 248344
rect 302436 247489 302464 248338
rect 302422 247480 302478 247489
rect 302422 247415 302478 247424
rect 302700 245608 302752 245614
rect 302700 245550 302752 245556
rect 302712 245177 302740 245550
rect 302698 245168 302754 245177
rect 302698 245103 302754 245112
rect 302516 244248 302568 244254
rect 302516 244190 302568 244196
rect 302528 243001 302556 244190
rect 302514 242992 302570 243001
rect 302514 242927 302570 242936
rect 302792 241460 302844 241466
rect 302792 241402 302844 241408
rect 302804 240825 302832 241402
rect 302790 240816 302846 240825
rect 302790 240751 302846 240760
rect 302792 238740 302844 238746
rect 302792 238682 302844 238688
rect 302804 238649 302832 238682
rect 302790 238640 302846 238649
rect 302790 238575 302846 238584
rect 302424 237380 302476 237386
rect 302424 237322 302476 237328
rect 302436 236473 302464 237322
rect 302422 236464 302478 236473
rect 302422 236399 302478 236408
rect 302700 234592 302752 234598
rect 302700 234534 302752 234540
rect 302712 234161 302740 234534
rect 302698 234152 302754 234161
rect 302698 234087 302754 234096
rect 302516 233232 302568 233238
rect 302516 233174 302568 233180
rect 302528 231985 302556 233174
rect 302514 231976 302570 231985
rect 302514 231911 302570 231920
rect 302792 230444 302844 230450
rect 302792 230386 302844 230392
rect 302804 229809 302832 230386
rect 302790 229800 302846 229809
rect 302790 229735 302846 229744
rect 302792 227724 302844 227730
rect 302792 227666 302844 227672
rect 302804 227633 302832 227666
rect 302790 227624 302846 227633
rect 302790 227559 302846 227568
rect 302792 226296 302844 226302
rect 302792 226238 302844 226244
rect 302804 225457 302832 226238
rect 302790 225448 302846 225457
rect 302790 225383 302846 225392
rect 302700 223576 302752 223582
rect 302700 223518 302752 223524
rect 302712 223145 302740 223518
rect 302698 223136 302754 223145
rect 302698 223071 302754 223080
rect 302792 222148 302844 222154
rect 302792 222090 302844 222096
rect 302804 220969 302832 222090
rect 302790 220960 302846 220969
rect 302790 220895 302846 220904
rect 302792 219428 302844 219434
rect 302792 219370 302844 219376
rect 302804 218793 302832 219370
rect 302790 218784 302846 218793
rect 302790 218719 302846 218728
rect 302792 216640 302844 216646
rect 302790 216608 302792 216617
rect 302844 216608 302846 216617
rect 302790 216543 302846 216552
rect 302792 215280 302844 215286
rect 302792 215222 302844 215228
rect 302804 214441 302832 215222
rect 302790 214432 302846 214441
rect 302790 214367 302846 214376
rect 302608 212492 302660 212498
rect 302608 212434 302660 212440
rect 302620 212129 302648 212434
rect 302606 212120 302662 212129
rect 302606 212055 302662 212064
rect 302792 211132 302844 211138
rect 302792 211074 302844 211080
rect 302804 209953 302832 211074
rect 302790 209944 302846 209953
rect 302790 209879 302846 209888
rect 302792 208344 302844 208350
rect 302792 208286 302844 208292
rect 302804 207777 302832 208286
rect 302790 207768 302846 207777
rect 302790 207703 302846 207712
rect 302792 205624 302844 205630
rect 302790 205592 302792 205601
rect 302844 205592 302846 205601
rect 302790 205527 302846 205536
rect 302238 203416 302294 203425
rect 302238 203351 302294 203360
rect 302896 201249 302924 459410
rect 302988 438977 303016 459478
rect 302974 438968 303030 438977
rect 302974 438903 303030 438912
rect 304276 320142 304304 539582
rect 304368 324494 304396 542370
rect 304460 329458 304488 545090
rect 305734 543824 305790 543833
rect 305734 543759 305790 543768
rect 305642 539608 305698 539617
rect 305642 539543 305698 539552
rect 304448 329452 304500 329458
rect 304448 329394 304500 329400
rect 304356 324488 304408 324494
rect 304356 324430 304408 324436
rect 305656 322726 305684 539543
rect 305748 326942 305776 543759
rect 305840 331158 305868 546479
rect 307666 545184 307722 545193
rect 307666 545119 307668 545128
rect 307720 545119 307722 545128
rect 307668 545090 307720 545096
rect 307206 542464 307262 542473
rect 307206 542399 307208 542408
rect 307260 542399 307262 542408
rect 307208 542370 307260 542376
rect 307298 540424 307354 540433
rect 307298 540359 307354 540368
rect 307312 539617 307340 540359
rect 307666 539880 307722 539889
rect 307666 539815 307722 539824
rect 307680 539646 307708 539815
rect 307668 539640 307720 539646
rect 307298 539608 307354 539617
rect 307668 539582 307720 539588
rect 307298 539543 307354 539552
rect 307022 537568 307078 537577
rect 307022 537503 307078 537512
rect 305918 480312 305974 480321
rect 305918 480247 305974 480256
rect 305828 331152 305880 331158
rect 305828 331094 305880 331100
rect 305736 326936 305788 326942
rect 305736 326878 305788 326884
rect 305644 322720 305696 322726
rect 305644 322662 305696 322668
rect 304264 320136 304316 320142
rect 304264 320078 304316 320084
rect 305932 295934 305960 480247
rect 307036 318374 307064 537503
rect 388444 536852 388496 536858
rect 388444 536794 388496 536800
rect 307114 478136 307170 478145
rect 307114 478071 307170 478080
rect 307128 477562 307156 478071
rect 307116 477556 307168 477562
rect 307116 477498 307168 477504
rect 351826 459640 351882 459649
rect 351826 459575 351882 459584
rect 327906 459504 327962 459513
rect 327906 459439 327962 459448
rect 313738 458144 313794 458153
rect 313738 458079 313794 458088
rect 321558 458144 321614 458153
rect 321558 458079 321614 458088
rect 322938 458144 322994 458153
rect 322938 458079 322994 458088
rect 325698 458144 325754 458153
rect 325698 458079 325754 458088
rect 327078 458144 327134 458153
rect 327078 458079 327134 458088
rect 313752 457502 313780 458079
rect 317418 457872 317474 457881
rect 317418 457807 317474 457816
rect 313740 457496 313792 457502
rect 313740 457438 313792 457444
rect 309784 457428 309836 457434
rect 309784 457370 309836 457376
rect 308404 457020 308456 457026
rect 308404 456962 308456 456968
rect 307024 318368 307076 318374
rect 307024 318310 307076 318316
rect 305920 295928 305972 295934
rect 305920 295870 305972 295876
rect 308416 285326 308444 456962
rect 308404 285320 308456 285326
rect 308404 285262 308456 285268
rect 309796 223582 309824 457370
rect 312544 457292 312596 457298
rect 312544 457234 312596 457240
rect 309784 223576 309836 223582
rect 309784 223518 309836 223524
rect 312556 219434 312584 457234
rect 315304 457156 315356 457162
rect 315304 457098 315356 457104
rect 312544 219428 312596 219434
rect 312544 219370 312596 219376
rect 315316 216646 315344 457098
rect 317432 457026 317460 457807
rect 320270 457056 320326 457065
rect 317420 457020 317472 457026
rect 320270 456991 320326 457000
rect 317420 456962 317472 456968
rect 316038 456920 316094 456929
rect 316038 456855 316094 456864
rect 318798 456920 318854 456929
rect 318798 456855 318854 456864
rect 320178 456920 320234 456929
rect 320178 456855 320234 456864
rect 316052 315994 316080 456855
rect 316684 456816 316736 456822
rect 316684 456758 316736 456764
rect 316040 315988 316092 315994
rect 316040 315930 316092 315936
rect 315304 216640 315356 216646
rect 315304 216582 315356 216588
rect 316696 211138 316724 456758
rect 318812 287026 318840 456855
rect 320192 289814 320220 456855
rect 320284 292534 320312 456991
rect 320272 292528 320324 292534
rect 320272 292470 320324 292476
rect 320180 289808 320232 289814
rect 320180 289750 320232 289756
rect 318800 287020 318852 287026
rect 318800 286962 318852 286968
rect 316684 211132 316736 211138
rect 316684 211074 316736 211080
rect 321572 205630 321600 458079
rect 322202 458008 322258 458017
rect 322202 457943 322258 457952
rect 322216 457366 322244 457943
rect 322204 457360 322256 457366
rect 322204 457302 322256 457308
rect 322216 351898 322244 457302
rect 322204 351892 322256 351898
rect 322204 351834 322256 351840
rect 322952 208350 322980 458079
rect 323582 458008 323638 458017
rect 323582 457943 323638 457952
rect 323596 457094 323624 457943
rect 324962 457872 325018 457881
rect 324962 457807 325018 457816
rect 324318 457192 324374 457201
rect 324318 457127 324374 457136
rect 323584 457088 323636 457094
rect 323584 457030 323636 457036
rect 323492 434716 323544 434722
rect 323492 434658 323544 434664
rect 323504 434518 323532 434658
rect 323492 434512 323544 434518
rect 323492 434454 323544 434460
rect 323596 353258 323624 457030
rect 324332 456822 324360 457127
rect 324976 456958 325004 457807
rect 324964 456952 325016 456958
rect 324964 456894 325016 456900
rect 324320 456816 324372 456822
rect 324320 456758 324372 456764
rect 324976 356046 325004 456894
rect 324964 356040 325016 356046
rect 324964 355982 325016 355988
rect 323584 353252 323636 353258
rect 323584 353194 323636 353200
rect 325712 212498 325740 458079
rect 326342 457872 326398 457881
rect 326342 457807 326398 457816
rect 326356 456890 326384 457807
rect 326344 456884 326396 456890
rect 326344 456826 326396 456832
rect 326356 358766 326384 456826
rect 326344 358760 326396 358766
rect 326344 358702 326396 358708
rect 327092 215286 327120 458079
rect 327920 457230 327948 459439
rect 335360 458176 335412 458182
rect 329102 458144 329158 458153
rect 329102 458079 329104 458088
rect 329156 458079 329158 458088
rect 329930 458144 329986 458153
rect 329930 458079 329986 458088
rect 331862 458144 331918 458153
rect 331862 458079 331918 458088
rect 333150 458144 333206 458153
rect 333150 458079 333206 458088
rect 334070 458144 334126 458153
rect 334070 458079 334126 458088
rect 335358 458144 335360 458153
rect 344744 458176 344796 458182
rect 335412 458144 335414 458153
rect 336554 458144 336610 458153
rect 335414 458102 335492 458130
rect 335358 458079 335414 458088
rect 329104 458050 329156 458056
rect 327908 457224 327960 457230
rect 327908 457166 327960 457172
rect 328458 457192 328514 457201
rect 327920 454073 327948 457166
rect 328458 457127 328460 457136
rect 328512 457127 328514 457136
rect 328460 457098 328512 457104
rect 327722 454064 327778 454073
rect 327722 453999 327778 454008
rect 327906 454064 327962 454073
rect 327906 453999 327962 454008
rect 327736 444446 327764 453999
rect 327632 444440 327684 444446
rect 327552 444388 327632 444394
rect 327552 444382 327684 444388
rect 327724 444440 327776 444446
rect 327724 444382 327776 444388
rect 327552 444366 327672 444382
rect 327552 437594 327580 444366
rect 327552 437566 327672 437594
rect 327644 437458 327672 437566
rect 327552 437430 327672 437458
rect 327552 434722 327580 437430
rect 327540 434716 327592 434722
rect 327540 434658 327592 434664
rect 327632 434716 327684 434722
rect 327632 434658 327684 434664
rect 327724 434716 327776 434722
rect 327724 434658 327776 434664
rect 327644 423706 327672 434658
rect 327736 434518 327764 434658
rect 327724 434512 327776 434518
rect 327724 434454 327776 434460
rect 327540 423700 327592 423706
rect 327540 423642 327592 423648
rect 327632 423700 327684 423706
rect 327632 423642 327684 423648
rect 327552 413982 327580 423642
rect 327540 413976 327592 413982
rect 327540 413918 327592 413924
rect 327724 413976 327776 413982
rect 327724 413918 327776 413924
rect 327736 404394 327764 413918
rect 327540 404388 327592 404394
rect 327540 404330 327592 404336
rect 327724 404388 327776 404394
rect 327724 404330 327776 404336
rect 327552 394670 327580 404330
rect 327540 394664 327592 394670
rect 327540 394606 327592 394612
rect 327632 394664 327684 394670
rect 327632 394606 327684 394612
rect 327644 385082 327672 394606
rect 327632 385076 327684 385082
rect 327632 385018 327684 385024
rect 327816 385076 327868 385082
rect 327816 385018 327868 385024
rect 327828 376786 327856 385018
rect 327632 376780 327684 376786
rect 327632 376722 327684 376728
rect 327816 376780 327868 376786
rect 327816 376722 327868 376728
rect 327644 369866 327672 376722
rect 327644 369838 327856 369866
rect 327828 367033 327856 369838
rect 327814 367024 327870 367033
rect 327814 366959 327870 366968
rect 328090 367024 328146 367033
rect 328090 366959 328146 366968
rect 328104 360194 328132 366959
rect 329116 362914 329144 458050
rect 329286 458008 329342 458017
rect 329286 457943 329342 457952
rect 329300 457162 329328 457943
rect 329838 457328 329894 457337
rect 329838 457263 329840 457272
rect 329892 457263 329894 457272
rect 329840 457234 329892 457240
rect 329288 457156 329340 457162
rect 329288 457098 329340 457104
rect 329300 364342 329328 457098
rect 329288 364336 329340 364342
rect 329288 364278 329340 364284
rect 329104 362908 329156 362914
rect 329104 362850 329156 362856
rect 328092 360188 328144 360194
rect 328092 360130 328144 360136
rect 329944 222154 329972 458079
rect 331876 457910 331904 458079
rect 331312 457904 331364 457910
rect 330482 457872 330538 457881
rect 331312 457846 331364 457852
rect 331864 457904 331916 457910
rect 331864 457846 331916 457852
rect 330482 457807 330538 457816
rect 330496 456822 330524 457807
rect 331218 457736 331274 457745
rect 331218 457671 331274 457680
rect 331232 457434 331260 457671
rect 331220 457428 331272 457434
rect 331220 457370 331272 457376
rect 331324 457366 331352 457846
rect 333164 457774 333192 458079
rect 332600 457768 332652 457774
rect 332600 457710 332652 457716
rect 333152 457768 333204 457774
rect 333152 457710 333204 457716
rect 331312 457360 331364 457366
rect 331312 457302 331364 457308
rect 332612 457094 332640 457710
rect 334084 457570 334112 458079
rect 334072 457564 334124 457570
rect 334072 457506 334124 457512
rect 332600 457088 332652 457094
rect 332600 457030 332652 457036
rect 334084 456958 334112 457506
rect 335358 457192 335414 457201
rect 335358 457127 335414 457136
rect 334072 456952 334124 456958
rect 332598 456920 332654 456929
rect 332598 456855 332654 456864
rect 333978 456920 334034 456929
rect 334072 456894 334124 456900
rect 333978 456855 334034 456864
rect 330484 456816 330536 456822
rect 330484 456758 330536 456764
rect 330496 367062 330524 456758
rect 330484 367056 330536 367062
rect 330484 366998 330536 367004
rect 332612 226302 332640 456855
rect 333992 227730 334020 456855
rect 335372 230450 335400 457127
rect 335464 456890 335492 458102
rect 336554 458079 336610 458088
rect 338026 458144 338082 458153
rect 338026 458079 338028 458088
rect 336568 457978 336596 458079
rect 338080 458079 338082 458088
rect 339038 458144 339094 458153
rect 339038 458079 339094 458088
rect 339866 458144 339922 458153
rect 339866 458079 339922 458088
rect 341246 458144 341302 458153
rect 341246 458079 341302 458088
rect 342258 458144 342314 458153
rect 342258 458079 342314 458088
rect 343638 458144 343694 458153
rect 344742 458144 344744 458153
rect 344796 458144 344798 458153
rect 343638 458079 343694 458088
rect 344376 458108 344428 458114
rect 338028 458050 338080 458056
rect 336556 457972 336608 457978
rect 336556 457914 336608 457920
rect 336568 457230 336596 457914
rect 338040 457706 338068 458050
rect 339052 457842 339080 458079
rect 339040 457836 339092 457842
rect 339040 457778 339092 457784
rect 338028 457700 338080 457706
rect 338028 457642 338080 457648
rect 336556 457224 336608 457230
rect 336556 457166 336608 457172
rect 339052 457162 339080 457778
rect 339880 457638 339908 458079
rect 341260 457910 341288 458079
rect 341248 457904 341300 457910
rect 341248 457846 341300 457852
rect 340880 457836 340932 457842
rect 340880 457778 340932 457784
rect 339868 457632 339920 457638
rect 339868 457574 339920 457580
rect 339040 457156 339092 457162
rect 339040 457098 339092 457104
rect 336830 457056 336886 457065
rect 336830 456991 336886 457000
rect 336738 456920 336794 456929
rect 335452 456884 335504 456890
rect 336738 456855 336794 456864
rect 335452 456826 335504 456832
rect 336752 233238 336780 456855
rect 336844 234598 336872 456991
rect 338118 456920 338174 456929
rect 338118 456855 338174 456864
rect 339498 456920 339554 456929
rect 339498 456855 339554 456864
rect 338132 237386 338160 456855
rect 339512 238746 339540 456855
rect 339880 456822 339908 457574
rect 340892 457434 340920 457778
rect 340880 457428 340932 457434
rect 340880 457370 340932 457376
rect 340878 457192 340934 457201
rect 340878 457127 340934 457136
rect 339868 456816 339920 456822
rect 339868 456758 339920 456764
rect 340892 241466 340920 457127
rect 342272 244254 342300 458079
rect 343548 458040 343600 458046
rect 342534 458008 342590 458017
rect 343548 457982 343600 457988
rect 342534 457943 342590 457952
rect 342548 457774 342576 457943
rect 343560 457774 343588 457982
rect 342536 457768 342588 457774
rect 342536 457710 342588 457716
rect 343548 457768 343600 457774
rect 343548 457710 343600 457716
rect 342904 457360 342956 457366
rect 342904 457302 342956 457308
rect 342916 371210 342944 457302
rect 342904 371204 342956 371210
rect 342904 371146 342956 371152
rect 343652 245614 343680 458079
rect 344742 458079 344798 458088
rect 345018 458144 345074 458153
rect 345018 458079 345074 458088
rect 346398 458144 346454 458153
rect 346398 458079 346454 458088
rect 347778 458144 347834 458153
rect 347778 458079 347834 458088
rect 349158 458144 349214 458153
rect 349158 458079 349214 458088
rect 344376 458050 344428 458056
rect 344388 458017 344416 458050
rect 344374 458008 344430 458017
rect 344374 457943 344430 457952
rect 343730 457736 343786 457745
rect 343730 457671 343786 457680
rect 343744 248402 343772 457671
rect 344388 457570 344416 457943
rect 344376 457564 344428 457570
rect 344376 457506 344428 457512
rect 345032 249762 345060 458079
rect 345938 458008 345994 458017
rect 345938 457943 345940 457952
rect 345992 457943 345994 457952
rect 345940 457914 345992 457920
rect 346412 252550 346440 458079
rect 346858 458008 346914 458017
rect 346858 457943 346914 457952
rect 346872 457706 346900 457943
rect 346860 457700 346912 457706
rect 346860 457642 346912 457648
rect 347044 457020 347096 457026
rect 347044 456962 347096 456968
rect 347056 415410 347084 456962
rect 347044 415404 347096 415410
rect 347044 415346 347096 415352
rect 347792 255270 347820 458079
rect 348238 458008 348294 458017
rect 348238 457943 348294 457952
rect 348252 457434 348280 457943
rect 348240 457428 348292 457434
rect 348240 457370 348292 457376
rect 349172 256698 349200 458079
rect 351840 458046 351868 459575
rect 358818 459504 358874 459513
rect 358818 459439 358874 459448
rect 353300 458176 353352 458182
rect 351918 458144 351974 458153
rect 353298 458144 353300 458153
rect 354036 458176 354088 458182
rect 353352 458144 353354 458153
rect 351918 458079 351920 458088
rect 351972 458079 351974 458088
rect 352748 458108 352800 458114
rect 351920 458050 351972 458056
rect 354036 458118 354088 458124
rect 353298 458079 353354 458088
rect 352748 458050 352800 458056
rect 351828 458040 351880 458046
rect 349250 458008 349306 458017
rect 349250 457943 349306 457952
rect 350538 458008 350594 458017
rect 351828 457982 351880 457988
rect 350538 457943 350594 457952
rect 349264 457774 349292 457943
rect 350552 457910 350580 457943
rect 350540 457904 350592 457910
rect 350540 457846 350592 457852
rect 350632 457904 350684 457910
rect 350632 457846 350684 457852
rect 349252 457768 349304 457774
rect 349252 457710 349304 457716
rect 349712 457768 349764 457774
rect 349712 457710 349764 457716
rect 349264 457638 349292 457710
rect 349252 457632 349304 457638
rect 349252 457574 349304 457580
rect 349724 457434 349752 457710
rect 350644 457638 350672 457846
rect 350632 457632 350684 457638
rect 350632 457574 350684 457580
rect 349712 457428 349764 457434
rect 349712 457370 349764 457376
rect 349804 457292 349856 457298
rect 349804 457234 349856 457240
rect 349816 418130 349844 457234
rect 351184 457224 351236 457230
rect 351184 457166 351236 457172
rect 350538 456920 350594 456929
rect 350538 456855 350594 456864
rect 349804 418124 349856 418130
rect 349804 418066 349856 418072
rect 350552 259418 350580 456855
rect 351196 419490 351224 457166
rect 352564 457156 352616 457162
rect 352564 457098 352616 457104
rect 352010 457056 352066 457065
rect 352010 456991 352066 457000
rect 351918 456920 351974 456929
rect 351918 456855 351974 456864
rect 351184 419484 351236 419490
rect 351184 419426 351236 419432
rect 351932 260846 351960 456855
rect 352024 263566 352052 456991
rect 352576 422278 352604 457098
rect 352656 457088 352708 457094
rect 352656 457030 352708 457036
rect 352668 423638 352696 457030
rect 352760 426426 352788 458050
rect 353944 458040 353996 458046
rect 353944 457982 353996 457988
rect 353668 457972 353720 457978
rect 353668 457914 353720 457920
rect 353680 457570 353708 457914
rect 353668 457564 353720 457570
rect 353668 457506 353720 457512
rect 353298 457192 353354 457201
rect 353298 457127 353354 457136
rect 352748 426420 352800 426426
rect 352748 426362 352800 426368
rect 352656 423632 352708 423638
rect 352656 423574 352708 423580
rect 352564 422272 352616 422278
rect 352564 422214 352616 422220
rect 353312 266354 353340 457127
rect 353956 429146 353984 457982
rect 354048 430574 354076 458118
rect 356058 458008 356114 458017
rect 356058 457943 356114 457952
rect 356072 457910 356100 457943
rect 356060 457904 356112 457910
rect 355046 457872 355102 457881
rect 356060 457846 356112 457852
rect 355046 457807 355102 457816
rect 355060 457570 355088 457807
rect 357438 457736 357494 457745
rect 357438 457671 357440 457680
rect 357492 457671 357494 457680
rect 357440 457642 357492 457648
rect 358832 457638 358860 459439
rect 359464 457700 359516 457706
rect 359464 457642 359516 457648
rect 358820 457632 358872 457638
rect 358820 457574 358872 457580
rect 355048 457564 355100 457570
rect 355048 457506 355100 457512
rect 358084 457564 358136 457570
rect 358084 457506 358136 457512
rect 355324 457428 355376 457434
rect 355324 457370 355376 457376
rect 354678 456920 354734 456929
rect 354678 456855 354734 456864
rect 354036 430568 354088 430574
rect 354036 430510 354088 430516
rect 353944 429140 353996 429146
rect 353944 429082 353996 429088
rect 354692 267714 354720 456855
rect 355336 373998 355364 457370
rect 356058 456920 356114 456929
rect 357438 456920 357494 456929
rect 356058 456855 356114 456864
rect 356704 456884 356756 456890
rect 355324 373992 355376 373998
rect 355324 373934 355376 373940
rect 356072 270502 356100 456855
rect 357438 456855 357494 456864
rect 356704 456826 356756 456832
rect 356716 375358 356744 456826
rect 356704 375352 356756 375358
rect 356704 375294 356756 375300
rect 357452 271862 357480 456855
rect 358096 378146 358124 457506
rect 358818 456920 358874 456929
rect 358818 456855 358874 456864
rect 358084 378140 358136 378146
rect 358084 378082 358136 378088
rect 358832 274650 358860 456855
rect 359476 380866 359504 457642
rect 359464 380860 359516 380866
rect 359464 380802 359516 380808
rect 388456 300830 388484 536794
rect 389192 489569 389220 547862
rect 399484 546508 399536 546514
rect 399484 546450 399536 546456
rect 398104 545148 398156 545154
rect 398104 545090 398156 545096
rect 395344 543788 395396 543794
rect 395344 543730 395396 543736
rect 393964 542428 394016 542434
rect 393964 542370 394016 542376
rect 392584 539708 392636 539714
rect 392584 539650 392636 539656
rect 391204 539640 391256 539646
rect 391204 539582 391256 539588
rect 389178 489560 389234 489569
rect 389178 489495 389234 489504
rect 389178 480992 389234 481001
rect 389178 480927 389234 480936
rect 389192 459474 389220 480927
rect 389180 459468 389232 459474
rect 389180 459410 389232 459416
rect 391216 303618 391244 539582
rect 392596 304978 392624 539650
rect 393976 307766 394004 542370
rect 395356 309126 395384 543730
rect 398116 311846 398144 545090
rect 399496 314634 399524 546450
rect 429580 543833 429608 550598
rect 516416 550316 516468 550322
rect 516416 550258 516468 550264
rect 516428 549953 516456 550258
rect 516414 549944 516470 549953
rect 516414 549879 516470 549888
rect 437478 546544 437534 546553
rect 437478 546479 437480 546488
rect 437532 546479 437534 546488
rect 437480 546450 437532 546456
rect 437478 545184 437534 545193
rect 437478 545119 437480 545128
rect 437532 545119 437534 545128
rect 437480 545090 437532 545096
rect 429566 543824 429622 543833
rect 429566 543759 429622 543768
rect 437478 543824 437534 543833
rect 437478 543759 437480 543768
rect 437532 543759 437534 543768
rect 437480 543730 437532 543736
rect 429382 543688 429438 543697
rect 429382 543623 429438 543632
rect 429396 540977 429424 543623
rect 437478 542464 437534 542473
rect 437478 542399 437480 542408
rect 437532 542399 437534 542408
rect 437480 542370 437532 542376
rect 429198 540968 429254 540977
rect 429198 540903 429254 540912
rect 429382 540968 429438 540977
rect 429382 540903 429438 540912
rect 429212 531350 429240 540903
rect 437570 540424 437626 540433
rect 437570 540359 437626 540368
rect 437478 539880 437534 539889
rect 437478 539815 437534 539824
rect 437492 539646 437520 539815
rect 437584 539714 437612 540359
rect 437572 539708 437624 539714
rect 437572 539650 437624 539656
rect 437480 539640 437532 539646
rect 437480 539582 437532 539588
rect 437478 537568 437534 537577
rect 437478 537503 437534 537512
rect 437492 536858 437520 537503
rect 437480 536852 437532 536858
rect 437480 536794 437532 536800
rect 429200 531344 429252 531350
rect 429200 531286 429252 531292
rect 429476 531344 429528 531350
rect 429476 531286 429528 531292
rect 429488 524482 429516 531286
rect 429476 524476 429528 524482
rect 429476 524418 429528 524424
rect 429568 524408 429620 524414
rect 429568 524350 429620 524356
rect 429580 521665 429608 524350
rect 429382 521656 429438 521665
rect 429382 521591 429438 521600
rect 429566 521656 429622 521665
rect 429566 521591 429622 521600
rect 429396 512038 429424 521591
rect 429384 512032 429436 512038
rect 429384 511974 429436 511980
rect 429660 512032 429712 512038
rect 429660 511974 429712 511980
rect 429672 502382 429700 511974
rect 429476 502376 429528 502382
rect 429476 502318 429528 502324
rect 429660 502376 429712 502382
rect 429660 502318 429712 502324
rect 429488 485858 429516 502318
rect 518912 489569 518940 550695
rect 559024 550662 559052 553318
rect 558920 550656 558972 550662
rect 558920 550598 558972 550604
rect 559012 550656 559064 550662
rect 559012 550598 559064 550604
rect 558932 543794 558960 550598
rect 580262 545592 580318 545601
rect 580262 545527 580318 545536
rect 558920 543788 558972 543794
rect 558920 543730 558972 543736
rect 559012 543652 559064 543658
rect 559012 543594 559064 543600
rect 559024 534070 559052 543594
rect 559012 534064 559064 534070
rect 559012 534006 559064 534012
rect 559196 534064 559248 534070
rect 559196 534006 559248 534012
rect 559208 524482 559236 534006
rect 559196 524476 559248 524482
rect 559196 524418 559248 524424
rect 559288 524408 559340 524414
rect 559288 524350 559340 524356
rect 559300 521665 559328 524350
rect 559102 521656 559158 521665
rect 559102 521591 559158 521600
rect 559286 521656 559342 521665
rect 559286 521591 559342 521600
rect 559116 512038 559144 521591
rect 559104 512032 559156 512038
rect 559104 511974 559156 511980
rect 559380 512032 559432 512038
rect 559380 511974 559432 511980
rect 559392 502382 559420 511974
rect 559196 502376 559248 502382
rect 559196 502318 559248 502324
rect 559380 502376 559432 502382
rect 559380 502318 559432 502324
rect 559208 492833 559236 502318
rect 559194 492824 559250 492833
rect 559194 492759 559250 492768
rect 559102 492688 559158 492697
rect 559102 492623 559104 492632
rect 559156 492623 559158 492632
rect 559196 492652 559248 492658
rect 559104 492594 559156 492600
rect 559196 492594 559248 492600
rect 518898 489560 518954 489569
rect 518898 489495 518954 489504
rect 429476 485852 429528 485858
rect 429476 485794 429528 485800
rect 559208 485790 559236 492594
rect 429568 485784 429620 485790
rect 429568 485726 429620 485732
rect 559104 485784 559156 485790
rect 559104 485726 559156 485732
rect 559196 485784 559248 485790
rect 559196 485726 559248 485732
rect 429580 483002 429608 485726
rect 559116 483018 559144 485726
rect 429568 482996 429620 483002
rect 429568 482938 429620 482944
rect 429660 482996 429712 483002
rect 559116 482990 559236 483018
rect 429660 482938 429712 482944
rect 402244 480276 402296 480282
rect 402244 480218 402296 480224
rect 399484 314628 399536 314634
rect 399484 314570 399536 314576
rect 398104 311840 398156 311846
rect 398104 311782 398156 311788
rect 395344 309120 395396 309126
rect 395344 309062 395396 309068
rect 393964 307760 394016 307766
rect 393964 307702 394016 307708
rect 392584 304972 392636 304978
rect 392584 304914 392636 304920
rect 391204 303612 391256 303618
rect 391204 303554 391256 303560
rect 388444 300824 388496 300830
rect 388444 300766 388496 300772
rect 402256 293962 402284 480218
rect 429672 476134 429700 482938
rect 437478 480312 437534 480321
rect 437478 480247 437480 480256
rect 437532 480247 437534 480256
rect 437480 480218 437532 480224
rect 438122 478000 438178 478009
rect 438122 477935 438178 477944
rect 429660 476128 429712 476134
rect 429660 476070 429712 476076
rect 429568 476060 429620 476066
rect 429568 476002 429620 476008
rect 429580 473362 429608 476002
rect 429580 473334 429700 473362
rect 429672 463729 429700 473334
rect 429474 463720 429530 463729
rect 429474 463655 429530 463664
rect 429658 463720 429714 463729
rect 429658 463655 429714 463664
rect 429488 447234 429516 463655
rect 438136 459542 438164 477935
rect 559208 476134 559236 482990
rect 559012 476128 559064 476134
rect 559196 476128 559248 476134
rect 559064 476076 559144 476082
rect 559012 476070 559144 476076
rect 559196 476070 559248 476076
rect 559024 476054 559144 476070
rect 559116 473346 559144 476054
rect 559104 473340 559156 473346
rect 559104 473282 559156 473288
rect 559196 473340 559248 473346
rect 559196 473282 559248 473288
rect 559208 466478 559236 473282
rect 559196 466472 559248 466478
rect 559196 466414 559248 466420
rect 559104 466404 559156 466410
rect 559104 466346 559156 466352
rect 559116 463706 559144 466346
rect 559116 463678 559236 463706
rect 438124 459536 438176 459542
rect 438124 459478 438176 459484
rect 483018 459504 483074 459513
rect 483074 459462 483152 459490
rect 483018 459439 483074 459448
rect 461766 458144 461822 458153
rect 461766 458079 461822 458088
rect 463054 458144 463110 458153
rect 463054 458079 463110 458088
rect 464986 458144 465042 458153
rect 464986 458079 465042 458088
rect 465170 458144 465226 458153
rect 465170 458079 465226 458088
rect 468758 458144 468814 458153
rect 468758 458079 468814 458088
rect 469954 458144 470010 458153
rect 469954 458079 470010 458088
rect 471794 458144 471850 458153
rect 471794 458079 471850 458088
rect 472254 458144 472310 458153
rect 472254 458079 472310 458088
rect 473450 458144 473506 458153
rect 473450 458079 473506 458088
rect 474830 458144 474886 458153
rect 474830 458079 474886 458088
rect 475474 458144 475530 458153
rect 475474 458079 475530 458088
rect 476946 458144 477002 458153
rect 476946 458079 477002 458088
rect 478326 458144 478382 458153
rect 478326 458079 478382 458088
rect 479430 458144 479486 458153
rect 479430 458079 479486 458088
rect 483018 458144 483074 458153
rect 483018 458079 483020 458088
rect 442998 458008 443054 458017
rect 442998 457943 443054 457952
rect 460202 458008 460258 458017
rect 460202 457943 460258 457952
rect 443012 457502 443040 457943
rect 460216 457910 460244 457943
rect 460204 457904 460256 457910
rect 458178 457872 458234 457881
rect 460204 457846 460256 457852
rect 458178 457807 458234 457816
rect 453488 457768 453540 457774
rect 453488 457710 453540 457716
rect 453304 457632 453356 457638
rect 453304 457574 453356 457580
rect 443000 457496 443052 457502
rect 443000 457438 443052 457444
rect 443644 457496 443696 457502
rect 443644 457438 443696 457444
rect 452658 457464 452714 457473
rect 429476 447228 429528 447234
rect 429476 447170 429528 447176
rect 429476 447092 429528 447098
rect 429476 447034 429528 447040
rect 429488 444446 429516 447034
rect 429384 444440 429436 444446
rect 429384 444382 429436 444388
rect 429476 444440 429528 444446
rect 429476 444382 429528 444388
rect 429396 439686 429424 444382
rect 429384 439680 429436 439686
rect 429384 439622 429436 439628
rect 443656 382226 443684 457438
rect 452658 457399 452714 457408
rect 452672 457366 452700 457399
rect 452660 457360 452712 457366
rect 452660 457302 452712 457308
rect 450542 457192 450598 457201
rect 450542 457127 450598 457136
rect 446402 457056 446458 457065
rect 446402 456991 446458 457000
rect 445758 456920 445814 456929
rect 445758 456855 445814 456864
rect 443644 382220 443696 382226
rect 443644 382162 443696 382168
rect 445772 298110 445800 456855
rect 445760 298104 445812 298110
rect 445760 298046 445812 298052
rect 402244 293956 402296 293962
rect 402244 293898 402296 293904
rect 446416 277370 446444 456991
rect 447782 456920 447838 456929
rect 447782 456855 447838 456864
rect 449162 456920 449218 456929
rect 449162 456855 449218 456864
rect 447796 278730 447824 456855
rect 449176 281518 449204 456855
rect 450556 282878 450584 457127
rect 453316 456929 453344 457574
rect 453500 456929 453528 457710
rect 458192 457706 458220 457807
rect 458180 457700 458232 457706
rect 458180 457642 458232 457648
rect 456798 457600 456854 457609
rect 456798 457535 456800 457544
rect 456852 457535 456854 457544
rect 459558 457600 459614 457609
rect 459558 457535 459614 457544
rect 456800 457506 456852 457512
rect 459572 457502 459600 457535
rect 459560 457496 459612 457502
rect 454038 457464 454094 457473
rect 459560 457438 459612 457444
rect 454038 457399 454040 457408
rect 454092 457399 454094 457408
rect 454684 457428 454736 457434
rect 454040 457370 454092 457376
rect 454684 457370 454736 457376
rect 454696 457201 454724 457370
rect 454682 457192 454738 457201
rect 454682 457127 454738 457136
rect 458822 457192 458878 457201
rect 458822 457127 458878 457136
rect 459374 457192 459430 457201
rect 459374 457127 459430 457136
rect 452750 456920 452806 456929
rect 452750 456855 452806 456864
rect 453302 456920 453358 456929
rect 453302 456855 453358 456864
rect 453486 456920 453542 456929
rect 453486 456855 453542 456864
rect 452764 369850 452792 456855
rect 452752 369844 452804 369850
rect 452752 369786 452804 369792
rect 453316 333946 453344 456855
rect 453500 336734 453528 456855
rect 454696 338094 454724 457127
rect 456062 457056 456118 457065
rect 456062 456991 456118 457000
rect 456706 457056 456762 457065
rect 456706 456991 456762 457000
rect 455418 456920 455474 456929
rect 455418 456855 455420 456864
rect 455472 456855 455474 456864
rect 455420 456826 455472 456832
rect 456076 340882 456104 456991
rect 456720 456890 456748 456991
rect 457442 456920 457498 456929
rect 456708 456884 456760 456890
rect 457442 456855 457498 456864
rect 458086 456920 458142 456929
rect 458086 456855 458142 456864
rect 456708 456826 456760 456832
rect 457456 342242 457484 456855
rect 458100 456822 458128 456855
rect 458088 456816 458140 456822
rect 458088 456758 458140 456764
rect 458836 345030 458864 457127
rect 459388 456958 459416 457127
rect 459376 456952 459428 456958
rect 459376 456894 459428 456900
rect 460216 347750 460244 457846
rect 460386 457736 460442 457745
rect 460386 457671 460388 457680
rect 460440 457671 460442 457680
rect 460388 457642 460440 457648
rect 460400 349110 460428 457642
rect 461780 457638 461808 458079
rect 463068 457774 463096 458079
rect 465000 457842 465028 458079
rect 464988 457836 465040 457842
rect 464988 457778 465040 457784
rect 463056 457768 463108 457774
rect 463056 457710 463108 457716
rect 461768 457632 461820 457638
rect 461768 457574 461820 457580
rect 465000 457434 465028 457778
rect 465184 457570 465212 458079
rect 468022 458008 468078 458017
rect 468022 457943 468078 457952
rect 466642 457872 466698 457881
rect 466642 457807 466698 457816
rect 465172 457564 465224 457570
rect 465172 457506 465224 457512
rect 464988 457428 465040 457434
rect 464988 457370 465040 457376
rect 464344 457360 464396 457366
rect 464344 457302 464396 457308
rect 461030 457192 461086 457201
rect 461030 457127 461086 457136
rect 460938 456920 460994 456929
rect 460938 456855 460994 456864
rect 460952 385014 460980 456855
rect 461044 386374 461072 457127
rect 462318 456920 462374 456929
rect 462318 456855 462374 456864
rect 463698 456920 463754 456929
rect 463698 456855 463754 456864
rect 462332 389162 462360 456855
rect 463712 390522 463740 456855
rect 464356 433294 464384 457302
rect 465078 456920 465134 456929
rect 465184 456890 465212 457506
rect 465724 457496 465776 457502
rect 465724 457438 465776 457444
rect 465078 456855 465134 456864
rect 465172 456884 465224 456890
rect 464344 433288 464396 433294
rect 464344 433230 464396 433236
rect 465092 393310 465120 456855
rect 465172 456826 465224 456832
rect 465736 434722 465764 457438
rect 466458 456920 466514 456929
rect 466656 456890 466684 457807
rect 467104 457428 467156 457434
rect 467104 457370 467156 457376
rect 466458 456855 466514 456864
rect 466644 456884 466696 456890
rect 465724 434716 465776 434722
rect 465724 434658 465776 434664
rect 466472 396030 466500 456855
rect 466644 456826 466696 456832
rect 467116 437442 467144 457370
rect 467930 457192 467986 457201
rect 467930 457127 467986 457136
rect 467838 456920 467894 456929
rect 467838 456855 467894 456864
rect 467104 437436 467156 437442
rect 467104 437378 467156 437384
rect 467852 397458 467880 456855
rect 467944 400178 467972 457127
rect 468036 456958 468064 457943
rect 468772 457910 468800 458079
rect 468760 457904 468812 457910
rect 468760 457846 468812 457852
rect 469968 457706 469996 458079
rect 471808 457978 471836 458079
rect 471796 457972 471848 457978
rect 471796 457914 471848 457920
rect 471164 457842 471560 457858
rect 471164 457836 471572 457842
rect 471164 457830 471520 457836
rect 469956 457700 470008 457706
rect 469956 457642 470008 457648
rect 468024 456952 468076 456958
rect 468024 456894 468076 456900
rect 469218 456920 469274 456929
rect 469218 456855 469274 456864
rect 470598 456920 470654 456929
rect 471164 456890 471192 457830
rect 471520 457778 471572 457784
rect 471336 457768 471388 457774
rect 471336 457710 471388 457716
rect 471348 457570 471376 457710
rect 471808 457638 471836 457914
rect 472268 457638 472296 458079
rect 473464 457774 473492 458079
rect 473452 457768 473504 457774
rect 473452 457710 473504 457716
rect 471796 457632 471848 457638
rect 471796 457574 471848 457580
rect 472256 457632 472308 457638
rect 472256 457574 472308 457580
rect 471244 457564 471296 457570
rect 471244 457506 471296 457512
rect 471336 457564 471388 457570
rect 471336 457506 471388 457512
rect 471256 456890 471284 457506
rect 471978 457192 472034 457201
rect 471978 457127 472034 457136
rect 470598 456855 470654 456864
rect 471152 456884 471204 456890
rect 469232 401606 469260 456855
rect 470612 404326 470640 456855
rect 471152 456826 471204 456832
rect 471244 456884 471296 456890
rect 471244 456826 471296 456832
rect 471992 407114 472020 457127
rect 473358 456920 473414 456929
rect 473358 456855 473414 456864
rect 474738 456920 474794 456929
rect 474844 456890 474872 458079
rect 475488 457842 475516 458079
rect 475476 457836 475528 457842
rect 475476 457778 475528 457784
rect 476960 457570 476988 458079
rect 478340 457910 478368 458079
rect 478328 457904 478380 457910
rect 478328 457846 478380 457852
rect 478878 457872 478934 457881
rect 478878 457807 478934 457816
rect 476304 457564 476356 457570
rect 476304 457506 476356 457512
rect 476948 457564 477000 457570
rect 476948 457506 477000 457512
rect 476118 457328 476174 457337
rect 476118 457263 476174 457272
rect 476132 457026 476160 457263
rect 476210 457192 476266 457201
rect 476210 457127 476266 457136
rect 476120 457020 476172 457026
rect 476120 456962 476172 456968
rect 474738 456855 474794 456864
rect 474832 456884 474884 456890
rect 473372 408474 473400 456855
rect 474752 411262 474780 456855
rect 474832 456826 474884 456832
rect 476224 412622 476252 457127
rect 476316 456958 476344 457506
rect 477498 457328 477554 457337
rect 477498 457263 477500 457272
rect 477552 457263 477554 457272
rect 477500 457234 477552 457240
rect 478892 457230 478920 457807
rect 479444 457706 479472 458079
rect 483072 458079 483074 458088
rect 483020 458050 483072 458056
rect 480442 458008 480498 458017
rect 480442 457943 480444 457952
rect 480496 457943 480498 457952
rect 480444 457914 480496 457920
rect 480534 457872 480590 457881
rect 480534 457807 480590 457816
rect 480260 457768 480312 457774
rect 480260 457710 480312 457716
rect 479432 457700 479484 457706
rect 479432 457642 479484 457648
rect 480272 457298 480300 457710
rect 480260 457292 480312 457298
rect 480260 457234 480312 457240
rect 478880 457224 478932 457230
rect 478880 457166 478932 457172
rect 480548 457162 480576 457807
rect 481638 457736 481694 457745
rect 481638 457671 481694 457680
rect 481652 457638 481680 457671
rect 481640 457632 481692 457638
rect 481640 457574 481692 457580
rect 483018 457464 483074 457473
rect 483018 457399 483074 457408
rect 481638 457192 481694 457201
rect 480536 457156 480588 457162
rect 481638 457127 481694 457136
rect 480536 457098 480588 457104
rect 481652 457094 481680 457127
rect 481640 457088 481692 457094
rect 481640 457030 481692 457036
rect 476304 456952 476356 456958
rect 476304 456894 476356 456900
rect 483032 456890 483060 457399
rect 483124 457298 483152 459462
rect 484400 458176 484452 458182
rect 483202 458144 483258 458153
rect 483202 458079 483258 458088
rect 484398 458144 484400 458153
rect 484452 458144 484454 458153
rect 484398 458079 484454 458088
rect 483216 458046 483244 458079
rect 483204 458040 483256 458046
rect 483204 457982 483256 457988
rect 487158 458008 487214 458017
rect 487158 457943 487214 457952
rect 487172 457910 487200 457943
rect 487160 457904 487212 457910
rect 484398 457872 484454 457881
rect 487160 457846 487212 457852
rect 484398 457807 484400 457816
rect 484452 457807 484454 457816
rect 484400 457778 484452 457784
rect 485778 457736 485834 457745
rect 485778 457671 485834 457680
rect 488538 457736 488594 457745
rect 488538 457671 488540 457680
rect 485792 457570 485820 457671
rect 488592 457671 488594 457680
rect 488540 457642 488592 457648
rect 487158 457600 487214 457609
rect 485780 457564 485832 457570
rect 487158 457535 487214 457544
rect 485780 457506 485832 457512
rect 487172 457502 487200 457535
rect 487160 457496 487212 457502
rect 485778 457464 485834 457473
rect 487160 457438 487212 457444
rect 488538 457464 488594 457473
rect 485778 457399 485834 457408
rect 488538 457399 488540 457408
rect 485792 457366 485820 457399
rect 488592 457399 488594 457408
rect 488540 457370 488592 457376
rect 485780 457360 485832 457366
rect 485780 457302 485832 457308
rect 483112 457292 483164 457298
rect 483112 457234 483164 457240
rect 483020 456884 483072 456890
rect 483020 456826 483072 456832
rect 559208 456822 559236 463678
rect 559012 456816 559064 456822
rect 559196 456816 559248 456822
rect 559064 456764 559196 456770
rect 559012 456758 559248 456764
rect 559024 456742 559236 456758
rect 559208 447234 559236 456742
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 559196 447228 559248 447234
rect 559196 447170 559248 447176
rect 559196 447092 559248 447098
rect 559196 447034 559248 447040
rect 559208 444446 559236 447034
rect 559104 444440 559156 444446
rect 559104 444382 559156 444388
rect 559196 444440 559248 444446
rect 559196 444382 559248 444388
rect 559116 439657 559144 444382
rect 580078 439920 580134 439929
rect 580078 439855 580134 439864
rect 559102 439648 559158 439657
rect 559102 439583 559158 439592
rect 580092 439006 580120 439855
rect 580080 439000 580132 439006
rect 580080 438942 580132 438948
rect 580276 438190 580304 545527
rect 580354 533896 580410 533905
rect 580354 533831 580410 533840
rect 580368 439618 580396 533831
rect 580446 510368 580502 510377
rect 580446 510303 580502 510312
rect 580356 439612 580408 439618
rect 580356 439554 580408 439560
rect 580460 439521 580488 510303
rect 580538 498672 580594 498681
rect 580538 498607 580594 498616
rect 580446 439512 580502 439521
rect 580446 439447 580502 439456
rect 580552 438326 580580 498607
rect 580722 486840 580778 486849
rect 580722 486775 580778 486784
rect 580736 439550 580764 486775
rect 580814 463448 580870 463457
rect 580814 463383 580870 463392
rect 580724 439544 580776 439550
rect 580724 439486 580776 439492
rect 580632 438932 580684 438938
rect 580632 438874 580684 438880
rect 580540 438320 580592 438326
rect 580540 438262 580592 438268
rect 580264 438184 580316 438190
rect 580264 438126 580316 438132
rect 580356 438048 580408 438054
rect 580356 437990 580408 437996
rect 476212 412616 476264 412622
rect 476212 412558 476264 412564
rect 474740 411256 474792 411262
rect 474740 411198 474792 411204
rect 473360 408468 473412 408474
rect 473360 408410 473412 408416
rect 471980 407108 472032 407114
rect 471980 407050 472032 407056
rect 580368 404841 580396 437990
rect 580448 437980 580500 437986
rect 580448 437922 580500 437928
rect 580460 416537 580488 437922
rect 580446 416528 580502 416537
rect 580446 416463 580502 416472
rect 580354 404832 580410 404841
rect 580354 404767 580410 404776
rect 470600 404320 470652 404326
rect 470600 404262 470652 404268
rect 469220 401600 469272 401606
rect 469220 401542 469272 401548
rect 467932 400172 467984 400178
rect 467932 400114 467984 400120
rect 467840 397452 467892 397458
rect 467840 397394 467892 397400
rect 466460 396024 466512 396030
rect 466460 395966 466512 395972
rect 465080 393304 465132 393310
rect 465080 393246 465132 393252
rect 580644 393009 580672 438874
rect 580828 438258 580856 463383
rect 580816 438252 580868 438258
rect 580816 438194 580868 438200
rect 580630 393000 580686 393009
rect 580630 392935 580686 392944
rect 463700 390516 463752 390522
rect 463700 390458 463752 390464
rect 462320 389156 462372 389162
rect 462320 389098 462372 389104
rect 461032 386368 461084 386374
rect 461032 386310 461084 386316
rect 460940 385008 460992 385014
rect 460940 384950 460992 384956
rect 580262 369608 580318 369617
rect 580262 369543 580318 369552
rect 460388 349104 460440 349110
rect 460388 349046 460440 349052
rect 460204 347744 460256 347750
rect 460204 347686 460256 347692
rect 458824 345024 458876 345030
rect 458824 344966 458876 344972
rect 457444 342236 457496 342242
rect 457444 342178 457496 342184
rect 456064 340876 456116 340882
rect 456064 340818 456116 340824
rect 454684 338088 454736 338094
rect 454684 338030 454736 338036
rect 453488 336728 453540 336734
rect 453488 336670 453540 336676
rect 453304 333940 453356 333946
rect 453304 333882 453356 333888
rect 450544 282872 450596 282878
rect 450544 282814 450596 282820
rect 449164 281512 449216 281518
rect 449164 281454 449216 281460
rect 447784 278724 447836 278730
rect 447784 278666 447836 278672
rect 446404 277364 446456 277370
rect 446404 277306 446456 277312
rect 358820 274644 358872 274650
rect 358820 274586 358872 274592
rect 357440 271856 357492 271862
rect 357440 271798 357492 271804
rect 356060 270496 356112 270502
rect 356060 270438 356112 270444
rect 354680 267708 354732 267714
rect 354680 267650 354732 267656
rect 353300 266348 353352 266354
rect 353300 266290 353352 266296
rect 352012 263560 352064 263566
rect 352012 263502 352064 263508
rect 351920 260840 351972 260846
rect 351920 260782 351972 260788
rect 350540 259412 350592 259418
rect 350540 259354 350592 259360
rect 349160 256692 349212 256698
rect 349160 256634 349212 256640
rect 347780 255264 347832 255270
rect 347780 255206 347832 255212
rect 346400 252544 346452 252550
rect 346400 252486 346452 252492
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 345020 249756 345072 249762
rect 345020 249698 345072 249704
rect 343732 248396 343784 248402
rect 343732 248338 343784 248344
rect 343640 245608 343692 245614
rect 343640 245550 343692 245556
rect 342260 244248 342312 244254
rect 342260 244190 342312 244196
rect 340880 241460 340932 241466
rect 340880 241402 340932 241408
rect 339500 238740 339552 238746
rect 339500 238682 339552 238688
rect 338120 237380 338172 237386
rect 338120 237322 338172 237328
rect 336832 234592 336884 234598
rect 336832 234534 336884 234540
rect 336740 233232 336792 233238
rect 336740 233174 336792 233180
rect 335360 230444 335412 230450
rect 335360 230386 335412 230392
rect 580078 228848 580134 228857
rect 580078 228783 580134 228792
rect 333980 227724 334032 227730
rect 333980 227666 334032 227672
rect 332600 226296 332652 226302
rect 332600 226238 332652 226244
rect 329932 222148 329984 222154
rect 329932 222090 329984 222096
rect 579986 217016 580042 217025
rect 579986 216951 580042 216960
rect 327080 215280 327132 215286
rect 327080 215222 327132 215228
rect 325700 212492 325752 212498
rect 325700 212434 325752 212440
rect 322940 208344 322992 208350
rect 322940 208286 322992 208292
rect 321560 205624 321612 205630
rect 321560 205566 321612 205572
rect 579896 205420 579948 205426
rect 579896 205362 579948 205368
rect 302882 201240 302938 201249
rect 302882 201175 302938 201184
rect 60752 200654 61042 200682
rect 59820 200456 59872 200462
rect 59820 200398 59872 200404
rect 57888 199912 57940 199918
rect 57888 199854 57940 199860
rect 57888 197804 57940 197810
rect 57888 197746 57940 197752
rect 57796 17944 57848 17950
rect 57796 17886 57848 17892
rect 56416 4752 56468 4758
rect 56416 4694 56468 4700
rect 55220 4412 55272 4418
rect 55220 4354 55272 4360
rect 55048 3046 55168 3074
rect 55048 2990 55076 3046
rect 54024 2984 54076 2990
rect 54024 2926 54076 2932
rect 55036 2984 55088 2990
rect 55036 2926 55088 2932
rect 55128 2984 55180 2990
rect 55128 2926 55180 2932
rect 54036 480 54064 2926
rect 55140 2786 55168 2926
rect 55128 2780 55180 2786
rect 55128 2722 55180 2728
rect 55232 480 55260 4354
rect 56428 480 56456 4694
rect 57900 3346 57928 197746
rect 60004 6656 60056 6662
rect 60004 6598 60056 6604
rect 58808 4480 58860 4486
rect 58808 4422 58860 4428
rect 57624 3318 57928 3346
rect 57624 480 57652 3318
rect 58820 480 58848 4422
rect 60016 480 60044 6598
rect 60752 3126 60780 200654
rect 579908 200530 579936 205362
rect 580000 200802 580028 216951
rect 579988 200796 580040 200802
rect 579988 200738 580040 200744
rect 580092 200598 580120 228783
rect 580184 205426 580212 252175
rect 580172 205420 580224 205426
rect 580172 205362 580224 205368
rect 580170 205320 580226 205329
rect 580170 205255 580226 205264
rect 580184 200666 580212 205255
rect 580276 200705 580304 369543
rect 580354 357912 580410 357921
rect 580354 357847 580410 357856
rect 580262 200696 580318 200705
rect 580172 200660 580224 200666
rect 580262 200631 580318 200640
rect 580172 200602 580224 200608
rect 580080 200592 580132 200598
rect 580080 200534 580132 200540
rect 579896 200524 579948 200530
rect 579896 200466 579948 200472
rect 580368 200462 580396 357847
rect 580446 346080 580502 346089
rect 580446 346015 580502 346024
rect 580356 200456 580408 200462
rect 580356 200398 580408 200404
rect 62224 200110 63158 200138
rect 64984 200110 65274 200138
rect 66272 200110 67390 200138
rect 62224 3126 62252 200110
rect 64788 197872 64840 197878
rect 64788 197814 64840 197820
rect 63592 6588 63644 6594
rect 63592 6530 63644 6536
rect 62396 4548 62448 4554
rect 62396 4490 62448 4496
rect 60740 3120 60792 3126
rect 60740 3062 60792 3068
rect 62212 3120 62264 3126
rect 62212 3062 62264 3068
rect 61200 3052 61252 3058
rect 61200 2994 61252 3000
rect 61212 480 61240 2994
rect 62408 480 62436 4490
rect 63604 480 63632 6530
rect 64800 480 64828 197814
rect 64984 3194 65012 200110
rect 65524 5500 65576 5506
rect 65524 5442 65576 5448
rect 65536 4758 65564 5442
rect 65524 4752 65576 4758
rect 65524 4694 65576 4700
rect 65984 4616 66036 4622
rect 65984 4558 66036 4564
rect 65616 4140 65668 4146
rect 65616 4082 65668 4088
rect 65156 3392 65208 3398
rect 65156 3334 65208 3340
rect 65168 3262 65196 3334
rect 65628 3330 65656 4082
rect 65616 3324 65668 3330
rect 65616 3266 65668 3272
rect 65156 3256 65208 3262
rect 65156 3198 65208 3204
rect 64972 3188 65024 3194
rect 64972 3130 65024 3136
rect 65996 480 66024 4558
rect 66272 3194 66300 200110
rect 69492 198490 69520 200124
rect 70504 200110 71622 200138
rect 73172 200110 73738 200138
rect 74552 200110 75854 200138
rect 69480 198484 69532 198490
rect 69480 198426 69532 198432
rect 69480 4684 69532 4690
rect 69480 4626 69532 4632
rect 66260 3188 66312 3194
rect 66260 3130 66312 3136
rect 68284 3188 68336 3194
rect 68284 3130 68336 3136
rect 67180 3120 67232 3126
rect 67180 3062 67232 3068
rect 67192 480 67220 3062
rect 68296 480 68324 3130
rect 69492 480 69520 4626
rect 70504 3398 70532 200110
rect 71688 198688 71740 198694
rect 71688 198630 71740 198636
rect 71700 3398 71728 198630
rect 72976 197940 73028 197946
rect 72976 197882 73028 197888
rect 72988 3398 73016 197882
rect 73068 4752 73120 4758
rect 73068 4694 73120 4700
rect 70492 3392 70544 3398
rect 70492 3334 70544 3340
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 71872 3392 71924 3398
rect 71872 3334 71924 3340
rect 72976 3392 73028 3398
rect 72976 3334 73028 3340
rect 70688 480 70716 3334
rect 71884 480 71912 3334
rect 73080 480 73108 4694
rect 73172 3262 73200 200110
rect 74552 3330 74580 200110
rect 77956 198422 77984 200124
rect 79968 198620 80020 198626
rect 79968 198562 80020 198568
rect 78588 198552 78640 198558
rect 78588 198494 78640 198500
rect 77944 198416 77996 198422
rect 77944 198358 77996 198364
rect 76656 5500 76708 5506
rect 76656 5442 76708 5448
rect 74540 3324 74592 3330
rect 74540 3266 74592 3272
rect 75460 3324 75512 3330
rect 75460 3266 75512 3272
rect 73160 3256 73212 3262
rect 73160 3198 73212 3204
rect 74264 3256 74316 3262
rect 74264 3198 74316 3204
rect 74276 480 74304 3198
rect 75472 480 75500 3266
rect 76668 480 76696 5442
rect 78600 3398 78628 198494
rect 79980 3398 80008 198562
rect 80072 198354 80100 200124
rect 81452 200110 82202 200138
rect 84212 200110 84318 200138
rect 80060 198348 80112 198354
rect 80060 198290 80112 198296
rect 80060 5568 80112 5574
rect 80060 5510 80112 5516
rect 80072 5370 80100 5510
rect 81452 5438 81480 200110
rect 81440 5432 81492 5438
rect 81440 5374 81492 5380
rect 83832 5432 83884 5438
rect 83832 5374 83884 5380
rect 80060 5364 80112 5370
rect 80060 5306 80112 5312
rect 80242 5264 80298 5273
rect 80242 5199 80298 5208
rect 77852 3392 77904 3398
rect 77852 3334 77904 3340
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 79048 3392 79100 3398
rect 79048 3334 79100 3340
rect 79968 3392 80020 3398
rect 79968 3334 80020 3340
rect 77864 480 77892 3334
rect 79060 480 79088 3334
rect 80256 480 80284 5199
rect 82636 4004 82688 4010
rect 82636 3946 82688 3952
rect 81440 3392 81492 3398
rect 81440 3334 81492 3340
rect 81452 480 81480 3334
rect 82648 480 82676 3946
rect 83844 480 83872 5374
rect 84212 4146 84240 200110
rect 85488 198484 85540 198490
rect 85488 198426 85540 198432
rect 85500 4146 85528 198426
rect 86512 198286 86540 200124
rect 86868 198416 86920 198422
rect 86868 198358 86920 198364
rect 86500 198280 86552 198286
rect 86500 198222 86552 198228
rect 86880 4146 86908 198358
rect 88628 198218 88656 200124
rect 89732 200110 90758 200138
rect 92492 200110 92874 200138
rect 88616 198212 88668 198218
rect 88616 198154 88668 198160
rect 89628 110832 89680 110838
rect 89626 110800 89628 110809
rect 89680 110800 89682 110809
rect 89626 110735 89682 110744
rect 89628 87304 89680 87310
rect 89626 87272 89628 87281
rect 89680 87272 89682 87281
rect 89626 87207 89682 87216
rect 89628 76288 89680 76294
rect 89626 76256 89628 76265
rect 89680 76256 89682 76265
rect 89626 76191 89682 76200
rect 88892 63912 88944 63918
rect 88890 63880 88892 63889
rect 88944 63880 88946 63889
rect 88890 63815 88946 63824
rect 88892 40384 88944 40390
rect 88890 40352 88892 40361
rect 88944 40352 88946 40361
rect 88890 40287 88946 40296
rect 89628 29368 89680 29374
rect 89626 29336 89628 29345
rect 89680 29336 89682 29345
rect 89626 29271 89682 29280
rect 89732 5302 89760 200110
rect 92388 198348 92440 198354
rect 92388 198290 92440 198296
rect 92400 193225 92428 198290
rect 92202 193216 92258 193225
rect 92202 193151 92258 193160
rect 92386 193216 92442 193225
rect 92386 193151 92442 193160
rect 92216 183598 92244 193151
rect 92204 183592 92256 183598
rect 92204 183534 92256 183540
rect 92388 183592 92440 183598
rect 92388 183534 92440 183540
rect 92400 173913 92428 183534
rect 92202 173904 92258 173913
rect 92202 173839 92258 173848
rect 92386 173904 92442 173913
rect 92386 173839 92442 173848
rect 92216 164257 92244 173839
rect 92202 164248 92258 164257
rect 92202 164183 92258 164192
rect 92386 164248 92442 164257
rect 92386 164183 92442 164192
rect 92400 154562 92428 164183
rect 92204 154556 92256 154562
rect 92204 154498 92256 154504
rect 92388 154556 92440 154562
rect 92388 154498 92440 154504
rect 92216 144945 92244 154498
rect 92202 144936 92258 144945
rect 92202 144871 92258 144880
rect 92386 144936 92442 144945
rect 92386 144871 92442 144880
rect 92400 135182 92428 144871
rect 92112 135176 92164 135182
rect 92112 135118 92164 135124
rect 92388 135176 92440 135182
rect 92388 135118 92440 135124
rect 92124 125633 92152 135118
rect 92110 125624 92166 125633
rect 92110 125559 92166 125568
rect 92386 125624 92442 125633
rect 92386 125559 92442 125568
rect 92400 115938 92428 125559
rect 92204 115932 92256 115938
rect 92204 115874 92256 115880
rect 92388 115932 92440 115938
rect 92388 115874 92440 115880
rect 92216 106350 92244 115874
rect 92204 106344 92256 106350
rect 92204 106286 92256 106292
rect 92388 106344 92440 106350
rect 92388 106286 92440 106292
rect 92400 96626 92428 106286
rect 92388 96620 92440 96626
rect 92388 96562 92440 96568
rect 92388 87032 92440 87038
rect 92388 86974 92440 86980
rect 92400 57934 92428 86974
rect 92204 57928 92256 57934
rect 92204 57870 92256 57876
rect 92388 57928 92440 57934
rect 92388 57870 92440 57876
rect 92216 48346 92244 57870
rect 92204 48340 92256 48346
rect 92204 48282 92256 48288
rect 92388 48340 92440 48346
rect 92388 48282 92440 48288
rect 92400 38622 92428 48282
rect 92204 38616 92256 38622
rect 92204 38558 92256 38564
rect 92388 38616 92440 38622
rect 92388 38558 92440 38564
rect 92216 29034 92244 38558
rect 92204 29028 92256 29034
rect 92204 28970 92256 28976
rect 92388 29028 92440 29034
rect 92388 28970 92440 28976
rect 92400 19310 92428 28970
rect 92204 19304 92256 19310
rect 92204 19246 92256 19252
rect 92388 19304 92440 19310
rect 92388 19246 92440 19252
rect 92216 9722 92244 19246
rect 92204 9716 92256 9722
rect 92204 9658 92256 9664
rect 92388 9716 92440 9722
rect 92388 9658 92440 9664
rect 91192 5364 91244 5370
rect 91192 5306 91244 5312
rect 89720 5296 89772 5302
rect 91204 5250 91232 5306
rect 89720 5238 89772 5244
rect 90928 5222 91232 5250
rect 87326 5128 87382 5137
rect 87326 5063 87382 5072
rect 84200 4140 84252 4146
rect 84200 4082 84252 4088
rect 84936 4140 84988 4146
rect 84936 4082 84988 4088
rect 85488 4140 85540 4146
rect 85488 4082 85540 4088
rect 86132 4140 86184 4146
rect 86132 4082 86184 4088
rect 86868 4140 86920 4146
rect 86868 4082 86920 4088
rect 86960 4140 87012 4146
rect 86960 4082 87012 4088
rect 84948 480 84976 4082
rect 86144 480 86172 4082
rect 86972 4010 87000 4082
rect 86960 4004 87012 4010
rect 86960 3946 87012 3952
rect 87340 480 87368 5063
rect 88524 4004 88576 4010
rect 88524 3946 88576 3952
rect 88536 480 88564 3946
rect 89718 3768 89774 3777
rect 89718 3703 89774 3712
rect 89732 480 89760 3703
rect 90928 480 90956 5222
rect 92400 3210 92428 9658
rect 92492 4078 92520 200110
rect 93768 198280 93820 198286
rect 93768 198222 93820 198228
rect 92572 96620 92624 96626
rect 92572 96562 92624 96568
rect 92584 87038 92612 96562
rect 92572 87032 92624 87038
rect 92572 86974 92624 86980
rect 93780 4078 93808 198222
rect 94976 198150 95004 200124
rect 94964 198144 95016 198150
rect 94964 198086 95016 198092
rect 97092 198082 97120 200124
rect 98012 200110 99222 200138
rect 100772 200110 101338 200138
rect 102152 200110 103454 200138
rect 97080 198076 97132 198082
rect 97080 198018 97132 198024
rect 96528 110832 96580 110838
rect 96526 110800 96528 110809
rect 96580 110800 96582 110809
rect 96526 110735 96582 110744
rect 96528 87304 96580 87310
rect 96526 87272 96528 87281
rect 96580 87272 96582 87281
rect 96526 87207 96582 87216
rect 96528 76288 96580 76294
rect 96526 76256 96528 76265
rect 96580 76256 96582 76265
rect 96526 76191 96582 76200
rect 96528 63912 96580 63918
rect 96526 63880 96528 63889
rect 96580 63880 96582 63889
rect 96526 63815 96582 63824
rect 96528 40384 96580 40390
rect 96526 40352 96528 40361
rect 96580 40352 96582 40361
rect 96526 40287 96582 40296
rect 96528 29368 96580 29374
rect 96526 29336 96528 29345
rect 96580 29336 96582 29345
rect 96526 29271 96582 29280
rect 98012 5234 98040 200110
rect 99196 198212 99248 198218
rect 99196 198154 99248 198160
rect 98000 5228 98052 5234
rect 98000 5170 98052 5176
rect 98828 5228 98880 5234
rect 98828 5170 98880 5176
rect 94502 4992 94558 5001
rect 94502 4927 94558 4936
rect 92480 4072 92532 4078
rect 92480 4014 92532 4020
rect 93308 4072 93360 4078
rect 93308 4014 93360 4020
rect 93768 4072 93820 4078
rect 93768 4014 93820 4020
rect 92400 3182 92520 3210
rect 92492 610 92520 3182
rect 92112 604 92164 610
rect 92112 546 92164 552
rect 92480 604 92532 610
rect 92480 546 92532 552
rect 92124 480 92152 546
rect 93320 480 93348 4014
rect 94516 480 94544 4927
rect 95700 4004 95752 4010
rect 95700 3946 95752 3952
rect 95712 480 95740 3946
rect 96894 3632 96950 3641
rect 96894 3567 96950 3576
rect 96908 480 96936 3567
rect 98840 2666 98868 5170
rect 98104 2638 98868 2666
rect 98104 480 98132 2638
rect 99208 626 99236 198154
rect 100668 198144 100720 198150
rect 100668 198086 100720 198092
rect 100680 626 100708 198086
rect 100772 3874 100800 200110
rect 101588 6520 101640 6526
rect 101588 6462 101640 6468
rect 100760 3868 100812 3874
rect 100760 3810 100812 3816
rect 99208 598 99328 626
rect 99300 480 99328 598
rect 100496 598 100708 626
rect 100496 480 100524 598
rect 101600 480 101628 6462
rect 102152 3942 102180 200110
rect 105556 198014 105584 200124
rect 107568 198076 107620 198082
rect 107568 198018 107620 198024
rect 105544 198008 105596 198014
rect 105544 197950 105596 197956
rect 107476 198008 107528 198014
rect 107476 197950 107528 197956
rect 103980 5568 104032 5574
rect 103980 5510 104032 5516
rect 103992 5302 104020 5510
rect 104084 5358 104296 5386
rect 103980 5296 104032 5302
rect 103980 5238 104032 5244
rect 104084 5166 104112 5358
rect 104268 5302 104296 5358
rect 104256 5296 104308 5302
rect 104256 5238 104308 5244
rect 106464 5296 106516 5302
rect 106464 5238 106516 5244
rect 104072 5160 104124 5166
rect 104072 5102 104124 5108
rect 106280 5160 106332 5166
rect 106476 5148 106504 5238
rect 106332 5120 106504 5148
rect 106280 5102 106332 5108
rect 105174 4856 105230 4865
rect 105174 4791 105230 4800
rect 102140 3936 102192 3942
rect 102140 3878 102192 3884
rect 102784 3936 102836 3942
rect 102784 3878 102836 3884
rect 102796 480 102824 3878
rect 103980 3868 104032 3874
rect 103980 3810 104032 3816
rect 103992 480 104020 3810
rect 105188 480 105216 4791
rect 106278 4040 106334 4049
rect 106278 3975 106334 3984
rect 106292 3942 106320 3975
rect 106280 3936 106332 3942
rect 106280 3878 106332 3884
rect 106372 3936 106424 3942
rect 106372 3878 106424 3884
rect 106384 480 106412 3878
rect 107488 3788 107516 197950
rect 107580 3942 107608 198018
rect 107672 5234 107700 200124
rect 109052 200110 109894 200138
rect 111812 200110 112010 200138
rect 113192 200110 114126 200138
rect 115952 200110 116242 200138
rect 117332 200110 118358 200138
rect 120092 200110 120474 200138
rect 121472 200110 122590 200138
rect 124232 200110 124706 200138
rect 125612 200110 126822 200138
rect 128464 200110 128938 200138
rect 130304 200110 131054 200138
rect 132512 200110 133262 200138
rect 108764 6452 108816 6458
rect 108764 6394 108816 6400
rect 107660 5228 107712 5234
rect 107660 5170 107712 5176
rect 107568 3936 107620 3942
rect 107568 3878 107620 3884
rect 107488 3760 107608 3788
rect 107580 480 107608 3760
rect 108776 480 108804 6394
rect 109052 3806 109080 200110
rect 109408 5568 109460 5574
rect 109408 5510 109460 5516
rect 109420 5166 109448 5510
rect 109408 5160 109460 5166
rect 109408 5102 109460 5108
rect 109040 3800 109092 3806
rect 109040 3742 109092 3748
rect 109776 3800 109828 3806
rect 109776 3742 109828 3748
rect 109788 3602 109816 3742
rect 111812 3738 111840 200110
rect 112352 6384 112404 6390
rect 112352 6326 112404 6332
rect 111800 3732 111852 3738
rect 111800 3674 111852 3680
rect 109776 3596 109828 3602
rect 109776 3538 109828 3544
rect 111154 3496 111210 3505
rect 111154 3431 111210 3440
rect 109960 1964 110012 1970
rect 109960 1906 110012 1912
rect 109972 480 110000 1906
rect 111168 480 111196 3431
rect 112364 480 112392 6326
rect 113192 5030 113220 200110
rect 115846 198112 115902 198121
rect 115846 198047 115902 198056
rect 115860 5030 115888 198047
rect 113180 5024 113232 5030
rect 113180 4966 113232 4972
rect 114744 5024 114796 5030
rect 114744 4966 114796 4972
rect 115848 5024 115900 5030
rect 115848 4966 115900 4972
rect 114650 3904 114706 3913
rect 114650 3839 114706 3848
rect 114664 3806 114692 3839
rect 114652 3800 114704 3806
rect 114652 3742 114704 3748
rect 113548 3732 113600 3738
rect 113548 3674 113600 3680
rect 113560 480 113588 3674
rect 114756 480 114784 4966
rect 115662 4040 115718 4049
rect 115662 3975 115718 3984
rect 115676 3942 115704 3975
rect 115664 3936 115716 3942
rect 115664 3878 115716 3884
rect 115848 3800 115900 3806
rect 115848 3742 115900 3748
rect 115860 1970 115888 3742
rect 115952 3602 115980 200110
rect 117226 197976 117282 197985
rect 117226 197911 117282 197920
rect 116032 110560 116084 110566
rect 116030 110528 116032 110537
rect 116084 110528 116086 110537
rect 116030 110463 116086 110472
rect 116032 87032 116084 87038
rect 116030 87000 116032 87009
rect 116084 87000 116086 87009
rect 116030 86935 116086 86944
rect 116032 76016 116084 76022
rect 116030 75984 116032 75993
rect 116084 75984 116086 75993
rect 116030 75919 116086 75928
rect 116032 63640 116084 63646
rect 116030 63608 116032 63617
rect 116084 63608 116086 63617
rect 116030 63543 116086 63552
rect 116032 40112 116084 40118
rect 116030 40080 116032 40089
rect 116084 40080 116086 40089
rect 116030 40015 116086 40024
rect 116032 29096 116084 29102
rect 116030 29064 116032 29073
rect 116084 29064 116086 29073
rect 116030 28999 116086 29008
rect 116124 6316 116176 6322
rect 116124 6258 116176 6264
rect 115940 3596 115992 3602
rect 115940 3538 115992 3544
rect 116136 3482 116164 6258
rect 115952 3454 116164 3482
rect 115848 1964 115900 1970
rect 115848 1906 115900 1912
rect 115952 480 115980 3454
rect 117240 626 117268 197911
rect 117332 3913 117360 200110
rect 118790 110800 118846 110809
rect 118790 110735 118846 110744
rect 118804 110566 118832 110735
rect 118792 110560 118844 110566
rect 118792 110502 118844 110508
rect 118790 76256 118846 76265
rect 118790 76191 118846 76200
rect 118804 76022 118832 76191
rect 118792 76016 118844 76022
rect 118792 75958 118844 75964
rect 118790 63880 118846 63889
rect 118790 63815 118846 63824
rect 118804 63646 118832 63815
rect 118792 63640 118844 63646
rect 118792 63582 118844 63588
rect 118790 40352 118846 40361
rect 118790 40287 118846 40296
rect 118804 40118 118832 40287
rect 118792 40112 118844 40118
rect 118792 40054 118844 40060
rect 119436 6248 119488 6254
rect 119436 6190 119488 6196
rect 118528 5222 118832 5250
rect 118528 5098 118556 5222
rect 118608 5160 118660 5166
rect 118608 5102 118660 5108
rect 118516 5092 118568 5098
rect 118516 5034 118568 5040
rect 118620 4978 118648 5102
rect 118804 5098 118832 5222
rect 118792 5092 118844 5098
rect 118792 5034 118844 5040
rect 118884 5024 118936 5030
rect 118620 4972 118884 4978
rect 118620 4966 118936 4972
rect 118620 4950 118924 4966
rect 117318 3904 117374 3913
rect 117318 3839 117374 3848
rect 118240 3664 118292 3670
rect 118240 3606 118292 3612
rect 117148 598 117268 626
rect 117148 480 117176 598
rect 118252 480 118280 3606
rect 119448 480 119476 6190
rect 120092 4962 120120 200110
rect 120814 87272 120870 87281
rect 120814 87207 120870 87216
rect 120828 87038 120856 87207
rect 120816 87032 120868 87038
rect 120816 86974 120868 86980
rect 120814 29336 120870 29345
rect 120814 29271 120870 29280
rect 120828 29102 120856 29271
rect 120816 29096 120868 29102
rect 120816 29038 120868 29044
rect 120080 4956 120132 4962
rect 120080 4898 120132 4904
rect 120632 3596 120684 3602
rect 120632 3538 120684 3544
rect 120644 480 120672 3538
rect 121472 3534 121500 200110
rect 123024 6180 123076 6186
rect 123024 6122 123076 6128
rect 121460 3528 121512 3534
rect 121460 3470 121512 3476
rect 121828 3528 121880 3534
rect 121828 3470 121880 3476
rect 121840 480 121868 3470
rect 123036 480 123064 6122
rect 124232 3618 124260 200110
rect 125612 4894 125640 200110
rect 127624 197396 127676 197402
rect 127624 197338 127676 197344
rect 126612 5228 126664 5234
rect 126612 5170 126664 5176
rect 125600 4888 125652 4894
rect 125600 4830 125652 4836
rect 124140 3590 124260 3618
rect 124140 3466 124168 3590
rect 124128 3460 124180 3466
rect 124128 3402 124180 3408
rect 124220 3460 124272 3466
rect 124220 3402 124272 3408
rect 124232 480 124260 3402
rect 125414 3360 125470 3369
rect 125414 3295 125470 3304
rect 125428 480 125456 3295
rect 126624 480 126652 5170
rect 127636 5030 127664 197338
rect 128174 87272 128230 87281
rect 128358 87272 128414 87281
rect 128230 87230 128358 87258
rect 128174 87207 128230 87216
rect 128358 87207 128414 87216
rect 128174 29336 128230 29345
rect 128358 29336 128414 29345
rect 128230 29294 128358 29322
rect 128174 29271 128230 29280
rect 128358 29271 128414 29280
rect 127808 5160 127860 5166
rect 127808 5102 127860 5108
rect 127624 5024 127676 5030
rect 127624 4966 127676 4972
rect 127820 480 127848 5102
rect 128464 2854 128492 200110
rect 130304 197470 130332 200110
rect 130292 197464 130344 197470
rect 130292 197406 130344 197412
rect 130384 197464 130436 197470
rect 130384 197406 130436 197412
rect 130396 5098 130424 197406
rect 130384 5092 130436 5098
rect 130384 5034 130436 5040
rect 130200 5024 130252 5030
rect 130200 4966 130252 4972
rect 129004 4956 129056 4962
rect 129004 4898 129056 4904
rect 128452 2848 128504 2854
rect 128452 2790 128504 2796
rect 129016 480 129044 4898
rect 130212 480 130240 4966
rect 131396 4956 131448 4962
rect 131396 4898 131448 4904
rect 131408 480 131436 4898
rect 132512 4826 132540 200110
rect 135364 197538 135392 200124
rect 136652 200110 137494 200138
rect 139412 200110 139610 200138
rect 140792 200110 141726 200138
rect 135352 197532 135404 197538
rect 135352 197474 135404 197480
rect 135166 111072 135222 111081
rect 135166 111007 135222 111016
rect 135180 110673 135208 111007
rect 135166 110664 135222 110673
rect 135166 110599 135222 110608
rect 135166 76528 135222 76537
rect 135166 76463 135222 76472
rect 135180 76129 135208 76463
rect 135166 76120 135222 76129
rect 135166 76055 135222 76064
rect 135166 64152 135222 64161
rect 135166 64087 135222 64096
rect 135180 63753 135208 64087
rect 135166 63744 135222 63753
rect 135166 63679 135222 63688
rect 135166 40624 135222 40633
rect 135166 40559 135222 40568
rect 135180 40225 135208 40559
rect 135166 40216 135222 40225
rect 135166 40151 135222 40160
rect 134892 4888 134944 4894
rect 134892 4830 134944 4836
rect 132500 4820 132552 4826
rect 132500 4762 132552 4768
rect 132592 4820 132644 4826
rect 132592 4762 132644 4768
rect 132604 480 132632 4762
rect 134904 480 134932 4830
rect 136652 2922 136680 200110
rect 139412 4214 139440 200110
rect 140042 110936 140098 110945
rect 140042 110871 140098 110880
rect 140056 110537 140084 110871
rect 140042 110528 140098 110537
rect 140042 110463 140098 110472
rect 140042 76392 140098 76401
rect 140042 76327 140098 76336
rect 140056 75993 140084 76327
rect 140042 75984 140098 75993
rect 140042 75919 140098 75928
rect 140042 64016 140098 64025
rect 140042 63951 140098 63960
rect 140056 63617 140084 63951
rect 140042 63608 140098 63617
rect 140042 63543 140098 63552
rect 140042 40488 140098 40497
rect 140042 40423 140098 40432
rect 140056 40089 140084 40423
rect 140042 40080 140098 40089
rect 140042 40015 140098 40024
rect 139400 4208 139452 4214
rect 139400 4150 139452 4156
rect 140792 2990 140820 200110
rect 143828 197606 143856 200124
rect 144932 200110 145958 200138
rect 143816 197600 143868 197606
rect 143816 197542 143868 197548
rect 143446 87408 143502 87417
rect 143446 87343 143502 87352
rect 143460 87009 143488 87343
rect 143446 87000 143502 87009
rect 143446 86935 143502 86944
rect 143446 29472 143502 29481
rect 143446 29407 143502 29416
rect 143460 29073 143488 29407
rect 143446 29064 143502 29073
rect 143446 28999 143502 29008
rect 144932 4282 144960 200110
rect 148060 197470 148088 200124
rect 150176 197674 150204 200124
rect 151832 200110 152306 200138
rect 153212 200110 154422 200138
rect 150164 197668 150216 197674
rect 150164 197610 150216 197616
rect 148048 197464 148100 197470
rect 148048 197406 148100 197412
rect 147588 110696 147640 110702
rect 147586 110664 147588 110673
rect 147640 110664 147642 110673
rect 147586 110599 147642 110608
rect 145564 87168 145616 87174
rect 145564 87110 145616 87116
rect 145576 87009 145604 87110
rect 145562 87000 145618 87009
rect 145562 86935 145618 86944
rect 147588 76152 147640 76158
rect 147586 76120 147588 76129
rect 147640 76120 147642 76129
rect 147586 76055 147642 76064
rect 147588 63776 147640 63782
rect 147586 63744 147588 63753
rect 147640 63744 147642 63753
rect 147586 63679 147642 63688
rect 147588 40248 147640 40254
rect 147586 40216 147588 40225
rect 147640 40216 147642 40225
rect 147586 40151 147642 40160
rect 145012 29096 145064 29102
rect 145010 29064 145012 29073
rect 145064 29064 145066 29073
rect 145010 28999 145066 29008
rect 151832 4350 151860 200110
rect 153212 6730 153240 200110
rect 156524 197742 156552 200124
rect 156512 197736 156564 197742
rect 156512 197678 156564 197684
rect 154486 110800 154542 110809
rect 154486 110735 154542 110744
rect 154500 110702 154528 110735
rect 154488 110696 154540 110702
rect 154488 110638 154540 110644
rect 154486 87272 154542 87281
rect 154486 87207 154542 87216
rect 154500 87174 154528 87207
rect 154488 87168 154540 87174
rect 154488 87110 154540 87116
rect 154486 76256 154542 76265
rect 154486 76191 154542 76200
rect 154500 76158 154528 76191
rect 154488 76152 154540 76158
rect 154488 76094 154540 76100
rect 154486 63880 154542 63889
rect 154486 63815 154542 63824
rect 154500 63782 154528 63815
rect 154488 63776 154540 63782
rect 154488 63718 154540 63724
rect 154486 40352 154542 40361
rect 154486 40287 154542 40296
rect 154500 40254 154528 40287
rect 154488 40248 154540 40254
rect 154488 40190 154540 40196
rect 154486 29336 154542 29345
rect 154486 29271 154542 29280
rect 154500 29102 154528 29271
rect 154488 29096 154540 29102
rect 154488 29038 154540 29044
rect 153200 6724 153252 6730
rect 153200 6666 153252 6672
rect 158732 4418 158760 200124
rect 160848 197402 160876 200124
rect 162964 197810 162992 200124
rect 164252 200110 165094 200138
rect 167012 200110 167210 200138
rect 168392 200110 169326 200138
rect 171152 200110 171442 200138
rect 172532 200110 173558 200138
rect 162952 197804 163004 197810
rect 162952 197746 163004 197752
rect 160836 197396 160888 197402
rect 160836 197338 160888 197344
rect 164252 4486 164280 200110
rect 167012 6662 167040 200110
rect 167000 6656 167052 6662
rect 167000 6598 167052 6604
rect 164240 4480 164292 4486
rect 164240 4422 164292 4428
rect 158720 4412 158772 4418
rect 158720 4354 158772 4360
rect 151820 4344 151872 4350
rect 151820 4286 151872 4292
rect 144920 4276 144972 4282
rect 144920 4218 144972 4224
rect 168392 3058 168420 200110
rect 171152 4554 171180 200110
rect 172532 6594 172560 200110
rect 175660 197878 175688 200124
rect 176672 200110 177790 200138
rect 179432 200110 179906 200138
rect 180812 200110 182114 200138
rect 183572 200110 184230 200138
rect 175648 197872 175700 197878
rect 175648 197814 175700 197820
rect 172520 6588 172572 6594
rect 172520 6530 172572 6536
rect 176672 4622 176700 200110
rect 176660 4616 176712 4622
rect 176660 4558 176712 4564
rect 171140 4548 171192 4554
rect 171140 4490 171192 4496
rect 179432 3126 179460 200110
rect 180812 3194 180840 200110
rect 183572 4690 183600 200110
rect 186332 198694 186360 200124
rect 186320 198688 186372 198694
rect 186320 198630 186372 198636
rect 188448 197946 188476 200124
rect 190472 200110 190578 200138
rect 191852 200110 192694 200138
rect 194612 200110 194810 200138
rect 195992 200110 196926 200138
rect 188436 197940 188488 197946
rect 188436 197882 188488 197888
rect 190472 4758 190500 200110
rect 190460 4752 190512 4758
rect 190460 4694 190512 4700
rect 183560 4684 183612 4690
rect 183560 4626 183612 4632
rect 191852 3262 191880 200110
rect 194612 3330 194640 200110
rect 195992 5506 196020 200110
rect 199028 198558 199056 200124
rect 201144 198626 201172 200124
rect 202892 200110 203274 200138
rect 204272 200110 205482 200138
rect 207032 200110 207598 200138
rect 208412 200110 209714 200138
rect 201132 198620 201184 198626
rect 201132 198562 201184 198568
rect 199016 198552 199068 198558
rect 199016 198494 199068 198500
rect 195980 5500 196032 5506
rect 195980 5442 196032 5448
rect 202892 5273 202920 200110
rect 202878 5264 202934 5273
rect 202878 5199 202934 5208
rect 204272 3398 204300 200110
rect 207032 4146 207060 200110
rect 208412 5438 208440 200110
rect 211816 198490 211844 200124
rect 211804 198484 211856 198490
rect 211804 198426 211856 198432
rect 213932 198422 213960 200124
rect 215312 200110 216062 200138
rect 218072 200110 218178 200138
rect 219452 200110 220294 200138
rect 222212 200110 222410 200138
rect 213920 198416 213972 198422
rect 213920 198358 213972 198364
rect 208400 5432 208452 5438
rect 208400 5374 208452 5380
rect 215312 5137 215340 200110
rect 215298 5128 215354 5137
rect 215298 5063 215354 5072
rect 207020 4140 207072 4146
rect 207020 4082 207072 4088
rect 218072 4078 218100 200110
rect 218060 4072 218112 4078
rect 218060 4014 218112 4020
rect 219452 3777 219480 200110
rect 222212 5370 222240 200110
rect 224512 198354 224540 200124
rect 224500 198348 224552 198354
rect 224500 198290 224552 198296
rect 226628 198286 226656 200124
rect 227732 200110 228758 200138
rect 230492 200110 230966 200138
rect 231872 200110 233082 200138
rect 234632 200110 235198 200138
rect 226616 198280 226668 198286
rect 226616 198222 226668 198228
rect 222200 5364 222252 5370
rect 222200 5306 222252 5312
rect 227732 5001 227760 200110
rect 227718 4992 227774 5001
rect 227718 4927 227774 4936
rect 230492 4010 230520 200110
rect 230480 4004 230532 4010
rect 230480 3946 230532 3952
rect 219438 3768 219494 3777
rect 219438 3703 219494 3712
rect 231872 3641 231900 200110
rect 234632 5302 234660 200110
rect 237300 198218 237328 200124
rect 237288 198212 237340 198218
rect 237288 198154 237340 198160
rect 239416 198150 239444 200124
rect 239404 198144 239456 198150
rect 239404 198086 239456 198092
rect 241532 6526 241560 200124
rect 242912 200110 243662 200138
rect 245672 200110 245778 200138
rect 247052 200110 247894 200138
rect 241520 6520 241572 6526
rect 241520 6462 241572 6468
rect 234620 5296 234672 5302
rect 234620 5238 234672 5244
rect 242912 3942 242940 200110
rect 242900 3936 242952 3942
rect 242900 3878 242952 3884
rect 245672 3874 245700 200110
rect 247052 4865 247080 200110
rect 249996 198082 250024 200124
rect 249984 198076 250036 198082
rect 249984 198018 250036 198024
rect 252112 198014 252140 200124
rect 253952 200110 254334 200138
rect 255332 200110 256450 200138
rect 258092 200110 258566 200138
rect 259472 200110 260682 200138
rect 262232 200110 262798 200138
rect 252100 198008 252152 198014
rect 252100 197950 252152 197956
rect 253952 6458 253980 200110
rect 253940 6452 253992 6458
rect 253940 6394 253992 6400
rect 247038 4856 247094 4865
rect 247038 4791 247094 4800
rect 245660 3868 245712 3874
rect 245660 3810 245712 3816
rect 255332 3806 255360 200110
rect 255320 3800 255372 3806
rect 255320 3742 255372 3748
rect 231858 3632 231914 3641
rect 231858 3567 231914 3576
rect 258092 3505 258120 200110
rect 259472 6390 259500 200110
rect 259460 6384 259512 6390
rect 259460 6326 259512 6332
rect 262232 3738 262260 200110
rect 264900 198121 264928 200124
rect 266372 200110 267030 200138
rect 264886 198112 264942 198121
rect 264886 198047 264942 198056
rect 266372 6322 266400 200110
rect 269132 197985 269160 200124
rect 270512 200110 271262 200138
rect 273272 200110 273378 200138
rect 274652 200110 275494 200138
rect 277412 200110 277702 200138
rect 278792 200110 279818 200138
rect 281552 200110 281934 200138
rect 282932 200110 284050 200138
rect 285692 200110 286166 200138
rect 287072 200110 288282 200138
rect 289832 200110 290398 200138
rect 291212 200110 292514 200138
rect 293972 200110 294630 200138
rect 269118 197976 269174 197985
rect 269118 197911 269174 197920
rect 266360 6316 266412 6322
rect 266360 6258 266412 6264
rect 262220 3732 262272 3738
rect 262220 3674 262272 3680
rect 270512 3670 270540 200110
rect 273272 6254 273300 200110
rect 273260 6248 273312 6254
rect 273260 6190 273312 6196
rect 270500 3664 270552 3670
rect 270500 3606 270552 3612
rect 274652 3602 274680 200110
rect 274640 3596 274692 3602
rect 274640 3538 274692 3544
rect 277412 3534 277440 200110
rect 278792 6186 278820 200110
rect 278780 6180 278832 6186
rect 278780 6122 278832 6128
rect 277400 3528 277452 3534
rect 258078 3496 258134 3505
rect 277400 3470 277452 3476
rect 281552 3466 281580 200110
rect 258078 3431 258134 3440
rect 281540 3460 281592 3466
rect 281540 3402 281592 3408
rect 204260 3392 204312 3398
rect 282932 3369 282960 200110
rect 285692 5234 285720 200110
rect 285680 5228 285732 5234
rect 285680 5170 285732 5176
rect 287072 5166 287100 200110
rect 287060 5160 287112 5166
rect 287060 5102 287112 5108
rect 289832 5030 289860 200110
rect 291212 5098 291240 200110
rect 291200 5092 291252 5098
rect 291200 5034 291252 5040
rect 289820 5024 289872 5030
rect 289820 4966 289872 4972
rect 293972 4962 294000 200110
rect 293960 4956 294012 4962
rect 293960 4898 294012 4904
rect 296732 4826 296760 200124
rect 298112 200110 298862 200138
rect 298112 4894 298140 200110
rect 580460 199918 580488 346015
rect 580538 322688 580594 322697
rect 580538 322623 580594 322632
rect 580552 200734 580580 322623
rect 580630 310856 580686 310865
rect 580630 310791 580686 310800
rect 580540 200728 580592 200734
rect 580540 200670 580592 200676
rect 580644 199986 580672 310791
rect 580722 299160 580778 299169
rect 580722 299095 580778 299104
rect 580736 200122 580764 299095
rect 580814 275768 580870 275777
rect 580814 275703 580870 275712
rect 580828 200870 580856 275703
rect 580906 263936 580962 263945
rect 580906 263871 580962 263880
rect 580816 200864 580868 200870
rect 580816 200806 580868 200812
rect 580724 200116 580776 200122
rect 580724 200058 580776 200064
rect 580920 200054 580948 263871
rect 580908 200048 580960 200054
rect 580908 199990 580960 199996
rect 580632 199980 580684 199986
rect 580632 199922 580684 199928
rect 580448 199912 580500 199918
rect 580448 199854 580500 199860
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 298100 4888 298152 4894
rect 298100 4830 298152 4836
rect 296720 4820 296772 4826
rect 296720 4762 296772 4768
rect 204260 3334 204312 3340
rect 282918 3360 282974 3369
rect 194600 3324 194652 3330
rect 282918 3295 282974 3304
rect 194600 3266 194652 3272
rect 191840 3256 191892 3262
rect 191840 3198 191892 3204
rect 180800 3188 180852 3194
rect 180800 3130 180852 3136
rect 179420 3120 179472 3126
rect 179420 3062 179472 3068
rect 168380 3052 168432 3058
rect 168380 2994 168432 3000
rect 140780 2984 140832 2990
rect 140780 2926 140832 2932
rect 136640 2916 136692 2922
rect 136640 2858 136692 2864
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 4802 682216 4858 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 4066 624824 4122 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 3422 567296 3478 567352
rect 3146 553016 3202 553072
rect 2962 481072 3018 481128
rect 3330 437960 3386 438016
rect 3146 423680 3202 423736
rect 2778 394984 2834 395040
rect 3054 366152 3110 366208
rect 3330 380568 3386 380624
rect 3606 538600 3662 538656
rect 3238 337456 3294 337512
rect 3054 294344 3110 294400
rect 3422 280100 3424 280120
rect 3424 280100 3476 280120
rect 3476 280100 3478 280120
rect 3422 280064 3478 280100
rect 2778 265648 2834 265704
rect 3422 251232 3478 251288
rect 3422 236952 3478 237008
rect 2778 222536 2834 222592
rect 3698 509904 3754 509960
rect 3790 495488 3846 495544
rect 3974 452376 4030 452432
rect 4066 323040 4122 323096
rect 3882 308760 3938 308816
rect 3514 208120 3570 208176
rect 3146 193840 3202 193896
rect 3238 179424 3294 179480
rect 2778 165008 2834 165064
rect 3146 150728 3202 150784
rect 3238 136312 3294 136368
rect 2778 122032 2834 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 3422 78920 3478 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 3422 7112 3478 7168
rect 19338 384820 19340 384840
rect 19340 384820 19392 384840
rect 19392 384820 19394 384840
rect 19338 384784 19394 384820
rect 22098 384784 22154 384840
rect 38658 384940 38714 384976
rect 38658 384920 38660 384940
rect 38660 384920 38712 384940
rect 38712 384920 38714 384940
rect 57518 546488 57574 546544
rect 57426 545128 57482 545184
rect 56874 543768 56930 543824
rect 56782 540368 56838 540424
rect 57334 542408 57390 542464
rect 57150 539552 57206 539608
rect 57058 537512 57114 537568
rect 56966 480256 57022 480312
rect 56874 442448 56930 442504
rect 57426 442312 57482 442368
rect 57518 442176 57574 442232
rect 56598 438932 56654 438968
rect 56598 438912 56600 438932
rect 56600 438912 56652 438932
rect 56652 438912 56654 438932
rect 42890 384940 42946 384976
rect 42890 384920 42892 384940
rect 42892 384920 42944 384940
rect 42944 384920 42946 384940
rect 56598 436092 56600 436112
rect 56600 436092 56652 436112
rect 56652 436092 56654 436112
rect 56598 436056 56654 436092
rect 56506 394732 56562 394768
rect 56506 394712 56508 394732
rect 56508 394712 56560 394732
rect 56560 394712 56562 394732
rect 56690 434732 56692 434752
rect 56692 434732 56744 434752
rect 56744 434732 56746 434752
rect 56690 434696 56746 434732
rect 56690 431996 56746 432032
rect 56690 431976 56692 431996
rect 56692 431976 56744 431996
rect 56744 431976 56746 431996
rect 56690 400968 56746 401024
rect 56690 398928 56746 398984
rect 56690 396752 56746 396808
rect 56598 392536 56654 392592
rect 56598 390496 56654 390552
rect 56598 387776 56654 387832
rect 56598 387640 56654 387696
rect 56598 386280 56654 386336
rect 56598 384104 56654 384160
rect 56598 382064 56654 382120
rect 56598 380024 56654 380080
rect 56598 377848 56654 377904
rect 56598 375808 56654 375864
rect 56598 373632 56654 373688
rect 56598 371592 56654 371648
rect 56598 369416 56654 369472
rect 56598 367376 56654 367432
rect 56598 365200 56654 365256
rect 56598 363160 56654 363216
rect 56598 360984 56654 361040
rect 56598 358944 56654 359000
rect 56598 356768 56654 356824
rect 56598 354728 56654 354784
rect 56598 352552 56654 352608
rect 56598 350512 56654 350568
rect 56598 348336 56654 348392
rect 56598 346332 56600 346352
rect 56600 346332 56652 346352
rect 56652 346332 56654 346352
rect 56598 346296 56654 346332
rect 56782 327256 56838 327312
rect 56874 321000 56930 321056
rect 56966 314744 57022 314800
rect 57150 430480 57206 430536
rect 57150 428440 57206 428496
rect 57150 426264 57206 426320
rect 57150 424224 57206 424280
rect 57150 422048 57206 422104
rect 57150 420008 57206 420064
rect 57150 417832 57206 417888
rect 57150 415792 57206 415848
rect 57150 413616 57206 413672
rect 57150 411576 57206 411632
rect 57150 409400 57206 409456
rect 57150 407360 57206 407416
rect 57150 405184 57206 405240
rect 57150 403144 57206 403200
rect 57058 308352 57114 308408
rect 57242 268368 57298 268424
rect 57334 259936 57390 259992
rect 57426 253680 57482 253736
rect 57702 333648 57758 333704
rect 57794 331472 57850 331528
rect 57610 261976 57666 262032
rect 57886 318960 57942 319016
rect 57978 270408 58034 270464
rect 58162 439320 58218 439376
rect 58070 264152 58126 264208
rect 58438 344120 58494 344176
rect 58530 342080 58586 342136
rect 58622 337864 58678 337920
rect 58714 335688 58770 335744
rect 58806 329432 58862 329488
rect 58898 323040 58954 323096
rect 58990 316784 59046 316840
rect 59082 312568 59138 312624
rect 59174 310528 59230 310584
rect 59266 304136 59322 304192
rect 59542 339904 59598 339960
rect 59450 325216 59506 325272
rect 59358 293664 59414 293720
rect 59726 603336 59782 603392
rect 59726 596264 59782 596320
rect 59634 287272 59690 287328
rect 59818 579536 59874 579592
rect 59818 570152 59874 570208
rect 133694 553444 133750 553480
rect 133694 553424 133696 553444
rect 133696 553424 133748 553444
rect 133748 553424 133750 553444
rect 59818 478527 59874 478583
rect 77298 459448 77354 459504
rect 74170 458088 74226 458144
rect 75826 458088 75882 458144
rect 79966 458108 80022 458144
rect 79966 458088 79968 458108
rect 79968 458088 80020 458108
rect 80020 458088 80022 458108
rect 73066 457700 73122 457736
rect 73066 457680 73068 457700
rect 73068 457680 73120 457700
rect 73120 457680 73122 457700
rect 81898 458088 81954 458144
rect 82818 458088 82874 458144
rect 84198 458088 84254 458144
rect 85486 458088 85542 458144
rect 86314 458124 86316 458144
rect 86316 458124 86368 458144
rect 86368 458124 86370 458144
rect 86314 458088 86370 458124
rect 81346 457952 81402 458008
rect 78586 457836 78642 457872
rect 78586 457816 78588 457836
rect 78588 457816 78640 457836
rect 78640 457816 78642 457836
rect 63682 457544 63738 457600
rect 77206 457564 77262 457600
rect 87878 458088 87934 458144
rect 89074 458108 89130 458144
rect 89074 458088 89076 458108
rect 89076 458088 89128 458108
rect 89128 458088 89130 458108
rect 90178 458088 90234 458144
rect 91098 458108 91154 458144
rect 91098 458088 91100 458108
rect 91100 458088 91152 458108
rect 91152 458088 91154 458108
rect 92478 458088 92534 458144
rect 93582 458088 93638 458144
rect 94778 458088 94834 458144
rect 95790 458088 95846 458144
rect 97170 458088 97226 458144
rect 98550 458088 98606 458144
rect 99470 458088 99526 458144
rect 100666 458088 100722 458144
rect 101954 458088 102010 458144
rect 102782 458088 102838 458144
rect 103426 458088 103482 458144
rect 104254 458088 104310 458144
rect 104806 458088 104862 458144
rect 105358 458124 105360 458144
rect 105360 458124 105412 458144
rect 105412 458124 105414 458144
rect 105358 458088 105414 458124
rect 106186 458088 106242 458144
rect 107566 458088 107622 458144
rect 100574 457952 100630 458008
rect 77206 457544 77208 457564
rect 77208 457544 77260 457564
rect 77260 457544 77262 457564
rect 59726 281016 59782 281072
rect 58346 276800 58402 276856
rect 58254 272584 58310 272640
rect 58162 257896 58218 257952
rect 57794 255720 57850 255776
rect 57518 251504 57574 251560
rect 57886 245248 57942 245304
rect 56874 243072 56930 243128
rect 56782 219952 56838 220008
rect 56690 217776 56746 217832
rect 56598 215736 56654 215792
rect 57702 241032 57758 241088
rect 57242 238856 57298 238912
rect 57150 234640 57206 234696
rect 56966 232600 57022 232656
rect 57058 230424 57114 230480
rect 57610 236816 57666 236872
rect 57518 226208 57574 226264
rect 57426 224168 57482 224224
rect 57334 221992 57390 222048
rect 57794 228384 57850 228440
rect 57794 201048 57850 201104
rect 59818 204992 59874 205048
rect 73158 457408 73214 457464
rect 75918 457408 75974 457464
rect 71778 457136 71834 457192
rect 70214 457000 70270 457056
rect 67546 456864 67602 456920
rect 68834 456864 68890 456920
rect 70122 456864 70178 456920
rect 71686 456864 71742 456920
rect 74722 457000 74778 457056
rect 77298 457136 77354 457192
rect 95146 457136 95202 457192
rect 99286 457136 99342 457192
rect 78770 457000 78826 457056
rect 93766 457000 93822 457056
rect 78678 456864 78734 456920
rect 80058 456864 80114 456920
rect 81438 456864 81494 456920
rect 82818 456864 82874 456920
rect 84198 456864 84254 456920
rect 86222 456864 86278 456920
rect 86866 456864 86922 456920
rect 88246 456864 88302 456920
rect 89626 456864 89682 456920
rect 91006 456864 91062 456920
rect 92386 456864 92442 456920
rect 93674 456864 93730 456920
rect 96526 456864 96582 456920
rect 97906 456864 97962 456920
rect 101862 457816 101918 457872
rect 102046 457952 102102 458008
rect 106278 457988 106280 458008
rect 106280 457988 106332 458008
rect 106332 457988 106334 458008
rect 106278 457952 106334 457988
rect 108762 458088 108818 458144
rect 110326 458088 110382 458144
rect 107658 457952 107714 458008
rect 108946 457952 109002 458008
rect 478510 700712 478566 700768
rect 494794 700576 494850 700632
rect 527178 700440 527234 700496
rect 543462 700304 543518 700360
rect 289818 673804 289874 673840
rect 289818 673784 289820 673804
rect 289820 673784 289872 673804
rect 289872 673784 289874 673804
rect 292670 673512 292726 673568
rect 580170 697992 580226 698048
rect 580170 686296 580226 686352
rect 553306 673920 553362 673976
rect 553490 673920 553546 673976
rect 540978 673804 541034 673840
rect 540978 673784 540980 673804
rect 540980 673784 541032 673804
rect 541032 673784 541034 673804
rect 548614 673512 548670 673568
rect 425058 650276 425114 650312
rect 425058 650256 425060 650276
rect 425060 650256 425112 650276
rect 425112 650256 425114 650276
rect 560298 673940 560354 673976
rect 560298 673920 560300 673940
rect 560300 673920 560352 673940
rect 560352 673920 560354 673940
rect 565174 673784 565230 673840
rect 572718 673784 572774 673840
rect 572626 673648 572682 673704
rect 553306 650392 553362 650448
rect 553490 650392 553546 650448
rect 540978 650276 541034 650312
rect 540978 650256 540980 650276
rect 540980 650256 541032 650276
rect 541032 650256 541034 650276
rect 434534 650120 434590 650176
rect 548614 649984 548670 650040
rect 560298 650412 560354 650448
rect 560298 650392 560300 650412
rect 560300 650392 560352 650412
rect 560352 650392 560354 650412
rect 565174 650256 565230 650312
rect 572718 650256 572774 650312
rect 572626 650120 572682 650176
rect 580170 639376 580226 639432
rect 289818 626884 289874 626920
rect 289818 626864 289820 626884
rect 289820 626864 289872 626884
rect 289872 626864 289874 626884
rect 292670 626592 292726 626648
rect 425058 626884 425114 626920
rect 425058 626864 425060 626884
rect 425060 626864 425112 626884
rect 425112 626864 425114 626884
rect 427910 626592 427966 626648
rect 553306 627000 553362 627056
rect 553490 627000 553546 627056
rect 540978 626884 541034 626920
rect 540978 626864 540980 626884
rect 540980 626864 541032 626884
rect 541032 626864 541034 626884
rect 548614 626592 548670 626648
rect 560298 627020 560354 627056
rect 560298 627000 560300 627020
rect 560300 627000 560352 627020
rect 560352 627000 560354 627020
rect 565174 626864 565230 626920
rect 572718 626864 572774 626920
rect 572626 626728 572682 626784
rect 289818 603356 289874 603392
rect 289818 603336 289820 603356
rect 289820 603336 289872 603356
rect 289872 603336 289874 603356
rect 292670 603064 292726 603120
rect 559102 608640 559158 608696
rect 559378 608640 559434 608696
rect 425058 603356 425114 603392
rect 425058 603336 425060 603356
rect 425060 603336 425112 603356
rect 425112 603336 425114 603356
rect 553398 603472 553454 603528
rect 441526 603336 441582 603392
rect 540978 603356 541034 603392
rect 540978 603336 540980 603356
rect 540980 603336 541032 603356
rect 541032 603336 541034 603356
rect 429934 603200 429990 603256
rect 548614 603064 548670 603120
rect 553306 603064 553362 603120
rect 441526 602928 441582 602984
rect 560298 603492 560354 603528
rect 560298 603472 560300 603492
rect 560300 603472 560352 603492
rect 560352 603472 560354 603492
rect 565174 603336 565230 603392
rect 572718 603336 572774 603392
rect 572626 603200 572682 603256
rect 580170 592456 580226 592512
rect 580170 580760 580226 580816
rect 259182 553444 259238 553480
rect 259182 553424 259184 553444
rect 259184 553424 259236 553444
rect 259236 553424 259238 553444
rect 263782 553444 263838 553480
rect 263782 553424 263784 553444
rect 263784 553424 263836 553444
rect 263836 553424 263838 553444
rect 378506 553444 378562 553480
rect 378506 553424 378508 553444
rect 378508 553424 378560 553444
rect 378560 553424 378562 553444
rect 382922 553444 382978 553480
rect 382922 553424 382924 553444
rect 382924 553424 382976 553444
rect 382976 553424 382978 553444
rect 139398 549888 139454 549944
rect 266450 549888 266506 549944
rect 270406 549344 270462 549400
rect 389178 549888 389234 549944
rect 187698 546508 187754 546544
rect 187698 546488 187700 546508
rect 187700 546488 187752 546508
rect 187752 546488 187754 546508
rect 139398 489504 139454 489560
rect 187698 545148 187754 545184
rect 187698 545128 187700 545148
rect 187700 545128 187752 545148
rect 187752 545128 187754 545148
rect 187698 543788 187754 543824
rect 187698 543768 187700 543788
rect 187700 543768 187752 543788
rect 187752 543768 187754 543788
rect 187698 542544 187754 542600
rect 187790 540368 187846 540424
rect 187698 539824 187754 539880
rect 188342 537512 188398 537568
rect 162950 442448 163006 442504
rect 165250 442312 165306 442368
rect 167458 442176 167514 442232
rect 299478 531256 299534 531312
rect 299662 531292 299664 531312
rect 299664 531292 299716 531312
rect 299716 531292 299718 531312
rect 299662 531256 299718 531292
rect 299478 511944 299534 512000
rect 299662 511944 299718 512000
rect 269118 484472 269174 484528
rect 299478 482976 299534 483032
rect 299754 482976 299810 483032
rect 188986 480256 189042 480312
rect 188894 477944 188950 478000
rect 193862 458088 193918 458144
rect 197358 457952 197414 458008
rect 198738 457952 198794 458008
rect 200210 458088 200266 458144
rect 195978 457544 196034 457600
rect 207662 457952 207718 458008
rect 208214 457952 208270 458008
rect 201498 457700 201554 457736
rect 201498 457680 201500 457700
rect 201500 457680 201552 457700
rect 201552 457680 201554 457700
rect 206282 457272 206338 457328
rect 206834 457272 206890 457328
rect 202142 457136 202198 457192
rect 202786 457136 202842 457192
rect 204902 457000 204958 457056
rect 205454 457000 205510 457056
rect 203522 456864 203578 456920
rect 204166 456864 204222 456920
rect 205546 456864 205602 456920
rect 206926 457136 206982 457192
rect 209686 457700 209742 457736
rect 209686 457680 209688 457700
rect 209688 457680 209740 457700
rect 209740 457680 209742 457700
rect 209042 457428 209098 457464
rect 209042 457408 209044 457428
rect 209044 457408 209096 457428
rect 209096 457408 209098 457428
rect 208306 456864 208362 456920
rect 210514 458088 210570 458144
rect 212446 458088 212502 458144
rect 213090 458088 213146 458144
rect 214010 458088 214066 458144
rect 215298 458124 215300 458144
rect 215300 458124 215352 458144
rect 215352 458124 215354 458144
rect 215298 458088 215354 458124
rect 216678 458088 216734 458144
rect 209686 456864 209742 456920
rect 210974 457136 211030 457192
rect 211066 456864 211122 456920
rect 212446 456864 212502 456920
rect 213826 456864 213882 456920
rect 215206 457156 215262 457192
rect 215206 457136 215208 457156
rect 215208 457136 215260 457156
rect 215260 457136 215262 457156
rect 217598 458088 217654 458144
rect 218886 458088 218942 458144
rect 216586 457408 216642 457464
rect 220174 458088 220230 458144
rect 221370 458088 221426 458144
rect 222566 458088 222622 458144
rect 217966 457136 218022 457192
rect 220726 457136 220782 457192
rect 217874 456864 217930 456920
rect 219346 456864 219402 456920
rect 223670 458108 223726 458144
rect 223670 458088 223672 458108
rect 223672 458088 223724 458108
rect 223724 458088 223726 458108
rect 224314 458088 224370 458144
rect 225878 458088 225934 458144
rect 222106 456864 222162 456920
rect 223486 456864 223542 456920
rect 226246 457000 226302 457056
rect 224866 456864 224922 456920
rect 226154 456864 226210 456920
rect 227166 458088 227222 458144
rect 228362 458088 228418 458144
rect 229558 458088 229614 458144
rect 231858 458108 231914 458144
rect 231858 458088 231860 458108
rect 231860 458088 231912 458108
rect 231912 458088 231914 458108
rect 233238 458088 233294 458144
rect 234618 457972 234674 458008
rect 234618 457952 234620 457972
rect 234620 457952 234672 457972
rect 234672 457952 234674 457972
rect 231858 457836 231914 457872
rect 231858 457816 231860 457836
rect 231860 457816 231912 457836
rect 231912 457816 231914 457836
rect 235998 457816 236054 457872
rect 237378 457700 237434 457736
rect 237378 457680 237380 457700
rect 237380 457680 237432 457700
rect 237432 457680 237434 457700
rect 238758 457680 238814 457736
rect 230478 457564 230534 457600
rect 230478 457544 230480 457564
rect 230480 457544 230532 457564
rect 230532 457544 230534 457564
rect 233054 457000 233110 457056
rect 227626 456864 227682 456920
rect 229006 456864 229062 456920
rect 230386 456864 230442 456920
rect 231766 456864 231822 456920
rect 233146 456864 233202 456920
rect 234526 456864 234582 456920
rect 235906 456864 235962 456920
rect 237286 456864 237342 456920
rect 238666 456864 238722 456920
rect 240046 456864 240102 456920
rect 233146 442448 233202 442504
rect 234526 442312 234582 442368
rect 237286 442176 237342 442232
rect 240046 441632 240102 441688
rect 248694 441632 248750 441688
rect 287518 442448 287574 442504
rect 289726 442312 289782 442368
rect 294326 442176 294382 442232
rect 507858 553444 507914 553480
rect 507858 553424 507860 553444
rect 507860 553424 507912 553444
rect 507912 553424 507914 553444
rect 513378 553424 513434 553480
rect 580170 557232 580226 557288
rect 518898 550704 518954 550760
rect 305826 546488 305882 546544
rect 302790 436736 302846 436792
rect 302790 434560 302846 434616
rect 302790 432384 302846 432440
rect 302790 430208 302846 430264
rect 302790 427896 302846 427952
rect 302790 425720 302846 425776
rect 302790 423580 302792 423600
rect 302792 423580 302844 423600
rect 302844 423580 302846 423600
rect 302790 423544 302846 423580
rect 302790 421368 302846 421424
rect 302790 419192 302846 419248
rect 302790 416880 302846 416936
rect 302790 414704 302846 414760
rect 302790 412564 302792 412584
rect 302792 412564 302844 412584
rect 302844 412564 302846 412584
rect 302790 412528 302846 412564
rect 302790 410352 302846 410408
rect 302790 408176 302846 408232
rect 302790 405864 302846 405920
rect 302698 403688 302754 403744
rect 302790 401548 302792 401568
rect 302792 401548 302844 401568
rect 302844 401548 302846 401568
rect 302790 401512 302846 401548
rect 302790 399336 302846 399392
rect 302790 397160 302846 397216
rect 302514 394848 302570 394904
rect 302698 392672 302754 392728
rect 302790 390516 302846 390552
rect 302790 390496 302792 390516
rect 302792 390496 302844 390516
rect 302844 390496 302846 390516
rect 302790 388320 302846 388376
rect 302514 386144 302570 386200
rect 302514 383832 302570 383888
rect 302790 381656 302846 381712
rect 302606 379480 302662 379536
rect 302790 377304 302846 377360
rect 302790 375128 302846 375184
rect 302790 372952 302846 373008
rect 302330 370640 302386 370696
rect 302606 368464 302662 368520
rect 302790 366288 302846 366344
rect 302514 364112 302570 364168
rect 302422 361936 302478 361992
rect 302330 359624 302386 359680
rect 302514 357448 302570 357504
rect 302790 355272 302846 355328
rect 302790 353096 302846 353152
rect 302422 350920 302478 350976
rect 302698 348608 302754 348664
rect 302514 346432 302570 346488
rect 302790 344256 302846 344312
rect 302790 342080 302846 342136
rect 302422 339904 302478 339960
rect 302698 337592 302754 337648
rect 302514 335416 302570 335472
rect 302790 333240 302846 333296
rect 302514 331100 302516 331120
rect 302516 331100 302568 331120
rect 302568 331100 302570 331120
rect 302514 331064 302570 331100
rect 302330 328888 302386 328944
rect 302514 326576 302570 326632
rect 302330 324436 302332 324456
rect 302332 324436 302384 324456
rect 302384 324436 302386 324456
rect 302330 324400 302386 324436
rect 302330 322224 302386 322280
rect 302330 320084 302332 320104
rect 302332 320084 302384 320104
rect 302384 320084 302386 320104
rect 302330 320048 302386 320084
rect 302698 317872 302754 317928
rect 302790 315696 302846 315752
rect 302790 313384 302846 313440
rect 302698 311208 302754 311264
rect 302790 309068 302792 309088
rect 302792 309068 302844 309088
rect 302844 309068 302846 309088
rect 302790 309032 302846 309068
rect 302790 306856 302846 306912
rect 302790 304680 302846 304736
rect 302790 302368 302846 302424
rect 302698 300192 302754 300248
rect 302790 298052 302792 298072
rect 302792 298052 302844 298072
rect 302844 298052 302846 298072
rect 302790 298016 302846 298052
rect 302606 295876 302608 295896
rect 302608 295876 302660 295896
rect 302660 295876 302662 295896
rect 302606 295840 302662 295876
rect 302790 293664 302846 293720
rect 302514 291352 302570 291408
rect 302698 289176 302754 289232
rect 302790 287020 302846 287056
rect 302790 287000 302792 287020
rect 302792 287000 302844 287020
rect 302844 287000 302846 287020
rect 302698 284824 302754 284880
rect 302514 282648 302570 282704
rect 302514 280336 302570 280392
rect 302330 278160 302386 278216
rect 302606 275984 302662 276040
rect 302790 273808 302846 273864
rect 302514 271632 302570 271688
rect 302514 269320 302570 269376
rect 302330 267144 302386 267200
rect 302606 264968 302662 265024
rect 302790 262792 302846 262848
rect 302514 260616 302570 260672
rect 302422 258440 302478 258496
rect 302330 256128 302386 256184
rect 302514 253952 302570 254008
rect 302790 251776 302846 251832
rect 302790 249600 302846 249656
rect 302422 247424 302478 247480
rect 302698 245112 302754 245168
rect 302514 242936 302570 242992
rect 302790 240760 302846 240816
rect 302790 238584 302846 238640
rect 302422 236408 302478 236464
rect 302698 234096 302754 234152
rect 302514 231920 302570 231976
rect 302790 229744 302846 229800
rect 302790 227568 302846 227624
rect 302790 225392 302846 225448
rect 302698 223080 302754 223136
rect 302790 220904 302846 220960
rect 302790 218728 302846 218784
rect 302790 216588 302792 216608
rect 302792 216588 302844 216608
rect 302844 216588 302846 216608
rect 302790 216552 302846 216588
rect 302790 214376 302846 214432
rect 302606 212064 302662 212120
rect 302790 209888 302846 209944
rect 302790 207712 302846 207768
rect 302790 205572 302792 205592
rect 302792 205572 302844 205592
rect 302844 205572 302846 205592
rect 302790 205536 302846 205572
rect 302238 203360 302294 203416
rect 302974 438912 303030 438968
rect 305734 543768 305790 543824
rect 305642 539552 305698 539608
rect 307666 545148 307722 545184
rect 307666 545128 307668 545148
rect 307668 545128 307720 545148
rect 307720 545128 307722 545148
rect 307206 542428 307262 542464
rect 307206 542408 307208 542428
rect 307208 542408 307260 542428
rect 307260 542408 307262 542428
rect 307298 540368 307354 540424
rect 307666 539824 307722 539880
rect 307298 539552 307354 539608
rect 307022 537512 307078 537568
rect 305918 480256 305974 480312
rect 307114 478080 307170 478136
rect 351826 459584 351882 459640
rect 327906 459448 327962 459504
rect 313738 458088 313794 458144
rect 321558 458088 321614 458144
rect 322938 458088 322994 458144
rect 325698 458088 325754 458144
rect 327078 458088 327134 458144
rect 317418 457816 317474 457872
rect 320270 457000 320326 457056
rect 316038 456864 316094 456920
rect 318798 456864 318854 456920
rect 320178 456864 320234 456920
rect 322202 457952 322258 458008
rect 323582 457952 323638 458008
rect 324962 457816 325018 457872
rect 324318 457136 324374 457192
rect 326342 457816 326398 457872
rect 329102 458108 329158 458144
rect 329102 458088 329104 458108
rect 329104 458088 329156 458108
rect 329156 458088 329158 458108
rect 329930 458088 329986 458144
rect 331862 458088 331918 458144
rect 333150 458088 333206 458144
rect 334070 458088 334126 458144
rect 335358 458124 335360 458144
rect 335360 458124 335412 458144
rect 335412 458124 335414 458144
rect 335358 458088 335414 458124
rect 328458 457156 328514 457192
rect 328458 457136 328460 457156
rect 328460 457136 328512 457156
rect 328512 457136 328514 457156
rect 327722 454008 327778 454064
rect 327906 454008 327962 454064
rect 327814 366968 327870 367024
rect 328090 366968 328146 367024
rect 329286 457952 329342 458008
rect 329838 457292 329894 457328
rect 329838 457272 329840 457292
rect 329840 457272 329892 457292
rect 329892 457272 329894 457292
rect 330482 457816 330538 457872
rect 331218 457680 331274 457736
rect 335358 457136 335414 457192
rect 332598 456864 332654 456920
rect 333978 456864 334034 456920
rect 336554 458088 336610 458144
rect 338026 458108 338082 458144
rect 338026 458088 338028 458108
rect 338028 458088 338080 458108
rect 338080 458088 338082 458108
rect 339038 458088 339094 458144
rect 339866 458088 339922 458144
rect 341246 458088 341302 458144
rect 342258 458088 342314 458144
rect 343638 458088 343694 458144
rect 344742 458124 344744 458144
rect 344744 458124 344796 458144
rect 344796 458124 344798 458144
rect 336830 457000 336886 457056
rect 336738 456864 336794 456920
rect 338118 456864 338174 456920
rect 339498 456864 339554 456920
rect 340878 457136 340934 457192
rect 342534 457952 342590 458008
rect 344742 458088 344798 458124
rect 345018 458088 345074 458144
rect 346398 458088 346454 458144
rect 347778 458088 347834 458144
rect 349158 458088 349214 458144
rect 344374 457952 344430 458008
rect 343730 457680 343786 457736
rect 345938 457972 345994 458008
rect 345938 457952 345940 457972
rect 345940 457952 345992 457972
rect 345992 457952 345994 457972
rect 346858 457952 346914 458008
rect 348238 457952 348294 458008
rect 358818 459448 358874 459504
rect 351918 458108 351974 458144
rect 353298 458124 353300 458144
rect 353300 458124 353352 458144
rect 353352 458124 353354 458144
rect 351918 458088 351920 458108
rect 351920 458088 351972 458108
rect 351972 458088 351974 458108
rect 353298 458088 353354 458124
rect 349250 457952 349306 458008
rect 350538 457952 350594 458008
rect 350538 456864 350594 456920
rect 352010 457000 352066 457056
rect 351918 456864 351974 456920
rect 353298 457136 353354 457192
rect 356058 457952 356114 458008
rect 355046 457816 355102 457872
rect 357438 457700 357494 457736
rect 357438 457680 357440 457700
rect 357440 457680 357492 457700
rect 357492 457680 357494 457700
rect 354678 456864 354734 456920
rect 356058 456864 356114 456920
rect 357438 456864 357494 456920
rect 358818 456864 358874 456920
rect 389178 489504 389234 489560
rect 389178 480936 389234 480992
rect 516414 549888 516470 549944
rect 437478 546508 437534 546544
rect 437478 546488 437480 546508
rect 437480 546488 437532 546508
rect 437532 546488 437534 546508
rect 437478 545148 437534 545184
rect 437478 545128 437480 545148
rect 437480 545128 437532 545148
rect 437532 545128 437534 545148
rect 429566 543768 429622 543824
rect 437478 543788 437534 543824
rect 437478 543768 437480 543788
rect 437480 543768 437532 543788
rect 437532 543768 437534 543788
rect 429382 543632 429438 543688
rect 437478 542428 437534 542464
rect 437478 542408 437480 542428
rect 437480 542408 437532 542428
rect 437532 542408 437534 542428
rect 429198 540912 429254 540968
rect 429382 540912 429438 540968
rect 437570 540368 437626 540424
rect 437478 539824 437534 539880
rect 437478 537512 437534 537568
rect 429382 521600 429438 521656
rect 429566 521600 429622 521656
rect 580262 545536 580318 545592
rect 559102 521600 559158 521656
rect 559286 521600 559342 521656
rect 559194 492768 559250 492824
rect 559102 492652 559158 492688
rect 559102 492632 559104 492652
rect 559104 492632 559156 492652
rect 559156 492632 559158 492652
rect 518898 489504 518954 489560
rect 437478 480276 437534 480312
rect 437478 480256 437480 480276
rect 437480 480256 437532 480276
rect 437532 480256 437534 480276
rect 438122 477944 438178 478000
rect 429474 463664 429530 463720
rect 429658 463664 429714 463720
rect 483018 459448 483074 459504
rect 461766 458088 461822 458144
rect 463054 458088 463110 458144
rect 464986 458088 465042 458144
rect 465170 458088 465226 458144
rect 468758 458088 468814 458144
rect 469954 458088 470010 458144
rect 471794 458088 471850 458144
rect 472254 458088 472310 458144
rect 473450 458088 473506 458144
rect 474830 458088 474886 458144
rect 475474 458088 475530 458144
rect 476946 458088 477002 458144
rect 478326 458088 478382 458144
rect 479430 458088 479486 458144
rect 483018 458108 483074 458144
rect 483018 458088 483020 458108
rect 483020 458088 483072 458108
rect 483072 458088 483074 458108
rect 442998 457952 443054 458008
rect 460202 457952 460258 458008
rect 458178 457816 458234 457872
rect 452658 457408 452714 457464
rect 450542 457136 450598 457192
rect 446402 457000 446458 457056
rect 445758 456864 445814 456920
rect 447782 456864 447838 456920
rect 449162 456864 449218 456920
rect 456798 457564 456854 457600
rect 456798 457544 456800 457564
rect 456800 457544 456852 457564
rect 456852 457544 456854 457564
rect 459558 457544 459614 457600
rect 454038 457428 454094 457464
rect 454038 457408 454040 457428
rect 454040 457408 454092 457428
rect 454092 457408 454094 457428
rect 454682 457136 454738 457192
rect 458822 457136 458878 457192
rect 459374 457136 459430 457192
rect 452750 456864 452806 456920
rect 453302 456864 453358 456920
rect 453486 456864 453542 456920
rect 456062 457000 456118 457056
rect 456706 457000 456762 457056
rect 455418 456884 455474 456920
rect 455418 456864 455420 456884
rect 455420 456864 455472 456884
rect 455472 456864 455474 456884
rect 457442 456864 457498 456920
rect 458086 456864 458142 456920
rect 460386 457700 460442 457736
rect 460386 457680 460388 457700
rect 460388 457680 460440 457700
rect 460440 457680 460442 457700
rect 468022 457952 468078 458008
rect 466642 457816 466698 457872
rect 461030 457136 461086 457192
rect 460938 456864 460994 456920
rect 462318 456864 462374 456920
rect 463698 456864 463754 456920
rect 465078 456864 465134 456920
rect 466458 456864 466514 456920
rect 467930 457136 467986 457192
rect 467838 456864 467894 456920
rect 469218 456864 469274 456920
rect 470598 456864 470654 456920
rect 471978 457136 472034 457192
rect 473358 456864 473414 456920
rect 474738 456864 474794 456920
rect 478878 457816 478934 457872
rect 476118 457272 476174 457328
rect 476210 457136 476266 457192
rect 477498 457292 477554 457328
rect 477498 457272 477500 457292
rect 477500 457272 477552 457292
rect 477552 457272 477554 457292
rect 480442 457972 480498 458008
rect 480442 457952 480444 457972
rect 480444 457952 480496 457972
rect 480496 457952 480498 457972
rect 480534 457816 480590 457872
rect 481638 457680 481694 457736
rect 483018 457408 483074 457464
rect 481638 457136 481694 457192
rect 483202 458088 483258 458144
rect 484398 458124 484400 458144
rect 484400 458124 484452 458144
rect 484452 458124 484454 458144
rect 484398 458088 484454 458124
rect 487158 457952 487214 458008
rect 484398 457836 484454 457872
rect 484398 457816 484400 457836
rect 484400 457816 484452 457836
rect 484452 457816 484454 457836
rect 485778 457680 485834 457736
rect 488538 457700 488594 457736
rect 488538 457680 488540 457700
rect 488540 457680 488592 457700
rect 488592 457680 488594 457700
rect 487158 457544 487214 457600
rect 485778 457408 485834 457464
rect 488538 457428 488594 457464
rect 488538 457408 488540 457428
rect 488540 457408 488592 457428
rect 488592 457408 488594 457428
rect 580170 451696 580226 451752
rect 580078 439864 580134 439920
rect 559102 439592 559158 439648
rect 580354 533840 580410 533896
rect 580446 510312 580502 510368
rect 580538 498616 580594 498672
rect 580446 439456 580502 439512
rect 580722 486784 580778 486840
rect 580814 463392 580870 463448
rect 580446 416472 580502 416528
rect 580354 404776 580410 404832
rect 580630 392944 580686 393000
rect 580262 369552 580318 369608
rect 580170 252184 580226 252240
rect 580078 228792 580134 228848
rect 579986 216960 580042 217016
rect 302882 201184 302938 201240
rect 580170 205264 580226 205320
rect 580354 357856 580410 357912
rect 580262 200640 580318 200696
rect 580446 346024 580502 346080
rect 80242 5208 80298 5264
rect 89626 110780 89628 110800
rect 89628 110780 89680 110800
rect 89680 110780 89682 110800
rect 89626 110744 89682 110780
rect 89626 87252 89628 87272
rect 89628 87252 89680 87272
rect 89680 87252 89682 87272
rect 89626 87216 89682 87252
rect 89626 76236 89628 76256
rect 89628 76236 89680 76256
rect 89680 76236 89682 76256
rect 89626 76200 89682 76236
rect 88890 63860 88892 63880
rect 88892 63860 88944 63880
rect 88944 63860 88946 63880
rect 88890 63824 88946 63860
rect 88890 40332 88892 40352
rect 88892 40332 88944 40352
rect 88944 40332 88946 40352
rect 88890 40296 88946 40332
rect 89626 29316 89628 29336
rect 89628 29316 89680 29336
rect 89680 29316 89682 29336
rect 89626 29280 89682 29316
rect 92202 193160 92258 193216
rect 92386 193160 92442 193216
rect 92202 173848 92258 173904
rect 92386 173848 92442 173904
rect 92202 164192 92258 164248
rect 92386 164192 92442 164248
rect 92202 144880 92258 144936
rect 92386 144880 92442 144936
rect 92110 125568 92166 125624
rect 92386 125568 92442 125624
rect 87326 5072 87382 5128
rect 89718 3712 89774 3768
rect 96526 110780 96528 110800
rect 96528 110780 96580 110800
rect 96580 110780 96582 110800
rect 96526 110744 96582 110780
rect 96526 87252 96528 87272
rect 96528 87252 96580 87272
rect 96580 87252 96582 87272
rect 96526 87216 96582 87252
rect 96526 76236 96528 76256
rect 96528 76236 96580 76256
rect 96580 76236 96582 76256
rect 96526 76200 96582 76236
rect 96526 63860 96528 63880
rect 96528 63860 96580 63880
rect 96580 63860 96582 63880
rect 96526 63824 96582 63860
rect 96526 40332 96528 40352
rect 96528 40332 96580 40352
rect 96580 40332 96582 40352
rect 96526 40296 96582 40332
rect 96526 29316 96528 29336
rect 96528 29316 96580 29336
rect 96580 29316 96582 29336
rect 96526 29280 96582 29316
rect 94502 4936 94558 4992
rect 96894 3576 96950 3632
rect 105174 4800 105230 4856
rect 106278 3984 106334 4040
rect 111154 3440 111210 3496
rect 115846 198056 115902 198112
rect 114650 3848 114706 3904
rect 115662 3984 115718 4040
rect 117226 197920 117282 197976
rect 116030 110508 116032 110528
rect 116032 110508 116084 110528
rect 116084 110508 116086 110528
rect 116030 110472 116086 110508
rect 116030 86980 116032 87000
rect 116032 86980 116084 87000
rect 116084 86980 116086 87000
rect 116030 86944 116086 86980
rect 116030 75964 116032 75984
rect 116032 75964 116084 75984
rect 116084 75964 116086 75984
rect 116030 75928 116086 75964
rect 116030 63588 116032 63608
rect 116032 63588 116084 63608
rect 116084 63588 116086 63608
rect 116030 63552 116086 63588
rect 116030 40060 116032 40080
rect 116032 40060 116084 40080
rect 116084 40060 116086 40080
rect 116030 40024 116086 40060
rect 116030 29044 116032 29064
rect 116032 29044 116084 29064
rect 116084 29044 116086 29064
rect 116030 29008 116086 29044
rect 118790 110744 118846 110800
rect 118790 76200 118846 76256
rect 118790 63824 118846 63880
rect 118790 40296 118846 40352
rect 117318 3848 117374 3904
rect 120814 87216 120870 87272
rect 120814 29280 120870 29336
rect 125414 3304 125470 3360
rect 128174 87216 128230 87272
rect 128358 87216 128414 87272
rect 128174 29280 128230 29336
rect 128358 29280 128414 29336
rect 135166 111016 135222 111072
rect 135166 110608 135222 110664
rect 135166 76472 135222 76528
rect 135166 76064 135222 76120
rect 135166 64096 135222 64152
rect 135166 63688 135222 63744
rect 135166 40568 135222 40624
rect 135166 40160 135222 40216
rect 140042 110880 140098 110936
rect 140042 110472 140098 110528
rect 140042 76336 140098 76392
rect 140042 75928 140098 75984
rect 140042 63960 140098 64016
rect 140042 63552 140098 63608
rect 140042 40432 140098 40488
rect 140042 40024 140098 40080
rect 143446 87352 143502 87408
rect 143446 86944 143502 87000
rect 143446 29416 143502 29472
rect 143446 29008 143502 29064
rect 147586 110644 147588 110664
rect 147588 110644 147640 110664
rect 147640 110644 147642 110664
rect 147586 110608 147642 110644
rect 145562 86944 145618 87000
rect 147586 76100 147588 76120
rect 147588 76100 147640 76120
rect 147640 76100 147642 76120
rect 147586 76064 147642 76100
rect 147586 63724 147588 63744
rect 147588 63724 147640 63744
rect 147640 63724 147642 63744
rect 147586 63688 147642 63724
rect 147586 40196 147588 40216
rect 147588 40196 147640 40216
rect 147640 40196 147642 40216
rect 147586 40160 147642 40196
rect 145010 29044 145012 29064
rect 145012 29044 145064 29064
rect 145064 29044 145066 29064
rect 145010 29008 145066 29044
rect 154486 110744 154542 110800
rect 154486 87216 154542 87272
rect 154486 76200 154542 76256
rect 154486 63824 154542 63880
rect 154486 40296 154542 40352
rect 154486 29280 154542 29336
rect 202878 5208 202934 5264
rect 215298 5072 215354 5128
rect 227718 4936 227774 4992
rect 219438 3712 219494 3768
rect 247038 4800 247094 4856
rect 231858 3576 231914 3632
rect 264886 198056 264942 198112
rect 269118 197920 269174 197976
rect 258078 3440 258134 3496
rect 580538 322632 580594 322688
rect 580630 310800 580686 310856
rect 580722 299104 580778 299160
rect 580814 275712 580870 275768
rect 580906 263880 580962 263936
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 17584 579858 17640
rect 282918 3304 282974 3360
<< metal3 >>
rect 57462 700708 57468 700772
rect 57532 700770 57538 700772
rect 478505 700770 478571 700773
rect 57532 700768 478571 700770
rect 57532 700712 478510 700768
rect 478566 700712 478571 700768
rect 57532 700710 478571 700712
rect 57532 700708 57538 700710
rect 478505 700707 478571 700710
rect 57646 700572 57652 700636
rect 57716 700634 57722 700636
rect 494789 700634 494855 700637
rect 57716 700632 494855 700634
rect 57716 700576 494794 700632
rect 494850 700576 494855 700632
rect 57716 700574 494855 700576
rect 57716 700572 57722 700574
rect 494789 700571 494855 700574
rect 59118 700436 59124 700500
rect 59188 700498 59194 700500
rect 527173 700498 527239 700501
rect 59188 700496 527239 700498
rect 59188 700440 527178 700496
rect 527234 700440 527239 700496
rect 59188 700438 527239 700440
rect 59188 700436 59194 700438
rect 527173 700435 527239 700438
rect 57830 700300 57836 700364
rect 57900 700362 57906 700364
rect 543457 700362 543523 700365
rect 57900 700360 543523 700362
rect 57900 700304 543462 700360
rect 543518 700304 543523 700360
rect 57900 700302 543523 700304
rect 57900 700300 57906 700302
rect 543457 700299 543523 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 4797 682274 4863 682277
rect -960 682272 4863 682274
rect -960 682216 4802 682272
rect 4858 682216 4863 682272
rect -960 682214 4863 682216
rect -960 682124 480 682214
rect 4797 682211 4863 682214
rect 583520 674658 584960 674748
rect 583342 674598 584960 674658
rect 550582 673916 550588 673980
rect 550652 673978 550658 673980
rect 553301 673978 553367 673981
rect 550652 673976 553367 673978
rect 550652 673920 553306 673976
rect 553362 673920 553367 673976
rect 550652 673918 553367 673920
rect 550652 673916 550658 673918
rect 553301 673915 553367 673918
rect 553485 673978 553551 673981
rect 560293 673978 560359 673981
rect 553485 673976 560359 673978
rect 553485 673920 553490 673976
rect 553546 673920 560298 673976
rect 560354 673920 560359 673976
rect 553485 673918 560359 673920
rect 553485 673915 553551 673918
rect 560293 673915 560359 673918
rect 57278 673780 57284 673844
rect 57348 673842 57354 673844
rect 289813 673842 289879 673845
rect 57348 673782 64890 673842
rect 57348 673780 57354 673782
rect 64830 673706 64890 673782
rect 74582 673782 84210 673842
rect 64830 673646 74458 673706
rect 74398 673570 74458 673646
rect 74582 673570 74642 673782
rect 84150 673706 84210 673782
rect 93902 673782 103530 673842
rect 84150 673646 93778 673706
rect 74398 673510 74642 673570
rect 93718 673570 93778 673646
rect 93902 673570 93962 673782
rect 103470 673706 103530 673782
rect 113222 673782 122850 673842
rect 103470 673646 113098 673706
rect 93718 673510 93962 673570
rect 113038 673570 113098 673646
rect 113222 673570 113282 673782
rect 122790 673706 122850 673782
rect 132542 673782 142170 673842
rect 122790 673646 132418 673706
rect 113038 673510 113282 673570
rect 132358 673570 132418 673646
rect 132542 673570 132602 673782
rect 142110 673706 142170 673782
rect 151862 673782 161490 673842
rect 142110 673646 151738 673706
rect 132358 673510 132602 673570
rect 151678 673570 151738 673646
rect 151862 673570 151922 673782
rect 161430 673706 161490 673782
rect 171182 673782 180810 673842
rect 161430 673646 171058 673706
rect 151678 673510 151922 673570
rect 170998 673570 171058 673646
rect 171182 673570 171242 673782
rect 180750 673706 180810 673782
rect 190502 673782 200130 673842
rect 180750 673646 190378 673706
rect 170998 673510 171242 673570
rect 190318 673570 190378 673646
rect 190502 673570 190562 673782
rect 200070 673706 200130 673782
rect 209822 673782 219450 673842
rect 200070 673646 209698 673706
rect 190318 673510 190562 673570
rect 209638 673570 209698 673646
rect 209822 673570 209882 673782
rect 219390 673706 219450 673782
rect 229142 673782 238770 673842
rect 219390 673646 229018 673706
rect 209638 673510 209882 673570
rect 228958 673570 229018 673646
rect 229142 673570 229202 673782
rect 238710 673706 238770 673782
rect 248462 673782 258090 673842
rect 238710 673646 248338 673706
rect 228958 673510 229202 673570
rect 248278 673570 248338 673646
rect 248462 673570 248522 673782
rect 258030 673706 258090 673782
rect 267782 673782 277410 673842
rect 258030 673646 267658 673706
rect 248278 673510 248522 673570
rect 267598 673570 267658 673646
rect 267782 673570 267842 673782
rect 277350 673706 277410 673782
rect 287102 673840 289879 673842
rect 287102 673784 289818 673840
rect 289874 673784 289879 673840
rect 287102 673782 289879 673784
rect 277350 673646 286978 673706
rect 267598 673510 267842 673570
rect 286918 673570 286978 673646
rect 287102 673570 287162 673782
rect 289813 673779 289879 673782
rect 299422 673780 299428 673844
rect 299492 673842 299498 673844
rect 540973 673842 541039 673845
rect 299492 673782 316050 673842
rect 299492 673780 299498 673782
rect 315990 673706 316050 673782
rect 325742 673782 335370 673842
rect 315990 673646 325618 673706
rect 286918 673510 287162 673570
rect 292665 673570 292731 673573
rect 299422 673570 299428 673572
rect 292665 673568 299428 673570
rect 292665 673512 292670 673568
rect 292726 673512 299428 673568
rect 292665 673510 299428 673512
rect 292665 673507 292731 673510
rect 299422 673508 299428 673510
rect 299492 673508 299498 673572
rect 325558 673570 325618 673646
rect 325742 673570 325802 673782
rect 335310 673706 335370 673782
rect 345062 673782 354690 673842
rect 335310 673646 344938 673706
rect 325558 673510 325802 673570
rect 344878 673570 344938 673646
rect 345062 673570 345122 673782
rect 354630 673706 354690 673782
rect 364382 673782 374010 673842
rect 354630 673646 364258 673706
rect 344878 673510 345122 673570
rect 364198 673570 364258 673646
rect 364382 673570 364442 673782
rect 373950 673706 374010 673782
rect 383702 673782 393330 673842
rect 373950 673646 383578 673706
rect 364198 673510 364442 673570
rect 383518 673570 383578 673646
rect 383702 673570 383762 673782
rect 393270 673706 393330 673782
rect 403022 673782 412650 673842
rect 393270 673646 402898 673706
rect 383518 673510 383762 673570
rect 402838 673570 402898 673646
rect 403022 673570 403082 673782
rect 412590 673706 412650 673782
rect 431910 673782 441538 673842
rect 412590 673646 422218 673706
rect 402838 673510 403082 673570
rect 422158 673570 422218 673646
rect 431910 673570 431970 673782
rect 422158 673510 431970 673570
rect 441478 673570 441538 673782
rect 441662 673782 451290 673842
rect 441662 673570 441722 673782
rect 451230 673706 451290 673782
rect 460982 673782 470610 673842
rect 451230 673646 460858 673706
rect 441478 673510 441722 673570
rect 460798 673570 460858 673646
rect 460982 673570 461042 673782
rect 470550 673706 470610 673782
rect 480302 673782 489930 673842
rect 470550 673646 480178 673706
rect 460798 673510 461042 673570
rect 480118 673570 480178 673646
rect 480302 673570 480362 673782
rect 489870 673706 489930 673782
rect 499622 673782 509250 673842
rect 489870 673646 499498 673706
rect 480118 673510 480362 673570
rect 499438 673570 499498 673646
rect 499622 673570 499682 673782
rect 509190 673706 509250 673782
rect 518942 673782 528570 673842
rect 509190 673646 518818 673706
rect 499438 673510 499682 673570
rect 518758 673570 518818 673646
rect 518942 673570 519002 673782
rect 528510 673706 528570 673782
rect 538262 673840 541039 673842
rect 538262 673784 540978 673840
rect 541034 673784 541039 673840
rect 538262 673782 541039 673784
rect 528510 673646 538138 673706
rect 518758 673510 519002 673570
rect 538078 673570 538138 673646
rect 538262 673570 538322 673782
rect 540973 673779 541039 673782
rect 565169 673842 565235 673845
rect 572713 673842 572779 673845
rect 565169 673840 569970 673842
rect 565169 673784 565174 673840
rect 565230 673784 569970 673840
rect 565169 673782 569970 673784
rect 565169 673779 565235 673782
rect 569910 673706 569970 673782
rect 572713 673840 576962 673842
rect 572713 673784 572718 673840
rect 572774 673784 576962 673840
rect 572713 673782 576962 673784
rect 572713 673779 572779 673782
rect 572621 673706 572687 673709
rect 569910 673704 572687 673706
rect 569910 673648 572626 673704
rect 572682 673648 572687 673704
rect 569910 673646 572687 673648
rect 576902 673706 576962 673782
rect 583342 673706 583402 674598
rect 583520 674508 584960 674598
rect 576902 673646 583402 673706
rect 572621 673643 572687 673646
rect 538078 673510 538322 673570
rect 548609 673570 548675 673573
rect 550582 673570 550588 673572
rect 548609 673568 550588 673570
rect 548609 673512 548614 673568
rect 548670 673512 550588 673568
rect 548609 673510 550588 673512
rect 548609 673507 548675 673510
rect 550582 673508 550588 673510
rect 550652 673508 550658 673572
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 583520 651130 584960 651220
rect 583342 651070 584960 651130
rect 550582 650388 550588 650452
rect 550652 650450 550658 650452
rect 553301 650450 553367 650453
rect 550652 650448 553367 650450
rect 550652 650392 553306 650448
rect 553362 650392 553367 650448
rect 550652 650390 553367 650392
rect 550652 650388 550658 650390
rect 553301 650387 553367 650390
rect 553485 650450 553551 650453
rect 560293 650450 560359 650453
rect 553485 650448 560359 650450
rect 553485 650392 553490 650448
rect 553546 650392 560298 650448
rect 560354 650392 560359 650448
rect 553485 650390 560359 650392
rect 553485 650387 553551 650390
rect 560293 650387 560359 650390
rect 58198 650252 58204 650316
rect 58268 650314 58274 650316
rect 58268 650254 64890 650314
rect 58268 650252 58274 650254
rect 64830 650178 64890 650254
rect 74582 650254 84210 650314
rect 64830 650118 74458 650178
rect 74398 650042 74458 650118
rect 74582 650042 74642 650254
rect 84150 650178 84210 650254
rect 93902 650254 103530 650314
rect 84150 650118 93778 650178
rect 74398 649982 74642 650042
rect 93718 650042 93778 650118
rect 93902 650042 93962 650254
rect 103470 650178 103530 650254
rect 113222 650254 122850 650314
rect 103470 650118 113098 650178
rect 93718 649982 93962 650042
rect 113038 650042 113098 650118
rect 113222 650042 113282 650254
rect 122790 650178 122850 650254
rect 132542 650254 142170 650314
rect 122790 650118 132418 650178
rect 113038 649982 113282 650042
rect 132358 650042 132418 650118
rect 132542 650042 132602 650254
rect 142110 650178 142170 650254
rect 151862 650254 161490 650314
rect 142110 650118 151738 650178
rect 132358 649982 132602 650042
rect 151678 650042 151738 650118
rect 151862 650042 151922 650254
rect 161430 650178 161490 650254
rect 171182 650254 180810 650314
rect 161430 650118 171058 650178
rect 151678 649982 151922 650042
rect 170998 650042 171058 650118
rect 171182 650042 171242 650254
rect 180750 650178 180810 650254
rect 190502 650254 200130 650314
rect 180750 650118 190378 650178
rect 170998 649982 171242 650042
rect 190318 650042 190378 650118
rect 190502 650042 190562 650254
rect 200070 650178 200130 650254
rect 209822 650254 219450 650314
rect 200070 650118 209698 650178
rect 190318 649982 190562 650042
rect 209638 650042 209698 650118
rect 209822 650042 209882 650254
rect 219390 650178 219450 650254
rect 229142 650254 238770 650314
rect 219390 650118 229018 650178
rect 209638 649982 209882 650042
rect 228958 650042 229018 650118
rect 229142 650042 229202 650254
rect 238710 650178 238770 650254
rect 248462 650254 258090 650314
rect 238710 650118 248338 650178
rect 228958 649982 229202 650042
rect 248278 650042 248338 650118
rect 248462 650042 248522 650254
rect 258030 650178 258090 650254
rect 267782 650254 277410 650314
rect 258030 650118 267658 650178
rect 248278 649982 248522 650042
rect 267598 650042 267658 650118
rect 267782 650042 267842 650254
rect 277350 650178 277410 650254
rect 287102 650254 292682 650314
rect 277350 650118 286978 650178
rect 267598 649982 267842 650042
rect 286918 650042 286978 650118
rect 287102 650042 287162 650254
rect 286918 649982 287162 650042
rect 292622 650042 292682 650254
rect 299422 650252 299428 650316
rect 299492 650314 299498 650316
rect 425053 650314 425119 650317
rect 540973 650314 541039 650317
rect 299492 650254 316050 650314
rect 299492 650252 299498 650254
rect 315990 650178 316050 650254
rect 325742 650254 335370 650314
rect 315990 650118 325618 650178
rect 299422 650042 299428 650044
rect 292622 649982 299428 650042
rect 299422 649980 299428 649982
rect 299492 649980 299498 650044
rect 325558 650042 325618 650118
rect 325742 650042 325802 650254
rect 335310 650178 335370 650254
rect 345062 650254 354690 650314
rect 335310 650118 344938 650178
rect 325558 649982 325802 650042
rect 344878 650042 344938 650118
rect 345062 650042 345122 650254
rect 354630 650178 354690 650254
rect 364382 650254 374010 650314
rect 354630 650118 364258 650178
rect 344878 649982 345122 650042
rect 364198 650042 364258 650118
rect 364382 650042 364442 650254
rect 373950 650178 374010 650254
rect 383702 650254 393330 650314
rect 373950 650118 383578 650178
rect 364198 649982 364442 650042
rect 383518 650042 383578 650118
rect 383702 650042 383762 650254
rect 393270 650178 393330 650254
rect 403022 650254 412650 650314
rect 393270 650118 402898 650178
rect 383518 649982 383762 650042
rect 402838 650042 402898 650118
rect 403022 650042 403082 650254
rect 412590 650178 412650 650254
rect 422342 650312 425119 650314
rect 422342 650256 425058 650312
rect 425114 650256 425119 650312
rect 422342 650254 425119 650256
rect 412590 650118 422218 650178
rect 402838 649982 403082 650042
rect 422158 650042 422218 650118
rect 422342 650042 422402 650254
rect 425053 650251 425119 650254
rect 437246 650254 451290 650314
rect 434529 650178 434595 650181
rect 437246 650178 437306 650254
rect 434529 650176 437306 650178
rect 434529 650120 434534 650176
rect 434590 650120 437306 650176
rect 434529 650118 437306 650120
rect 451230 650178 451290 650254
rect 460982 650254 470610 650314
rect 451230 650118 460858 650178
rect 434529 650115 434595 650118
rect 422158 649982 422402 650042
rect 460798 650042 460858 650118
rect 460982 650042 461042 650254
rect 470550 650178 470610 650254
rect 480302 650254 489930 650314
rect 470550 650118 480178 650178
rect 460798 649982 461042 650042
rect 480118 650042 480178 650118
rect 480302 650042 480362 650254
rect 489870 650178 489930 650254
rect 499622 650254 509250 650314
rect 489870 650118 499498 650178
rect 480118 649982 480362 650042
rect 499438 650042 499498 650118
rect 499622 650042 499682 650254
rect 509190 650178 509250 650254
rect 518942 650254 528570 650314
rect 509190 650118 518818 650178
rect 499438 649982 499682 650042
rect 518758 650042 518818 650118
rect 518942 650042 519002 650254
rect 528510 650178 528570 650254
rect 538262 650312 541039 650314
rect 538262 650256 540978 650312
rect 541034 650256 541039 650312
rect 538262 650254 541039 650256
rect 528510 650118 538138 650178
rect 518758 649982 519002 650042
rect 538078 650042 538138 650118
rect 538262 650042 538322 650254
rect 540973 650251 541039 650254
rect 565169 650314 565235 650317
rect 572713 650314 572779 650317
rect 565169 650312 569970 650314
rect 565169 650256 565174 650312
rect 565230 650256 569970 650312
rect 565169 650254 569970 650256
rect 565169 650251 565235 650254
rect 569910 650178 569970 650254
rect 572713 650312 576962 650314
rect 572713 650256 572718 650312
rect 572774 650256 576962 650312
rect 572713 650254 576962 650256
rect 572713 650251 572779 650254
rect 572621 650178 572687 650181
rect 569910 650176 572687 650178
rect 569910 650120 572626 650176
rect 572682 650120 572687 650176
rect 569910 650118 572687 650120
rect 576902 650178 576962 650254
rect 583342 650178 583402 651070
rect 583520 650980 584960 651070
rect 576902 650118 583402 650178
rect 572621 650115 572687 650118
rect 538078 649982 538322 650042
rect 548609 650042 548675 650045
rect 550582 650042 550588 650044
rect 548609 650040 550588 650042
rect 548609 649984 548614 650040
rect 548670 649984 550588 650040
rect 548609 649982 550588 649984
rect 548609 649979 548675 649982
rect 550582 649980 550588 649982
rect 550652 649980 550658 650044
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 583520 627738 584960 627828
rect 583342 627678 584960 627738
rect 550582 626996 550588 627060
rect 550652 627058 550658 627060
rect 553301 627058 553367 627061
rect 550652 627056 553367 627058
rect 550652 627000 553306 627056
rect 553362 627000 553367 627056
rect 550652 626998 553367 627000
rect 550652 626996 550658 626998
rect 553301 626995 553367 626998
rect 553485 627058 553551 627061
rect 560293 627058 560359 627061
rect 553485 627056 560359 627058
rect 553485 627000 553490 627056
rect 553546 627000 560298 627056
rect 560354 627000 560359 627056
rect 553485 626998 560359 627000
rect 553485 626995 553551 626998
rect 560293 626995 560359 626998
rect 58014 626860 58020 626924
rect 58084 626922 58090 626924
rect 289813 626922 289879 626925
rect 58084 626862 64890 626922
rect 58084 626860 58090 626862
rect 64830 626786 64890 626862
rect 74582 626862 84210 626922
rect 64830 626726 74458 626786
rect 74398 626650 74458 626726
rect 74582 626650 74642 626862
rect 84150 626786 84210 626862
rect 93902 626862 103530 626922
rect 84150 626726 93778 626786
rect 74398 626590 74642 626650
rect 93718 626650 93778 626726
rect 93902 626650 93962 626862
rect 103470 626786 103530 626862
rect 113222 626862 122850 626922
rect 103470 626726 113098 626786
rect 93718 626590 93962 626650
rect 113038 626650 113098 626726
rect 113222 626650 113282 626862
rect 122790 626786 122850 626862
rect 132542 626862 142170 626922
rect 122790 626726 132418 626786
rect 113038 626590 113282 626650
rect 132358 626650 132418 626726
rect 132542 626650 132602 626862
rect 142110 626786 142170 626862
rect 151862 626862 161490 626922
rect 142110 626726 151738 626786
rect 132358 626590 132602 626650
rect 151678 626650 151738 626726
rect 151862 626650 151922 626862
rect 161430 626786 161490 626862
rect 171182 626862 180810 626922
rect 161430 626726 171058 626786
rect 151678 626590 151922 626650
rect 170998 626650 171058 626726
rect 171182 626650 171242 626862
rect 180750 626786 180810 626862
rect 190502 626862 200130 626922
rect 180750 626726 190378 626786
rect 170998 626590 171242 626650
rect 190318 626650 190378 626726
rect 190502 626650 190562 626862
rect 200070 626786 200130 626862
rect 209822 626862 219450 626922
rect 200070 626726 209698 626786
rect 190318 626590 190562 626650
rect 209638 626650 209698 626726
rect 209822 626650 209882 626862
rect 219390 626786 219450 626862
rect 229142 626862 238770 626922
rect 219390 626726 229018 626786
rect 209638 626590 209882 626650
rect 228958 626650 229018 626726
rect 229142 626650 229202 626862
rect 238710 626786 238770 626862
rect 248462 626862 258090 626922
rect 238710 626726 248338 626786
rect 228958 626590 229202 626650
rect 248278 626650 248338 626726
rect 248462 626650 248522 626862
rect 258030 626786 258090 626862
rect 267782 626862 277410 626922
rect 258030 626726 267658 626786
rect 248278 626590 248522 626650
rect 267598 626650 267658 626726
rect 267782 626650 267842 626862
rect 277350 626786 277410 626862
rect 287102 626920 289879 626922
rect 287102 626864 289818 626920
rect 289874 626864 289879 626920
rect 287102 626862 289879 626864
rect 277350 626726 286978 626786
rect 267598 626590 267842 626650
rect 286918 626650 286978 626726
rect 287102 626650 287162 626862
rect 289813 626859 289879 626862
rect 299422 626860 299428 626924
rect 299492 626922 299498 626924
rect 425053 626922 425119 626925
rect 299492 626862 316050 626922
rect 299492 626860 299498 626862
rect 315990 626786 316050 626862
rect 325742 626862 335370 626922
rect 315990 626726 325618 626786
rect 286918 626590 287162 626650
rect 292665 626650 292731 626653
rect 299422 626650 299428 626652
rect 292665 626648 299428 626650
rect 292665 626592 292670 626648
rect 292726 626592 299428 626648
rect 292665 626590 299428 626592
rect 292665 626587 292731 626590
rect 299422 626588 299428 626590
rect 299492 626588 299498 626652
rect 325558 626650 325618 626726
rect 325742 626650 325802 626862
rect 335310 626786 335370 626862
rect 345062 626862 354690 626922
rect 335310 626726 344938 626786
rect 325558 626590 325802 626650
rect 344878 626650 344938 626726
rect 345062 626650 345122 626862
rect 354630 626786 354690 626862
rect 364382 626862 374010 626922
rect 354630 626726 364258 626786
rect 344878 626590 345122 626650
rect 364198 626650 364258 626726
rect 364382 626650 364442 626862
rect 373950 626786 374010 626862
rect 383702 626862 393330 626922
rect 373950 626726 383578 626786
rect 364198 626590 364442 626650
rect 383518 626650 383578 626726
rect 383702 626650 383762 626862
rect 393270 626786 393330 626862
rect 403022 626862 412650 626922
rect 393270 626726 402898 626786
rect 383518 626590 383762 626650
rect 402838 626650 402898 626726
rect 403022 626650 403082 626862
rect 412590 626786 412650 626862
rect 422342 626920 425119 626922
rect 422342 626864 425058 626920
rect 425114 626864 425119 626920
rect 422342 626862 425119 626864
rect 412590 626726 422218 626786
rect 402838 626590 403082 626650
rect 422158 626650 422218 626726
rect 422342 626650 422402 626862
rect 425053 626859 425119 626862
rect 434662 626860 434668 626924
rect 434732 626922 434738 626924
rect 540973 626922 541039 626925
rect 434732 626862 451290 626922
rect 434732 626860 434738 626862
rect 451230 626786 451290 626862
rect 460982 626862 470610 626922
rect 451230 626726 460858 626786
rect 422158 626590 422402 626650
rect 427905 626650 427971 626653
rect 434662 626650 434668 626652
rect 427905 626648 434668 626650
rect 427905 626592 427910 626648
rect 427966 626592 434668 626648
rect 427905 626590 434668 626592
rect 427905 626587 427971 626590
rect 434662 626588 434668 626590
rect 434732 626588 434738 626652
rect 460798 626650 460858 626726
rect 460982 626650 461042 626862
rect 470550 626786 470610 626862
rect 480302 626862 489930 626922
rect 470550 626726 480178 626786
rect 460798 626590 461042 626650
rect 480118 626650 480178 626726
rect 480302 626650 480362 626862
rect 489870 626786 489930 626862
rect 499622 626862 509250 626922
rect 489870 626726 499498 626786
rect 480118 626590 480362 626650
rect 499438 626650 499498 626726
rect 499622 626650 499682 626862
rect 509190 626786 509250 626862
rect 518942 626862 528570 626922
rect 509190 626726 518818 626786
rect 499438 626590 499682 626650
rect 518758 626650 518818 626726
rect 518942 626650 519002 626862
rect 528510 626786 528570 626862
rect 538262 626920 541039 626922
rect 538262 626864 540978 626920
rect 541034 626864 541039 626920
rect 538262 626862 541039 626864
rect 528510 626726 538138 626786
rect 518758 626590 519002 626650
rect 538078 626650 538138 626726
rect 538262 626650 538322 626862
rect 540973 626859 541039 626862
rect 565169 626922 565235 626925
rect 572713 626922 572779 626925
rect 565169 626920 569970 626922
rect 565169 626864 565174 626920
rect 565230 626864 569970 626920
rect 565169 626862 569970 626864
rect 565169 626859 565235 626862
rect 569910 626786 569970 626862
rect 572713 626920 576962 626922
rect 572713 626864 572718 626920
rect 572774 626864 576962 626920
rect 572713 626862 576962 626864
rect 572713 626859 572779 626862
rect 572621 626786 572687 626789
rect 569910 626784 572687 626786
rect 569910 626728 572626 626784
rect 572682 626728 572687 626784
rect 569910 626726 572687 626728
rect 576902 626786 576962 626862
rect 583342 626786 583402 627678
rect 583520 627588 584960 627678
rect 576902 626726 583402 626786
rect 572621 626723 572687 626726
rect 538078 626590 538322 626650
rect 548609 626650 548675 626653
rect 550582 626650 550588 626652
rect 548609 626648 550588 626650
rect 548609 626592 548614 626648
rect 548670 626592 550588 626648
rect 548609 626590 550588 626592
rect 548609 626587 548675 626590
rect 550582 626588 550588 626590
rect 550652 626588 550658 626652
rect -960 624882 480 624972
rect 4061 624882 4127 624885
rect -960 624880 4127 624882
rect -960 624824 4066 624880
rect 4122 624824 4127 624880
rect -960 624822 4127 624824
rect -960 624732 480 624822
rect 4061 624819 4127 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 559097 608698 559163 608701
rect 559373 608698 559439 608701
rect 559097 608696 559439 608698
rect 559097 608640 559102 608696
rect 559158 608640 559378 608696
rect 559434 608640 559439 608696
rect 559097 608638 559439 608640
rect 559097 608635 559163 608638
rect 559373 608635 559439 608638
rect 583520 604210 584960 604300
rect 583342 604150 584960 604210
rect 553393 603530 553459 603533
rect 560293 603530 560359 603533
rect 553393 603528 560359 603530
rect 553393 603472 553398 603528
rect 553454 603472 560298 603528
rect 560354 603472 560359 603528
rect 553393 603470 560359 603472
rect 553393 603467 553459 603470
rect 560293 603467 560359 603470
rect 59721 603394 59787 603397
rect 289813 603394 289879 603397
rect 59721 603392 64890 603394
rect 59721 603336 59726 603392
rect 59782 603336 64890 603392
rect 59721 603334 64890 603336
rect 59721 603331 59787 603334
rect 64830 603258 64890 603334
rect 74582 603334 84210 603394
rect 64830 603198 74458 603258
rect 74398 603122 74458 603198
rect 74582 603122 74642 603334
rect 84150 603258 84210 603334
rect 93902 603334 103530 603394
rect 84150 603198 93778 603258
rect 74398 603062 74642 603122
rect 93718 603122 93778 603198
rect 93902 603122 93962 603334
rect 103470 603258 103530 603334
rect 113222 603334 122850 603394
rect 103470 603198 113098 603258
rect 93718 603062 93962 603122
rect 113038 603122 113098 603198
rect 113222 603122 113282 603334
rect 122790 603258 122850 603334
rect 132542 603334 142170 603394
rect 122790 603198 132418 603258
rect 113038 603062 113282 603122
rect 132358 603122 132418 603198
rect 132542 603122 132602 603334
rect 142110 603258 142170 603334
rect 151862 603334 161490 603394
rect 142110 603198 151738 603258
rect 132358 603062 132602 603122
rect 151678 603122 151738 603198
rect 151862 603122 151922 603334
rect 161430 603258 161490 603334
rect 171182 603334 180810 603394
rect 161430 603198 171058 603258
rect 151678 603062 151922 603122
rect 170998 603122 171058 603198
rect 171182 603122 171242 603334
rect 180750 603258 180810 603334
rect 190502 603334 200130 603394
rect 180750 603198 190378 603258
rect 170998 603062 171242 603122
rect 190318 603122 190378 603198
rect 190502 603122 190562 603334
rect 200070 603258 200130 603334
rect 209822 603334 219450 603394
rect 200070 603198 209698 603258
rect 190318 603062 190562 603122
rect 209638 603122 209698 603198
rect 209822 603122 209882 603334
rect 219390 603258 219450 603334
rect 229142 603334 238770 603394
rect 219390 603198 229018 603258
rect 209638 603062 209882 603122
rect 228958 603122 229018 603198
rect 229142 603122 229202 603334
rect 238710 603258 238770 603334
rect 248462 603334 258090 603394
rect 238710 603198 248338 603258
rect 228958 603062 229202 603122
rect 248278 603122 248338 603198
rect 248462 603122 248522 603334
rect 258030 603258 258090 603334
rect 267782 603334 277410 603394
rect 258030 603198 267658 603258
rect 248278 603062 248522 603122
rect 267598 603122 267658 603198
rect 267782 603122 267842 603334
rect 277350 603258 277410 603334
rect 287102 603392 289879 603394
rect 287102 603336 289818 603392
rect 289874 603336 289879 603392
rect 287102 603334 289879 603336
rect 277350 603198 286978 603258
rect 267598 603062 267842 603122
rect 286918 603122 286978 603198
rect 287102 603122 287162 603334
rect 289813 603331 289879 603334
rect 299422 603332 299428 603396
rect 299492 603394 299498 603396
rect 425053 603394 425119 603397
rect 299492 603334 316050 603394
rect 299492 603332 299498 603334
rect 315990 603258 316050 603334
rect 325742 603334 335370 603394
rect 315990 603198 325618 603258
rect 286918 603062 287162 603122
rect 292665 603122 292731 603125
rect 299422 603122 299428 603124
rect 292665 603120 299428 603122
rect 292665 603064 292670 603120
rect 292726 603064 299428 603120
rect 292665 603062 299428 603064
rect 292665 603059 292731 603062
rect 299422 603060 299428 603062
rect 299492 603060 299498 603124
rect 325558 603122 325618 603198
rect 325742 603122 325802 603334
rect 335310 603258 335370 603334
rect 345062 603334 354690 603394
rect 335310 603198 344938 603258
rect 325558 603062 325802 603122
rect 344878 603122 344938 603198
rect 345062 603122 345122 603334
rect 354630 603258 354690 603334
rect 364382 603334 374010 603394
rect 354630 603198 364258 603258
rect 344878 603062 345122 603122
rect 364198 603122 364258 603198
rect 364382 603122 364442 603334
rect 373950 603258 374010 603334
rect 383702 603334 393330 603394
rect 373950 603198 383578 603258
rect 364198 603062 364442 603122
rect 383518 603122 383578 603198
rect 383702 603122 383762 603334
rect 393270 603258 393330 603334
rect 403022 603392 425119 603394
rect 403022 603336 425058 603392
rect 425114 603336 425119 603392
rect 403022 603334 425119 603336
rect 393270 603198 402898 603258
rect 383518 603062 383762 603122
rect 402838 603122 402898 603198
rect 403022 603122 403082 603334
rect 425053 603331 425119 603334
rect 441521 603394 441587 603397
rect 540973 603394 541039 603397
rect 441521 603392 451290 603394
rect 441521 603336 441526 603392
rect 441582 603336 451290 603392
rect 441521 603334 451290 603336
rect 441521 603331 441587 603334
rect 429929 603258 429995 603261
rect 434662 603258 434668 603260
rect 429929 603256 434668 603258
rect 429929 603200 429934 603256
rect 429990 603200 434668 603256
rect 429929 603198 434668 603200
rect 429929 603195 429995 603198
rect 434662 603196 434668 603198
rect 434732 603196 434738 603260
rect 451230 603258 451290 603334
rect 460982 603334 470610 603394
rect 451230 603198 460858 603258
rect 402838 603062 403082 603122
rect 460798 603122 460858 603198
rect 460982 603122 461042 603334
rect 470550 603258 470610 603334
rect 480302 603334 489930 603394
rect 470550 603198 480178 603258
rect 460798 603062 461042 603122
rect 480118 603122 480178 603198
rect 480302 603122 480362 603334
rect 489870 603258 489930 603334
rect 499622 603334 509250 603394
rect 489870 603198 499498 603258
rect 480118 603062 480362 603122
rect 499438 603122 499498 603198
rect 499622 603122 499682 603334
rect 509190 603258 509250 603334
rect 518942 603334 528570 603394
rect 509190 603198 518818 603258
rect 499438 603062 499682 603122
rect 518758 603122 518818 603198
rect 518942 603122 519002 603334
rect 528510 603258 528570 603334
rect 538262 603392 541039 603394
rect 538262 603336 540978 603392
rect 541034 603336 541039 603392
rect 538262 603334 541039 603336
rect 528510 603198 538138 603258
rect 518758 603062 519002 603122
rect 538078 603122 538138 603198
rect 538262 603122 538322 603334
rect 540973 603331 541039 603334
rect 565169 603394 565235 603397
rect 572713 603394 572779 603397
rect 565169 603392 569970 603394
rect 565169 603336 565174 603392
rect 565230 603336 569970 603392
rect 565169 603334 569970 603336
rect 565169 603331 565235 603334
rect 569910 603258 569970 603334
rect 572713 603392 576962 603394
rect 572713 603336 572718 603392
rect 572774 603336 576962 603392
rect 572713 603334 576962 603336
rect 572713 603331 572779 603334
rect 572621 603258 572687 603261
rect 569910 603256 572687 603258
rect 569910 603200 572626 603256
rect 572682 603200 572687 603256
rect 569910 603198 572687 603200
rect 576902 603258 576962 603334
rect 583342 603258 583402 604150
rect 583520 604060 584960 604150
rect 576902 603198 583402 603258
rect 572621 603195 572687 603198
rect 538078 603062 538322 603122
rect 548609 603122 548675 603125
rect 553301 603122 553367 603125
rect 548609 603120 553367 603122
rect 548609 603064 548614 603120
rect 548670 603064 553306 603120
rect 553362 603064 553367 603120
rect 548609 603062 553367 603064
rect 548609 603059 548675 603062
rect 553301 603059 553367 603062
rect 434662 602924 434668 602988
rect 434732 602986 434738 602988
rect 441521 602986 441587 602989
rect 434732 602984 441587 602986
rect 434732 602928 441526 602984
rect 441582 602928 441587 602984
rect 434732 602926 441587 602928
rect 434732 602924 434738 602926
rect 441521 602923 441587 602926
rect 59721 596322 59787 596325
rect 59126 596320 59787 596322
rect 59126 596264 59726 596320
rect 59782 596264 59787 596320
rect 59126 596262 59787 596264
rect 59126 596186 59186 596262
rect 59721 596259 59787 596262
rect 59486 596186 59492 596188
rect -960 596050 480 596140
rect 59126 596126 59492 596186
rect 59486 596124 59492 596126
rect 59556 596124 59562 596188
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 59302 581572 59308 581636
rect 59372 581634 59378 581636
rect 59854 581634 59860 581636
rect 59372 581574 59860 581634
rect 59372 581572 59378 581574
rect 59854 581572 59860 581574
rect 59924 581572 59930 581636
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 59813 579596 59879 579597
rect 59813 579594 59860 579596
rect 59768 579592 59860 579594
rect 59768 579536 59818 579592
rect 59768 579534 59860 579536
rect 59813 579532 59860 579534
rect 59924 579532 59930 579596
rect 59813 579531 59879 579532
rect 59813 570210 59879 570213
rect 59678 570208 59879 570210
rect 59678 570152 59818 570208
rect 59874 570152 59879 570208
rect 59678 570150 59879 570152
rect 59678 570076 59738 570150
rect 59813 570147 59879 570150
rect 59670 570012 59676 570076
rect 59740 570012 59746 570076
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 59670 563274 59676 563276
rect 59494 563214 59676 563274
rect 59494 563004 59554 563214
rect 59670 563212 59676 563214
rect 59740 563212 59746 563276
rect 59486 562940 59492 563004
rect 59556 562940 59562 563004
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect 133689 553484 133755 553485
rect 259177 553484 259243 553485
rect 263777 553484 263843 553485
rect 133638 553482 133644 553484
rect 133598 553422 133644 553482
rect 133708 553480 133755 553484
rect 259126 553482 259132 553484
rect 133750 553424 133755 553480
rect 133638 553420 133644 553422
rect 133708 553420 133755 553424
rect 259086 553422 259132 553482
rect 259196 553480 259243 553484
rect 263726 553482 263732 553484
rect 259238 553424 259243 553480
rect 259126 553420 259132 553422
rect 259196 553420 259243 553424
rect 263686 553422 263732 553482
rect 263796 553480 263843 553484
rect 263838 553424 263843 553480
rect 263726 553420 263732 553422
rect 263796 553420 263843 553424
rect 133689 553419 133755 553420
rect 259177 553419 259243 553420
rect 263777 553419 263843 553420
rect 378501 553484 378567 553485
rect 382917 553484 382983 553485
rect 507853 553484 507919 553485
rect 513373 553484 513439 553485
rect 378501 553480 378548 553484
rect 378612 553482 378618 553484
rect 378501 553424 378506 553480
rect 378501 553420 378548 553424
rect 378612 553422 378658 553482
rect 382917 553480 382964 553484
rect 383028 553482 383034 553484
rect 382917 553424 382922 553480
rect 378612 553420 378618 553422
rect 382917 553420 382964 553424
rect 383028 553422 383074 553482
rect 507853 553480 507900 553484
rect 507964 553482 507970 553484
rect 507853 553424 507858 553480
rect 383028 553420 383034 553422
rect 507853 553420 507900 553424
rect 507964 553422 508010 553482
rect 513373 553480 513420 553484
rect 513484 553482 513490 553484
rect 513373 553424 513378 553480
rect 507964 553420 507970 553422
rect 513373 553420 513420 553424
rect 513484 553422 513530 553482
rect 513484 553420 513490 553422
rect 378501 553419 378567 553420
rect 382917 553419 382983 553420
rect 507853 553419 507919 553420
rect 513373 553419 513439 553420
rect -960 553074 480 553164
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 129222 551108 129228 551172
rect 129292 551170 129298 551172
rect 132902 551170 132908 551172
rect 129292 551110 132908 551170
rect 129292 551108 129298 551110
rect 132902 551108 132908 551110
rect 132972 551108 132978 551172
rect 514150 550700 514156 550764
rect 514220 550762 514226 550764
rect 518893 550762 518959 550765
rect 514220 550760 518959 550762
rect 514220 550704 518898 550760
rect 518954 550704 518959 550760
rect 514220 550702 518959 550704
rect 514220 550700 514226 550702
rect 518893 550699 518959 550702
rect 139393 549946 139459 549949
rect 137142 549944 139459 549946
rect 137142 549888 139398 549944
rect 139454 549888 139459 549944
rect 137142 549886 139459 549888
rect 137142 549683 137202 549886
rect 139393 549883 139459 549886
rect 266445 549946 266511 549949
rect 389173 549946 389239 549949
rect 266445 549944 266554 549946
rect 266445 549888 266450 549944
rect 266506 549888 266554 549944
rect 266445 549883 266554 549888
rect 266494 549402 266554 549883
rect 387198 549944 389239 549946
rect 387198 549888 389178 549944
rect 389234 549888 389239 549944
rect 387198 549886 389239 549888
rect 387198 549683 387258 549886
rect 389173 549883 389239 549886
rect 516409 549946 516475 549949
rect 516409 549944 516610 549946
rect 516409 549888 516414 549944
rect 516470 549888 516610 549944
rect 516409 549886 516610 549888
rect 516409 549883 516475 549886
rect 516550 549683 516610 549886
rect 270401 549402 270467 549405
rect 266494 549400 270467 549402
rect 266494 549344 270406 549400
rect 270462 549344 270467 549400
rect 266494 549342 270467 549344
rect 270401 549339 270467 549342
rect 59494 546557 60076 546617
rect 189582 546557 190164 546617
rect 309550 546557 310132 546617
rect 439454 546557 440036 546617
rect 57513 546546 57579 546549
rect 59494 546546 59554 546557
rect 57513 546544 59554 546546
rect 57513 546488 57518 546544
rect 57574 546488 59554 546544
rect 57513 546486 59554 546488
rect 187693 546546 187759 546549
rect 189582 546546 189642 546557
rect 187693 546544 189642 546546
rect 187693 546488 187698 546544
rect 187754 546488 189642 546544
rect 187693 546486 189642 546488
rect 305821 546546 305887 546549
rect 309550 546546 309610 546557
rect 305821 546544 309610 546546
rect 305821 546488 305826 546544
rect 305882 546488 309610 546544
rect 305821 546486 309610 546488
rect 437473 546546 437539 546549
rect 439454 546546 439514 546557
rect 437473 546544 439514 546546
rect 437473 546488 437478 546544
rect 437534 546488 439514 546544
rect 437473 546486 439514 546488
rect 57513 546483 57579 546486
rect 187693 546483 187759 546486
rect 305821 546483 305887 546486
rect 437473 546483 437539 546486
rect 580257 545594 580323 545597
rect 583520 545594 584960 545684
rect 580257 545592 584960 545594
rect 580257 545536 580262 545592
rect 580318 545536 584960 545592
rect 580257 545534 584960 545536
rect 580257 545531 580323 545534
rect 57421 545186 57487 545189
rect 60046 545186 60106 545459
rect 57421 545184 60106 545186
rect 57421 545128 57426 545184
rect 57482 545128 60106 545184
rect 57421 545126 60106 545128
rect 187693 545186 187759 545189
rect 190134 545186 190194 545459
rect 187693 545184 190194 545186
rect 187693 545128 187698 545184
rect 187754 545128 190194 545184
rect 187693 545126 190194 545128
rect 307661 545186 307727 545189
rect 310102 545186 310162 545459
rect 307661 545184 310162 545186
rect 307661 545128 307666 545184
rect 307722 545128 310162 545184
rect 307661 545126 310162 545128
rect 437473 545186 437539 545189
rect 440006 545186 440066 545459
rect 583520 545444 584960 545534
rect 437473 545184 440066 545186
rect 437473 545128 437478 545184
rect 437534 545128 440066 545184
rect 437473 545126 440066 545128
rect 57421 545123 57487 545126
rect 187693 545123 187759 545126
rect 307661 545123 307727 545126
rect 437473 545123 437539 545126
rect 56869 543826 56935 543829
rect 187693 543826 187759 543829
rect 305729 543826 305795 543829
rect 429561 543826 429627 543829
rect 56869 543824 60106 543826
rect 56869 543768 56874 543824
rect 56930 543768 60106 543824
rect 56869 543766 60106 543768
rect 56869 543763 56935 543766
rect 60046 543759 60106 543766
rect 187693 543824 190194 543826
rect 187693 543768 187698 543824
rect 187754 543768 190194 543824
rect 187693 543766 190194 543768
rect 187693 543763 187759 543766
rect 190134 543759 190194 543766
rect 305729 543824 310162 543826
rect 305729 543768 305734 543824
rect 305790 543768 310162 543824
rect 305729 543766 310162 543768
rect 305729 543763 305795 543766
rect 310102 543759 310162 543766
rect 429518 543824 429627 543826
rect 429518 543768 429566 543824
rect 429622 543768 429627 543824
rect 429518 543763 429627 543768
rect 437473 543826 437539 543829
rect 437473 543824 440066 543826
rect 437473 543768 437478 543824
rect 437534 543768 440066 543824
rect 437473 543766 440066 543768
rect 437473 543763 437539 543766
rect 429377 543690 429443 543693
rect 429518 543690 429578 543763
rect 440006 543759 440066 543766
rect 429377 543688 429578 543690
rect 429377 543632 429382 543688
rect 429438 543632 429578 543688
rect 429377 543630 429578 543632
rect 429377 543627 429443 543630
rect 57329 542466 57395 542469
rect 60046 542466 60106 542631
rect 187693 542602 187759 542605
rect 190134 542602 190194 542631
rect 187693 542600 190194 542602
rect 187693 542544 187698 542600
rect 187754 542544 190194 542600
rect 187693 542542 190194 542544
rect 187693 542539 187759 542542
rect 57329 542464 60106 542466
rect 57329 542408 57334 542464
rect 57390 542408 60106 542464
rect 57329 542406 60106 542408
rect 307201 542466 307267 542469
rect 310102 542466 310162 542631
rect 307201 542464 310162 542466
rect 307201 542408 307206 542464
rect 307262 542408 310162 542464
rect 307201 542406 310162 542408
rect 437473 542466 437539 542469
rect 440006 542466 440066 542631
rect 437473 542464 440066 542466
rect 437473 542408 437478 542464
rect 437534 542408 440066 542464
rect 437473 542406 440066 542408
rect 57329 542403 57395 542406
rect 307201 542403 307267 542406
rect 437473 542403 437539 542406
rect 429193 540970 429259 540973
rect 429377 540970 429443 540973
rect 429193 540968 429443 540970
rect 56777 540426 56843 540429
rect 60046 540426 60106 540931
rect 56777 540424 60106 540426
rect 56777 540368 56782 540424
rect 56838 540368 60106 540424
rect 56777 540366 60106 540368
rect 187785 540426 187851 540429
rect 190134 540426 190194 540931
rect 187785 540424 190194 540426
rect 187785 540368 187790 540424
rect 187846 540368 190194 540424
rect 187785 540366 190194 540368
rect 307293 540426 307359 540429
rect 310102 540426 310162 540931
rect 429193 540912 429198 540968
rect 429254 540912 429382 540968
rect 429438 540912 429443 540968
rect 429193 540910 429443 540912
rect 429193 540907 429259 540910
rect 429377 540907 429443 540910
rect 307293 540424 310162 540426
rect 307293 540368 307298 540424
rect 307354 540368 310162 540424
rect 307293 540366 310162 540368
rect 437565 540426 437631 540429
rect 440006 540426 440066 540931
rect 437565 540424 440066 540426
rect 437565 540368 437570 540424
rect 437626 540368 440066 540424
rect 437565 540366 440066 540368
rect 56777 540363 56843 540366
rect 187785 540363 187851 540366
rect 307293 540363 307359 540366
rect 437565 540363 437631 540366
rect 187693 539882 187759 539885
rect 307661 539882 307727 539885
rect 437473 539882 437539 539885
rect 187693 539880 190194 539882
rect 187693 539824 187698 539880
rect 187754 539824 190194 539880
rect 187693 539822 190194 539824
rect 187693 539819 187759 539822
rect 190134 539803 190194 539822
rect 307661 539880 310162 539882
rect 307661 539824 307666 539880
rect 307722 539824 310162 539880
rect 307661 539822 310162 539824
rect 307661 539819 307727 539822
rect 310102 539803 310162 539822
rect 437473 539880 440066 539882
rect 437473 539824 437478 539880
rect 437534 539824 440066 539880
rect 437473 539822 440066 539824
rect 437473 539819 437539 539822
rect 440006 539803 440066 539822
rect 57145 539610 57211 539613
rect 60046 539610 60106 539803
rect 57145 539608 60106 539610
rect 57145 539552 57150 539608
rect 57206 539552 60106 539608
rect 57145 539550 60106 539552
rect 305637 539610 305703 539613
rect 307293 539610 307359 539613
rect 305637 539608 307359 539610
rect 305637 539552 305642 539608
rect 305698 539552 307298 539608
rect 307354 539552 307359 539608
rect 305637 539550 307359 539552
rect 57145 539547 57211 539550
rect 305637 539547 305703 539550
rect 307293 539547 307359 539550
rect -960 538658 480 538748
rect 3601 538658 3667 538661
rect -960 538656 3667 538658
rect -960 538600 3606 538656
rect 3662 538600 3667 538656
rect -960 538598 3667 538600
rect -960 538508 480 538598
rect 3601 538595 3667 538598
rect 57053 537570 57119 537573
rect 60046 537570 60106 538103
rect 57053 537568 60106 537570
rect 57053 537512 57058 537568
rect 57114 537512 60106 537568
rect 57053 537510 60106 537512
rect 188337 537570 188403 537573
rect 190134 537570 190194 538103
rect 188337 537568 190194 537570
rect 188337 537512 188342 537568
rect 188398 537512 190194 537568
rect 188337 537510 190194 537512
rect 307017 537570 307083 537573
rect 310102 537570 310162 538103
rect 307017 537568 310162 537570
rect 307017 537512 307022 537568
rect 307078 537512 310162 537568
rect 307017 537510 310162 537512
rect 437473 537570 437539 537573
rect 440006 537570 440066 538103
rect 437473 537568 440066 537570
rect 437473 537512 437478 537568
rect 437534 537512 440066 537568
rect 437473 537510 440066 537512
rect 57053 537507 57119 537510
rect 188337 537507 188403 537510
rect 307017 537507 307083 537510
rect 437473 537507 437539 537510
rect 580349 533898 580415 533901
rect 583520 533898 584960 533988
rect 580349 533896 584960 533898
rect 580349 533840 580354 533896
rect 580410 533840 584960 533896
rect 580349 533838 584960 533840
rect 580349 533835 580415 533838
rect 583520 533748 584960 533838
rect 299473 531314 299539 531317
rect 299657 531314 299723 531317
rect 299473 531312 299723 531314
rect 299473 531256 299478 531312
rect 299534 531256 299662 531312
rect 299718 531256 299723 531312
rect 299473 531254 299723 531256
rect 299473 531251 299539 531254
rect 299657 531251 299723 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 429377 521658 429443 521661
rect 429561 521658 429627 521661
rect 429377 521656 429627 521658
rect 429377 521600 429382 521656
rect 429438 521600 429566 521656
rect 429622 521600 429627 521656
rect 429377 521598 429627 521600
rect 429377 521595 429443 521598
rect 429561 521595 429627 521598
rect 559097 521658 559163 521661
rect 559281 521658 559347 521661
rect 559097 521656 559347 521658
rect 559097 521600 559102 521656
rect 559158 521600 559286 521656
rect 559342 521600 559347 521656
rect 559097 521598 559347 521600
rect 559097 521595 559163 521598
rect 559281 521595 559347 521598
rect 299473 512002 299539 512005
rect 299657 512002 299723 512005
rect 299473 512000 299723 512002
rect 299473 511944 299478 512000
rect 299534 511944 299662 512000
rect 299718 511944 299723 512000
rect 299473 511942 299723 511944
rect 299473 511939 299539 511942
rect 299657 511939 299723 511942
rect 580441 510370 580507 510373
rect 583520 510370 584960 510460
rect 580441 510368 584960 510370
rect 580441 510312 580446 510368
rect 580502 510312 584960 510368
rect 580441 510310 584960 510312
rect 580441 510307 580507 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3693 509962 3759 509965
rect -960 509960 3759 509962
rect -960 509904 3698 509960
rect 3754 509904 3759 509960
rect -960 509902 3759 509904
rect -960 509812 480 509902
rect 3693 509899 3759 509902
rect 580533 498674 580599 498677
rect 583520 498674 584960 498764
rect 580533 498672 584960 498674
rect 580533 498616 580538 498672
rect 580594 498616 584960 498672
rect 580533 498614 584960 498616
rect 580533 498611 580599 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3785 495546 3851 495549
rect -960 495544 3851 495546
rect -960 495488 3790 495544
rect 3846 495488 3851 495544
rect -960 495486 3851 495488
rect -960 495396 480 495486
rect 3785 495483 3851 495486
rect 559189 492826 559255 492829
rect 559054 492824 559255 492826
rect 559054 492768 559194 492824
rect 559250 492768 559255 492824
rect 559054 492766 559255 492768
rect 559054 492693 559114 492766
rect 559189 492763 559255 492766
rect 559054 492688 559163 492693
rect 559054 492632 559102 492688
rect 559158 492632 559163 492688
rect 559054 492630 559163 492632
rect 559097 492627 559163 492630
rect 139393 489562 139459 489565
rect 389173 489562 389239 489565
rect 518893 489562 518959 489565
rect 137142 489560 139459 489562
rect 137142 489504 139398 489560
rect 139454 489504 139459 489560
rect 137142 489502 139459 489504
rect -960 481130 480 481220
rect 2957 481130 3023 481133
rect -960 481128 3023 481130
rect -960 481072 2962 481128
rect 3018 481072 3023 481128
rect -960 481070 3023 481072
rect -960 480980 480 481070
rect 2957 481067 3023 481070
rect 137142 480928 137202 489502
rect 139393 489499 139459 489502
rect 387198 489560 389239 489562
rect 387198 489504 389178 489560
rect 389234 489504 389239 489560
rect 387198 489502 389239 489504
rect 266678 484914 266738 489412
rect 266678 484884 267260 484914
rect 266708 484854 267290 484884
rect 267230 484530 267290 484854
rect 269113 484530 269179 484533
rect 267230 484528 269179 484530
rect 267230 484472 269118 484528
rect 269174 484472 269179 484528
rect 267230 484470 269179 484472
rect 267230 480928 267290 484470
rect 269113 484467 269179 484470
rect 299473 483034 299539 483037
rect 299749 483034 299815 483037
rect 299473 483032 299815 483034
rect 299473 482976 299478 483032
rect 299534 482976 299754 483032
rect 299810 482976 299815 483032
rect 299473 482974 299815 482976
rect 299473 482971 299539 482974
rect 299749 482971 299815 482974
rect 387198 480994 387258 489502
rect 389173 489499 389239 489502
rect 517102 489560 518959 489562
rect 517102 489504 518898 489560
rect 518954 489504 518959 489560
rect 517102 489502 518959 489504
rect 517102 484914 517162 489502
rect 518893 489499 518959 489502
rect 580717 486842 580783 486845
rect 583520 486842 584960 486932
rect 580717 486840 584960 486842
rect 580717 486784 580722 486840
rect 580778 486784 584960 486840
rect 580717 486782 584960 486784
rect 580717 486779 580783 486782
rect 583520 486692 584960 486782
rect 516580 484884 517162 484914
rect 516550 484854 517132 484884
rect 389173 480994 389239 480997
rect 387198 480992 389239 480994
rect 387198 480936 389178 480992
rect 389234 480936 389239 480992
rect 387198 480934 389239 480936
rect 387198 480928 387258 480934
rect 389173 480931 389239 480934
rect 516550 480928 516610 484854
rect 56961 480314 57027 480317
rect 188981 480314 189047 480317
rect 305913 480314 305979 480317
rect 437473 480314 437539 480317
rect 56961 480312 60106 480314
rect 56961 480256 56966 480312
rect 57022 480256 60106 480312
rect 56961 480254 60106 480256
rect 188981 480312 190194 480314
rect 188981 480256 188986 480312
rect 189042 480256 190194 480312
rect 188981 480254 190194 480256
rect 305913 480312 310162 480314
rect 305913 480256 305918 480312
rect 305974 480256 310162 480312
rect 305913 480254 310162 480256
rect 437473 480312 440066 480314
rect 437473 480256 437478 480312
rect 437534 480256 440066 480312
rect 437473 480254 440066 480256
rect 56961 480251 57027 480254
rect 188981 480251 189047 480254
rect 305913 480251 305979 480254
rect 437473 480251 437539 480254
rect 59813 478585 59879 478588
rect 59813 478583 60076 478585
rect 59813 478527 59818 478583
rect 59874 478527 60076 478583
rect 59813 478525 60076 478527
rect 59813 478522 59879 478525
rect 188889 478002 188955 478005
rect 190134 478002 190194 478555
rect 307109 478138 307175 478141
rect 310102 478138 310162 478555
rect 307109 478136 310162 478138
rect 307109 478080 307114 478136
rect 307170 478080 310162 478136
rect 307109 478078 310162 478080
rect 307109 478075 307175 478078
rect 188889 478000 190194 478002
rect 188889 477944 188894 478000
rect 188950 477944 190194 478000
rect 188889 477942 190194 477944
rect 438117 478002 438183 478005
rect 440006 478002 440066 478555
rect 438117 478000 440066 478002
rect 438117 477944 438122 478000
rect 438178 477944 440066 478000
rect 438117 477942 440066 477944
rect 188889 477939 188955 477942
rect 438117 477939 438183 477942
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 429469 463722 429535 463725
rect 429653 463722 429719 463725
rect 429469 463720 429719 463722
rect 429469 463664 429474 463720
rect 429530 463664 429658 463720
rect 429714 463664 429719 463720
rect 429469 463662 429719 463664
rect 429469 463659 429535 463662
rect 429653 463659 429719 463662
rect 580809 463450 580875 463453
rect 583520 463450 584960 463540
rect 580809 463448 584960 463450
rect 580809 463392 580814 463448
rect 580870 463392 584960 463448
rect 580809 463390 584960 463392
rect 580809 463387 580875 463390
rect 583520 463300 584960 463390
rect 351821 459644 351887 459645
rect 351821 459642 351840 459644
rect 351748 459640 351840 459642
rect 351748 459584 351826 459640
rect 351748 459582 351840 459584
rect 351821 459580 351840 459582
rect 351904 459580 351910 459644
rect 351821 459579 351887 459580
rect 77293 459508 77359 459509
rect 77293 459506 77312 459508
rect 77220 459504 77312 459506
rect 77220 459448 77298 459504
rect 77220 459446 77312 459448
rect 77293 459444 77312 459446
rect 77376 459444 77382 459508
rect 327306 459444 327312 459508
rect 327376 459506 327382 459508
rect 327901 459506 327967 459509
rect 358813 459508 358879 459509
rect 483013 459508 483079 459509
rect 327376 459504 327967 459506
rect 327376 459448 327906 459504
rect 327962 459448 327967 459504
rect 327376 459446 327967 459448
rect 327376 459444 327382 459446
rect 77293 459443 77359 459444
rect 327901 459443 327967 459446
rect 328474 459444 328480 459508
rect 328544 459506 328550 459508
rect 328862 459506 328868 459508
rect 328544 459446 328868 459506
rect 328544 459444 328550 459446
rect 328862 459444 328868 459446
rect 328932 459444 328938 459508
rect 358813 459506 358848 459508
rect 358756 459504 358848 459506
rect 358756 459448 358818 459504
rect 358756 459446 358848 459448
rect 358813 459444 358848 459446
rect 358912 459444 358918 459508
rect 452634 459444 452640 459508
rect 452704 459506 452710 459508
rect 453062 459506 453068 459508
rect 452704 459446 453068 459506
rect 452704 459444 452710 459446
rect 453062 459444 453068 459446
rect 453132 459444 453138 459508
rect 483002 459444 483008 459508
rect 483072 459506 483079 459508
rect 483072 459504 483164 459506
rect 483074 459448 483164 459504
rect 483072 459446 483164 459448
rect 483072 459444 483079 459446
rect 358813 459443 358879 459444
rect 483013 459443 483079 459444
rect 73838 458084 73844 458148
rect 73908 458146 73914 458148
rect 74165 458146 74231 458149
rect 73908 458144 74231 458146
rect 73908 458088 74170 458144
rect 74226 458088 74231 458144
rect 73908 458086 74231 458088
rect 73908 458084 73914 458086
rect 74165 458083 74231 458086
rect 74942 458084 74948 458148
rect 75012 458146 75018 458148
rect 75821 458146 75887 458149
rect 75012 458144 75887 458146
rect 75012 458088 75826 458144
rect 75882 458088 75887 458144
rect 75012 458086 75887 458088
rect 75012 458084 75018 458086
rect 75821 458083 75887 458086
rect 79358 458084 79364 458148
rect 79428 458146 79434 458148
rect 79961 458146 80027 458149
rect 79428 458144 80027 458146
rect 79428 458088 79966 458144
rect 80022 458088 80027 458144
rect 79428 458086 80027 458088
rect 79428 458084 79434 458086
rect 79961 458083 80027 458086
rect 81893 458148 81959 458149
rect 82813 458148 82879 458149
rect 84193 458148 84259 458149
rect 85481 458148 85547 458149
rect 81893 458144 81940 458148
rect 82004 458146 82010 458148
rect 81893 458088 81898 458144
rect 81893 458084 81940 458088
rect 82004 458086 82050 458146
rect 82813 458144 82860 458148
rect 82924 458146 82930 458148
rect 82813 458088 82818 458144
rect 82004 458084 82010 458086
rect 82813 458084 82860 458088
rect 82924 458086 82970 458146
rect 82924 458084 82930 458086
rect 84142 458084 84148 458148
rect 84212 458146 84259 458148
rect 85430 458146 85436 458148
rect 84212 458144 84304 458146
rect 84254 458088 84304 458144
rect 84212 458086 84304 458088
rect 85390 458086 85436 458146
rect 85500 458144 85547 458148
rect 85542 458088 85547 458144
rect 84212 458084 84259 458086
rect 85430 458084 85436 458086
rect 85500 458084 85547 458088
rect 81893 458083 81959 458084
rect 82813 458083 82879 458084
rect 84193 458083 84259 458084
rect 85481 458083 85547 458084
rect 86309 458148 86375 458149
rect 87873 458148 87939 458149
rect 86309 458144 86356 458148
rect 86420 458146 86426 458148
rect 87822 458146 87828 458148
rect 86309 458088 86314 458144
rect 86309 458084 86356 458088
rect 86420 458086 86466 458146
rect 87782 458086 87828 458146
rect 87892 458144 87939 458148
rect 87934 458088 87939 458144
rect 86420 458084 86426 458086
rect 87822 458084 87828 458086
rect 87892 458084 87939 458088
rect 88926 458084 88932 458148
rect 88996 458146 89002 458148
rect 89069 458146 89135 458149
rect 88996 458144 89135 458146
rect 88996 458088 89074 458144
rect 89130 458088 89135 458144
rect 88996 458086 89135 458088
rect 88996 458084 89002 458086
rect 86309 458083 86375 458084
rect 87873 458083 87939 458084
rect 89069 458083 89135 458086
rect 90173 458148 90239 458149
rect 90173 458144 90220 458148
rect 90284 458146 90290 458148
rect 91093 458146 91159 458149
rect 92473 458148 92539 458149
rect 93577 458148 93643 458149
rect 91318 458146 91324 458148
rect 90173 458088 90178 458144
rect 90173 458084 90220 458088
rect 90284 458086 90330 458146
rect 91093 458144 91324 458146
rect 91093 458088 91098 458144
rect 91154 458088 91324 458144
rect 91093 458086 91324 458088
rect 90284 458084 90290 458086
rect 90173 458083 90239 458084
rect 91093 458083 91159 458086
rect 91318 458084 91324 458086
rect 91388 458084 91394 458148
rect 92422 458146 92428 458148
rect 92382 458086 92428 458146
rect 92492 458144 92539 458148
rect 92534 458088 92539 458144
rect 92422 458084 92428 458086
rect 92492 458084 92539 458088
rect 93526 458084 93532 458148
rect 93596 458146 93643 458148
rect 94773 458148 94839 458149
rect 95785 458148 95851 458149
rect 93596 458144 93688 458146
rect 93638 458088 93688 458144
rect 93596 458086 93688 458088
rect 94773 458144 94820 458148
rect 94884 458146 94890 458148
rect 95734 458146 95740 458148
rect 94773 458088 94778 458144
rect 93596 458084 93643 458086
rect 92473 458083 92539 458084
rect 93577 458083 93643 458084
rect 94773 458084 94820 458088
rect 94884 458086 94930 458146
rect 95694 458086 95740 458146
rect 95804 458144 95851 458148
rect 95846 458088 95851 458144
rect 94884 458084 94890 458086
rect 95734 458084 95740 458086
rect 95804 458084 95851 458088
rect 94773 458083 94839 458084
rect 95785 458083 95851 458084
rect 97165 458148 97231 458149
rect 97165 458144 97212 458148
rect 97276 458146 97282 458148
rect 97165 458088 97170 458144
rect 97165 458084 97212 458088
rect 97276 458086 97322 458146
rect 97276 458084 97282 458086
rect 98310 458084 98316 458148
rect 98380 458146 98386 458148
rect 98545 458146 98611 458149
rect 99465 458148 99531 458149
rect 99414 458146 99420 458148
rect 98380 458144 98611 458146
rect 98380 458088 98550 458144
rect 98606 458088 98611 458144
rect 98380 458086 98611 458088
rect 99374 458086 99420 458146
rect 99484 458144 99531 458148
rect 99526 458088 99531 458144
rect 98380 458084 98386 458086
rect 97165 458083 97231 458084
rect 98545 458083 98611 458086
rect 99414 458084 99420 458086
rect 99484 458084 99531 458088
rect 100150 458084 100156 458148
rect 100220 458146 100226 458148
rect 100661 458146 100727 458149
rect 101949 458148 102015 458149
rect 102777 458148 102843 458149
rect 101949 458146 101996 458148
rect 100220 458144 100727 458146
rect 100220 458088 100666 458144
rect 100722 458088 100727 458144
rect 100220 458086 100727 458088
rect 101904 458144 101996 458146
rect 101904 458088 101954 458144
rect 101904 458086 101996 458088
rect 100220 458084 100226 458086
rect 99465 458083 99531 458084
rect 100661 458083 100727 458086
rect 101949 458084 101996 458086
rect 102060 458084 102066 458148
rect 102726 458146 102732 458148
rect 102686 458086 102732 458146
rect 102796 458144 102843 458148
rect 102838 458088 102843 458144
rect 102726 458084 102732 458086
rect 102796 458084 102843 458088
rect 103094 458084 103100 458148
rect 103164 458146 103170 458148
rect 103421 458146 103487 458149
rect 104249 458148 104315 458149
rect 104801 458148 104867 458149
rect 105353 458148 105419 458149
rect 104198 458146 104204 458148
rect 103164 458144 103487 458146
rect 103164 458088 103426 458144
rect 103482 458088 103487 458144
rect 103164 458086 103487 458088
rect 104158 458086 104204 458146
rect 104268 458144 104315 458148
rect 104310 458088 104315 458144
rect 103164 458084 103170 458086
rect 101949 458083 102015 458084
rect 102777 458083 102843 458084
rect 103421 458083 103487 458086
rect 104198 458084 104204 458086
rect 104268 458084 104315 458088
rect 104750 458084 104756 458148
rect 104820 458146 104867 458148
rect 105302 458146 105308 458148
rect 104820 458144 104912 458146
rect 104862 458088 104912 458144
rect 104820 458086 104912 458088
rect 105262 458086 105308 458146
rect 105372 458144 105419 458148
rect 105414 458088 105419 458144
rect 104820 458084 104867 458086
rect 105302 458084 105308 458086
rect 105372 458084 105419 458088
rect 105486 458084 105492 458148
rect 105556 458146 105562 458148
rect 106181 458146 106247 458149
rect 105556 458144 106247 458146
rect 105556 458088 106186 458144
rect 106242 458088 106247 458144
rect 105556 458086 106247 458088
rect 105556 458084 105562 458086
rect 104249 458083 104315 458084
rect 104801 458083 104867 458084
rect 105353 458083 105419 458084
rect 106181 458083 106247 458086
rect 107142 458084 107148 458148
rect 107212 458146 107218 458148
rect 107561 458146 107627 458149
rect 108757 458148 108823 458149
rect 108757 458146 108804 458148
rect 107212 458144 107627 458146
rect 107212 458088 107566 458144
rect 107622 458088 107627 458144
rect 107212 458086 107627 458088
rect 108712 458144 108804 458146
rect 108712 458088 108762 458144
rect 108712 458086 108804 458088
rect 107212 458084 107218 458086
rect 107561 458083 107627 458086
rect 108757 458084 108804 458086
rect 108868 458084 108874 458148
rect 108982 458084 108988 458148
rect 109052 458146 109058 458148
rect 110321 458146 110387 458149
rect 193857 458148 193923 458149
rect 193806 458146 193812 458148
rect 109052 458144 110387 458146
rect 109052 458088 110326 458144
rect 110382 458088 110387 458144
rect 109052 458086 110387 458088
rect 193766 458086 193812 458146
rect 193876 458144 193923 458148
rect 200205 458148 200271 458149
rect 210509 458148 210575 458149
rect 200205 458146 200252 458148
rect 193918 458088 193923 458144
rect 109052 458084 109058 458086
rect 108757 458083 108823 458084
rect 110321 458083 110387 458086
rect 193806 458084 193812 458086
rect 193876 458084 193923 458088
rect 200160 458144 200252 458146
rect 200160 458088 200210 458144
rect 200160 458086 200252 458088
rect 193857 458083 193923 458084
rect 200205 458084 200252 458086
rect 200316 458084 200322 458148
rect 210509 458144 210556 458148
rect 210620 458146 210626 458148
rect 210509 458088 210514 458144
rect 210509 458084 210556 458088
rect 210620 458086 210666 458146
rect 210620 458084 210626 458086
rect 212022 458084 212028 458148
rect 212092 458146 212098 458148
rect 212441 458146 212507 458149
rect 212092 458144 212507 458146
rect 212092 458088 212446 458144
rect 212502 458088 212507 458144
rect 212092 458086 212507 458088
rect 212092 458084 212098 458086
rect 200205 458083 200271 458084
rect 210509 458083 210575 458084
rect 212441 458083 212507 458086
rect 213085 458148 213151 458149
rect 214005 458148 214071 458149
rect 215293 458148 215359 458149
rect 216673 458148 216739 458149
rect 217593 458148 217659 458149
rect 218881 458148 218947 458149
rect 220169 458148 220235 458149
rect 213085 458144 213132 458148
rect 213196 458146 213202 458148
rect 213085 458088 213090 458144
rect 213085 458084 213132 458088
rect 213196 458086 213242 458146
rect 214005 458144 214052 458148
rect 214116 458146 214122 458148
rect 214005 458088 214010 458144
rect 213196 458084 213202 458086
rect 214005 458084 214052 458088
rect 214116 458086 214162 458146
rect 215293 458144 215340 458148
rect 215404 458146 215410 458148
rect 216622 458146 216628 458148
rect 215293 458088 215298 458144
rect 214116 458084 214122 458086
rect 215293 458084 215340 458088
rect 215404 458086 215450 458146
rect 216582 458086 216628 458146
rect 216692 458144 216739 458148
rect 217542 458146 217548 458148
rect 216734 458088 216739 458144
rect 215404 458084 215410 458086
rect 216622 458084 216628 458086
rect 216692 458084 216739 458088
rect 217502 458086 217548 458146
rect 217612 458144 217659 458148
rect 218830 458146 218836 458148
rect 217654 458088 217659 458144
rect 217542 458084 217548 458086
rect 217612 458084 217659 458088
rect 218790 458086 218836 458146
rect 218900 458144 218947 458148
rect 220118 458146 220124 458148
rect 218942 458088 218947 458144
rect 218830 458084 218836 458086
rect 218900 458084 218947 458088
rect 220078 458086 220124 458146
rect 220188 458144 220235 458148
rect 220230 458088 220235 458144
rect 220118 458084 220124 458086
rect 220188 458084 220235 458088
rect 213085 458083 213151 458084
rect 214005 458083 214071 458084
rect 215293 458083 215359 458084
rect 216673 458083 216739 458084
rect 217593 458083 217659 458084
rect 218881 458083 218947 458084
rect 220169 458083 220235 458084
rect 221365 458148 221431 458149
rect 222561 458148 222627 458149
rect 223665 458148 223731 458149
rect 221365 458144 221412 458148
rect 221476 458146 221482 458148
rect 222510 458146 222516 458148
rect 221365 458088 221370 458144
rect 221365 458084 221412 458088
rect 221476 458086 221522 458146
rect 222470 458086 222516 458146
rect 222580 458144 222627 458148
rect 223614 458146 223620 458148
rect 222622 458088 222627 458144
rect 221476 458084 221482 458086
rect 222510 458084 222516 458086
rect 222580 458084 222627 458088
rect 223574 458086 223620 458146
rect 223684 458144 223731 458148
rect 223726 458088 223731 458144
rect 223614 458084 223620 458086
rect 223684 458084 223731 458088
rect 221365 458083 221431 458084
rect 222561 458083 222627 458084
rect 223665 458083 223731 458084
rect 224309 458148 224375 458149
rect 225873 458148 225939 458149
rect 227161 458148 227227 458149
rect 224309 458144 224356 458148
rect 224420 458146 224426 458148
rect 225822 458146 225828 458148
rect 224309 458088 224314 458144
rect 224309 458084 224356 458088
rect 224420 458086 224466 458146
rect 225782 458086 225828 458146
rect 225892 458144 225939 458148
rect 227110 458146 227116 458148
rect 225934 458088 225939 458144
rect 224420 458084 224426 458086
rect 225822 458084 225828 458086
rect 225892 458084 225939 458088
rect 227070 458086 227116 458146
rect 227180 458144 227227 458148
rect 227222 458088 227227 458144
rect 227110 458084 227116 458086
rect 227180 458084 227227 458088
rect 224309 458083 224375 458084
rect 225873 458083 225939 458084
rect 227161 458083 227227 458084
rect 228357 458148 228423 458149
rect 229553 458148 229619 458149
rect 228357 458144 228404 458148
rect 228468 458146 228474 458148
rect 229502 458146 229508 458148
rect 228357 458088 228362 458144
rect 228357 458084 228404 458088
rect 228468 458086 228514 458146
rect 229462 458086 229508 458146
rect 229572 458144 229619 458148
rect 229614 458088 229619 458144
rect 228468 458084 228474 458086
rect 229502 458084 229508 458086
rect 229572 458084 229619 458088
rect 228357 458083 228423 458084
rect 229553 458083 229619 458084
rect 231853 458146 231919 458149
rect 232814 458146 232820 458148
rect 231853 458144 232820 458146
rect 231853 458088 231858 458144
rect 231914 458088 232820 458144
rect 231853 458086 232820 458088
rect 231853 458083 231919 458086
rect 232814 458084 232820 458086
rect 232884 458084 232890 458148
rect 233233 458146 233299 458149
rect 313733 458148 313799 458149
rect 233550 458146 233556 458148
rect 233233 458144 233556 458146
rect 233233 458088 233238 458144
rect 233294 458088 233556 458144
rect 233233 458086 233556 458088
rect 233233 458083 233299 458086
rect 233550 458084 233556 458086
rect 233620 458084 233626 458148
rect 313733 458144 313780 458148
rect 313844 458146 313850 458148
rect 321553 458146 321619 458149
rect 322790 458146 322796 458148
rect 313733 458088 313738 458144
rect 313733 458084 313780 458088
rect 313844 458086 313890 458146
rect 321553 458144 322796 458146
rect 321553 458088 321558 458144
rect 321614 458088 322796 458144
rect 321553 458086 322796 458088
rect 313844 458084 313850 458086
rect 313733 458083 313799 458084
rect 321553 458083 321619 458086
rect 322790 458084 322796 458086
rect 322860 458084 322866 458148
rect 322933 458146 322999 458149
rect 323894 458146 323900 458148
rect 322933 458144 323900 458146
rect 322933 458088 322938 458144
rect 322994 458088 323900 458144
rect 322933 458086 323900 458088
rect 322933 458083 322999 458086
rect 323894 458084 323900 458086
rect 323964 458084 323970 458148
rect 325693 458146 325759 458149
rect 326286 458146 326292 458148
rect 325693 458144 326292 458146
rect 325693 458088 325698 458144
rect 325754 458088 326292 458144
rect 325693 458086 326292 458088
rect 325693 458083 325759 458086
rect 326286 458084 326292 458086
rect 326356 458084 326362 458148
rect 327073 458146 327139 458149
rect 327390 458146 327396 458148
rect 327073 458144 327396 458146
rect 327073 458088 327078 458144
rect 327134 458088 327396 458144
rect 327073 458086 327396 458088
rect 327073 458083 327139 458086
rect 327390 458084 327396 458086
rect 327460 458084 327466 458148
rect 328862 458084 328868 458148
rect 328932 458146 328938 458148
rect 329097 458146 329163 458149
rect 328932 458144 329163 458146
rect 328932 458088 329102 458144
rect 329158 458088 329163 458144
rect 328932 458086 329163 458088
rect 328932 458084 328938 458086
rect 329097 458083 329163 458086
rect 329925 458146 329991 458149
rect 331857 458148 331923 458149
rect 333145 458148 333211 458149
rect 334065 458148 334131 458149
rect 335353 458148 335419 458149
rect 330886 458146 330892 458148
rect 329925 458144 330892 458146
rect 329925 458088 329930 458144
rect 329986 458088 330892 458144
rect 329925 458086 330892 458088
rect 329925 458083 329991 458086
rect 330886 458084 330892 458086
rect 330956 458084 330962 458148
rect 331806 458146 331812 458148
rect 331766 458086 331812 458146
rect 331876 458144 331923 458148
rect 333094 458146 333100 458148
rect 331918 458088 331923 458144
rect 331806 458084 331812 458086
rect 331876 458084 331923 458088
rect 333054 458086 333100 458146
rect 333164 458144 333211 458148
rect 334014 458146 334020 458148
rect 333206 458088 333211 458144
rect 333094 458084 333100 458086
rect 333164 458084 333211 458088
rect 333974 458086 334020 458146
rect 334084 458144 334131 458148
rect 334126 458088 334131 458144
rect 334014 458084 334020 458086
rect 334084 458084 334131 458088
rect 335302 458084 335308 458148
rect 335372 458146 335419 458148
rect 336549 458148 336615 458149
rect 335372 458144 335464 458146
rect 335414 458088 335464 458144
rect 335372 458086 335464 458088
rect 336549 458144 336596 458148
rect 336660 458146 336666 458148
rect 336549 458088 336554 458144
rect 335372 458084 335419 458086
rect 331857 458083 331923 458084
rect 333145 458083 333211 458084
rect 334065 458083 334131 458084
rect 335353 458083 335419 458084
rect 336549 458084 336596 458088
rect 336660 458086 336706 458146
rect 336660 458084 336666 458086
rect 337694 458084 337700 458148
rect 337764 458146 337770 458148
rect 338021 458146 338087 458149
rect 339033 458148 339099 458149
rect 338982 458146 338988 458148
rect 337764 458144 338087 458146
rect 337764 458088 338026 458144
rect 338082 458088 338087 458144
rect 337764 458086 338087 458088
rect 338942 458086 338988 458146
rect 339052 458144 339099 458148
rect 339094 458088 339099 458144
rect 337764 458084 337770 458086
rect 336549 458083 336615 458084
rect 338021 458083 338087 458086
rect 338982 458084 338988 458086
rect 339052 458084 339099 458088
rect 339033 458083 339099 458084
rect 339861 458148 339927 458149
rect 341241 458148 341307 458149
rect 339861 458144 339908 458148
rect 339972 458146 339978 458148
rect 341190 458146 341196 458148
rect 339861 458088 339866 458144
rect 339861 458084 339908 458088
rect 339972 458086 340018 458146
rect 341150 458086 341196 458146
rect 341260 458144 341307 458148
rect 341302 458088 341307 458144
rect 339972 458084 339978 458086
rect 341190 458084 341196 458086
rect 341260 458084 341307 458088
rect 339861 458083 339927 458084
rect 341241 458083 341307 458084
rect 342253 458146 342319 458149
rect 342662 458146 342668 458148
rect 342253 458144 342668 458146
rect 342253 458088 342258 458144
rect 342314 458088 342668 458144
rect 342253 458086 342668 458088
rect 342253 458083 342319 458086
rect 342662 458084 342668 458086
rect 342732 458084 342738 458148
rect 343633 458146 343699 458149
rect 344737 458148 344803 458149
rect 343950 458146 343956 458148
rect 343633 458144 343956 458146
rect 343633 458088 343638 458144
rect 343694 458088 343956 458144
rect 343633 458086 343956 458088
rect 343633 458083 343699 458086
rect 343950 458084 343956 458086
rect 344020 458084 344026 458148
rect 344686 458146 344692 458148
rect 344646 458086 344692 458146
rect 344756 458144 344803 458148
rect 344798 458088 344803 458144
rect 344686 458084 344692 458086
rect 344756 458084 344803 458088
rect 344737 458083 344803 458084
rect 345013 458146 345079 458149
rect 346158 458146 346164 458148
rect 345013 458144 346164 458146
rect 345013 458088 345018 458144
rect 345074 458088 346164 458144
rect 345013 458086 346164 458088
rect 345013 458083 345079 458086
rect 346158 458084 346164 458086
rect 346228 458084 346234 458148
rect 346393 458146 346459 458149
rect 347262 458146 347268 458148
rect 346393 458144 347268 458146
rect 346393 458088 346398 458144
rect 346454 458088 347268 458144
rect 346393 458086 347268 458088
rect 346393 458083 346459 458086
rect 347262 458084 347268 458086
rect 347332 458084 347338 458148
rect 347773 458146 347839 458149
rect 348366 458146 348372 458148
rect 347773 458144 348372 458146
rect 347773 458088 347778 458144
rect 347834 458088 348372 458144
rect 347773 458086 348372 458088
rect 347773 458083 347839 458086
rect 348366 458084 348372 458086
rect 348436 458084 348442 458148
rect 349153 458146 349219 458149
rect 349654 458146 349660 458148
rect 349153 458144 349660 458146
rect 349153 458088 349158 458144
rect 349214 458088 349660 458144
rect 349153 458086 349660 458088
rect 349153 458083 349219 458086
rect 349654 458084 349660 458086
rect 349724 458084 349730 458148
rect 351913 458146 351979 458149
rect 352966 458146 352972 458148
rect 351913 458144 352972 458146
rect 351913 458088 351918 458144
rect 351974 458088 352972 458144
rect 351913 458086 352972 458088
rect 351913 458083 351979 458086
rect 352966 458084 352972 458086
rect 353036 458084 353042 458148
rect 353293 458146 353359 458149
rect 461761 458148 461827 458149
rect 463049 458148 463115 458149
rect 353518 458146 353524 458148
rect 353293 458144 353524 458146
rect 353293 458088 353298 458144
rect 353354 458088 353524 458144
rect 353293 458086 353524 458088
rect 353293 458083 353359 458086
rect 353518 458084 353524 458086
rect 353588 458084 353594 458148
rect 461710 458146 461716 458148
rect 461670 458086 461716 458146
rect 461780 458144 461827 458148
rect 462998 458146 463004 458148
rect 461822 458088 461827 458144
rect 461710 458084 461716 458086
rect 461780 458084 461827 458088
rect 462958 458086 463004 458146
rect 463068 458144 463115 458148
rect 463110 458088 463115 458144
rect 462998 458084 463004 458086
rect 463068 458084 463115 458088
rect 464286 458084 464292 458148
rect 464356 458146 464362 458148
rect 464981 458146 465047 458149
rect 464356 458144 465047 458146
rect 464356 458088 464986 458144
rect 465042 458088 465047 458144
rect 464356 458086 465047 458088
rect 464356 458084 464362 458086
rect 461761 458083 461827 458084
rect 463049 458083 463115 458084
rect 464981 458083 465047 458086
rect 465165 458148 465231 458149
rect 468753 458148 468819 458149
rect 465165 458144 465212 458148
rect 465276 458146 465282 458148
rect 468702 458146 468708 458148
rect 465165 458088 465170 458144
rect 465165 458084 465212 458088
rect 465276 458086 465322 458146
rect 468662 458086 468708 458146
rect 468772 458144 468819 458148
rect 468814 458088 468819 458144
rect 465276 458084 465282 458086
rect 468702 458084 468708 458086
rect 468772 458084 468819 458088
rect 465165 458083 465231 458084
rect 468753 458083 468819 458084
rect 469949 458148 470015 458149
rect 469949 458144 469996 458148
rect 470060 458146 470066 458148
rect 469949 458088 469954 458144
rect 469949 458084 469996 458088
rect 470060 458086 470106 458146
rect 470060 458084 470066 458086
rect 471278 458084 471284 458148
rect 471348 458146 471354 458148
rect 471789 458146 471855 458149
rect 472249 458148 472315 458149
rect 472198 458146 472204 458148
rect 471348 458144 471855 458146
rect 471348 458088 471794 458144
rect 471850 458088 471855 458144
rect 471348 458086 471855 458088
rect 472158 458086 472204 458146
rect 472268 458144 472315 458148
rect 472310 458088 472315 458144
rect 471348 458084 471354 458086
rect 469949 458083 470015 458084
rect 471789 458083 471855 458086
rect 472198 458084 472204 458086
rect 472268 458084 472315 458088
rect 472249 458083 472315 458084
rect 473445 458148 473511 458149
rect 474825 458148 474891 458149
rect 473445 458144 473492 458148
rect 473556 458146 473562 458148
rect 474774 458146 474780 458148
rect 473445 458088 473450 458144
rect 473445 458084 473492 458088
rect 473556 458086 473602 458146
rect 474734 458086 474780 458146
rect 474844 458144 474891 458148
rect 474886 458088 474891 458144
rect 473556 458084 473562 458086
rect 474774 458084 474780 458086
rect 474844 458084 474891 458088
rect 473445 458083 473511 458084
rect 474825 458083 474891 458084
rect 475469 458148 475535 458149
rect 476941 458148 477007 458149
rect 478321 458148 478387 458149
rect 479425 458148 479491 458149
rect 475469 458144 475516 458148
rect 475580 458146 475586 458148
rect 475469 458088 475474 458144
rect 475469 458084 475516 458088
rect 475580 458086 475626 458146
rect 476941 458144 476988 458148
rect 477052 458146 477058 458148
rect 478270 458146 478276 458148
rect 476941 458088 476946 458144
rect 475580 458084 475586 458086
rect 476941 458084 476988 458088
rect 477052 458086 477098 458146
rect 478230 458086 478276 458146
rect 478340 458144 478387 458148
rect 479374 458146 479380 458148
rect 478382 458088 478387 458144
rect 477052 458084 477058 458086
rect 478270 458084 478276 458086
rect 478340 458084 478387 458088
rect 479334 458086 479380 458146
rect 479444 458144 479491 458148
rect 483013 458148 483079 458149
rect 483013 458146 483060 458148
rect 479486 458088 479491 458144
rect 479374 458084 479380 458086
rect 479444 458084 479491 458088
rect 482968 458144 483060 458146
rect 482968 458088 483018 458144
rect 482968 458086 483060 458088
rect 475469 458083 475535 458084
rect 476941 458083 477007 458084
rect 478321 458083 478387 458084
rect 479425 458083 479491 458084
rect 483013 458084 483060 458086
rect 483124 458084 483130 458148
rect 483197 458146 483263 458149
rect 484158 458146 484164 458148
rect 483197 458144 484164 458146
rect 483197 458088 483202 458144
rect 483258 458088 484164 458144
rect 483197 458086 484164 458088
rect 483013 458083 483079 458084
rect 483197 458083 483263 458086
rect 484158 458084 484164 458086
rect 484228 458084 484234 458148
rect 484393 458146 484459 458149
rect 485446 458146 485452 458148
rect 484393 458144 485452 458146
rect 484393 458088 484398 458144
rect 484454 458088 485452 458144
rect 484393 458086 485452 458088
rect 484393 458083 484459 458086
rect 485446 458084 485452 458086
rect 485516 458084 485522 458148
rect 80646 457948 80652 458012
rect 80716 458010 80722 458012
rect 81341 458010 81407 458013
rect 100569 458012 100635 458013
rect 100518 458010 100524 458012
rect 80716 458008 81407 458010
rect 80716 457952 81346 458008
rect 81402 457952 81407 458008
rect 80716 457950 81407 457952
rect 100478 457950 100524 458010
rect 100588 458008 100635 458012
rect 100630 457952 100635 458008
rect 80716 457948 80722 457950
rect 81341 457947 81407 457950
rect 100518 457948 100524 457950
rect 100588 457948 100635 457952
rect 101438 457948 101444 458012
rect 101508 458010 101514 458012
rect 102041 458010 102107 458013
rect 101508 458008 102107 458010
rect 101508 457952 102046 458008
rect 102102 457952 102107 458008
rect 101508 457950 102107 457952
rect 101508 457948 101514 457950
rect 100569 457947 100635 457948
rect 102041 457947 102107 457950
rect 106273 458010 106339 458013
rect 107653 458012 107719 458013
rect 106406 458010 106412 458012
rect 106273 458008 106412 458010
rect 106273 457952 106278 458008
rect 106334 457952 106412 458008
rect 106273 457950 106412 457952
rect 106273 457947 106339 457950
rect 106406 457948 106412 457950
rect 106476 457948 106482 458012
rect 107653 458008 107700 458012
rect 107764 458010 107770 458012
rect 107653 457952 107658 458008
rect 107653 457948 107700 457952
rect 107764 457950 107810 458010
rect 107764 457948 107770 457950
rect 108430 457948 108436 458012
rect 108500 458010 108506 458012
rect 108941 458010 109007 458013
rect 108500 458008 109007 458010
rect 108500 457952 108946 458008
rect 109002 457952 109007 458008
rect 108500 457950 109007 457952
rect 108500 457948 108506 457950
rect 107653 457947 107719 457948
rect 108941 457947 109007 457950
rect 197353 458010 197419 458013
rect 197486 458010 197492 458012
rect 197353 458008 197492 458010
rect 197353 457952 197358 458008
rect 197414 457952 197492 458008
rect 197353 457950 197492 457952
rect 197353 457947 197419 457950
rect 197486 457948 197492 457950
rect 197556 457948 197562 458012
rect 198733 458010 198799 458013
rect 199142 458010 199148 458012
rect 198733 458008 199148 458010
rect 198733 457952 198738 458008
rect 198794 457952 199148 458008
rect 198733 457950 199148 457952
rect 198733 457947 198799 457950
rect 199142 457948 199148 457950
rect 199212 457948 199218 458012
rect 207054 457948 207060 458012
rect 207124 458010 207130 458012
rect 207657 458010 207723 458013
rect 208209 458010 208275 458013
rect 234613 458012 234679 458013
rect 234613 458010 234660 458012
rect 207124 458008 208275 458010
rect 207124 457952 207662 458008
rect 207718 457952 208214 458008
rect 208270 457952 208275 458008
rect 207124 457950 208275 457952
rect 234568 458008 234660 458010
rect 234568 457952 234618 458008
rect 234568 457950 234660 457952
rect 207124 457948 207130 457950
rect 207657 457947 207723 457950
rect 208209 457947 208275 457950
rect 234613 457948 234660 457950
rect 234724 457948 234730 458012
rect 322197 458010 322263 458013
rect 323577 458012 323643 458013
rect 322606 458010 322612 458012
rect 322197 458008 322612 458010
rect 322197 457952 322202 458008
rect 322258 457952 322612 458008
rect 322197 457950 322612 457952
rect 234613 457947 234679 457948
rect 322197 457947 322263 457950
rect 322606 457948 322612 457950
rect 322676 457948 322682 458012
rect 323526 458010 323532 458012
rect 323486 457950 323532 458010
rect 323596 458008 323643 458012
rect 323638 457952 323643 458008
rect 323526 457948 323532 457950
rect 323596 457948 323643 457952
rect 323577 457947 323643 457948
rect 329281 458010 329347 458013
rect 342529 458012 342595 458013
rect 329598 458010 329604 458012
rect 329281 458008 329604 458010
rect 329281 457952 329286 458008
rect 329342 457952 329604 458008
rect 329281 457950 329604 457952
rect 329281 457947 329347 457950
rect 329598 457948 329604 457950
rect 329668 457948 329674 458012
rect 342478 458010 342484 458012
rect 342438 457950 342484 458010
rect 342548 458008 342595 458012
rect 342590 457952 342595 458008
rect 342478 457948 342484 457950
rect 342548 457948 342595 457952
rect 343582 457948 343588 458012
rect 343652 458010 343658 458012
rect 344369 458010 344435 458013
rect 343652 458008 344435 458010
rect 343652 457952 344374 458008
rect 344430 457952 344435 458008
rect 343652 457950 344435 457952
rect 343652 457948 343658 457950
rect 342529 457947 342595 457948
rect 344369 457947 344435 457950
rect 345933 458012 345999 458013
rect 346853 458012 346919 458013
rect 348233 458012 348299 458013
rect 345933 458008 345980 458012
rect 346044 458010 346050 458012
rect 345933 457952 345938 458008
rect 345933 457948 345980 457952
rect 346044 457950 346090 458010
rect 346853 458008 346900 458012
rect 346964 458010 346970 458012
rect 348182 458010 348188 458012
rect 346853 457952 346858 458008
rect 346044 457948 346050 457950
rect 346853 457948 346900 457952
rect 346964 457950 347010 458010
rect 348142 457950 348188 458010
rect 348252 458008 348299 458012
rect 348294 457952 348299 458008
rect 346964 457948 346970 457950
rect 348182 457948 348188 457950
rect 348252 457948 348299 457952
rect 345933 457947 345999 457948
rect 346853 457947 346919 457948
rect 348233 457947 348299 457948
rect 349245 458010 349311 458013
rect 350533 458012 350599 458013
rect 349470 458010 349476 458012
rect 349245 458008 349476 458010
rect 349245 457952 349250 458008
rect 349306 457952 349476 458008
rect 349245 457950 349476 457952
rect 349245 457947 349311 457950
rect 349470 457948 349476 457950
rect 349540 457948 349546 458012
rect 350533 458010 350580 458012
rect 350488 458008 350580 458010
rect 350488 457952 350538 458008
rect 350488 457950 350580 457952
rect 350533 457948 350580 457950
rect 350644 457948 350650 458012
rect 356053 458010 356119 458013
rect 356462 458010 356468 458012
rect 356053 458008 356468 458010
rect 356053 457952 356058 458008
rect 356114 457952 356468 458008
rect 356053 457950 356468 457952
rect 350533 457947 350599 457948
rect 356053 457947 356119 457950
rect 356462 457948 356468 457950
rect 356532 457948 356538 458012
rect 442993 458010 443059 458013
rect 443126 458010 443132 458012
rect 442993 458008 443132 458010
rect 442993 457952 442998 458008
rect 443054 457952 443132 458008
rect 442993 457950 443132 457952
rect 442993 457947 443059 457950
rect 443126 457948 443132 457950
rect 443196 457948 443202 458012
rect 459502 457948 459508 458012
rect 459572 458010 459578 458012
rect 460197 458010 460263 458013
rect 459572 458008 460263 458010
rect 459572 457952 460202 458008
rect 460258 457952 460263 458008
rect 459572 457950 460263 457952
rect 459572 457948 459578 457950
rect 460197 457947 460263 457950
rect 467782 457948 467788 458012
rect 467852 458010 467858 458012
rect 468017 458010 468083 458013
rect 467852 458008 468083 458010
rect 467852 457952 468022 458008
rect 468078 457952 468083 458008
rect 467852 457950 468083 457952
rect 467852 457948 467858 457950
rect 468017 457947 468083 457950
rect 480437 458010 480503 458013
rect 480662 458010 480668 458012
rect 480437 458008 480668 458010
rect 480437 457952 480442 458008
rect 480498 457952 480668 458008
rect 480437 457950 480668 457952
rect 480437 457947 480503 457950
rect 480662 457948 480668 457950
rect 480732 457948 480738 458012
rect 487153 458010 487219 458013
rect 487654 458010 487660 458012
rect 487153 458008 487660 458010
rect 487153 457952 487158 458008
rect 487214 457952 487660 458008
rect 487153 457950 487660 457952
rect 487153 457947 487219 457950
rect 487654 457948 487660 457950
rect 487724 457948 487730 458012
rect 78438 457812 78444 457876
rect 78508 457874 78514 457876
rect 78581 457874 78647 457877
rect 101857 457876 101923 457877
rect 101806 457874 101812 457876
rect 78508 457872 78647 457874
rect 78508 457816 78586 457872
rect 78642 457816 78647 457872
rect 78508 457814 78647 457816
rect 101766 457814 101812 457874
rect 101876 457872 101923 457876
rect 231853 457876 231919 457877
rect 231853 457874 231900 457876
rect 101918 457816 101923 457872
rect 78508 457812 78514 457814
rect 78581 457811 78647 457814
rect 101806 457812 101812 457814
rect 101876 457812 101923 457816
rect 231808 457872 231900 457874
rect 231808 457816 231858 457872
rect 231808 457814 231900 457816
rect 101857 457811 101923 457812
rect 231853 457812 231900 457814
rect 231964 457812 231970 457876
rect 235993 457874 236059 457877
rect 317413 457876 317479 457877
rect 236494 457874 236500 457876
rect 235993 457872 236500 457874
rect 235993 457816 235998 457872
rect 236054 457816 236500 457872
rect 235993 457814 236500 457816
rect 231853 457811 231919 457812
rect 235993 457811 236059 457814
rect 236494 457812 236500 457814
rect 236564 457812 236570 457876
rect 317413 457874 317460 457876
rect 317368 457872 317460 457874
rect 317368 457816 317418 457872
rect 317368 457814 317460 457816
rect 317413 457812 317460 457814
rect 317524 457812 317530 457876
rect 324814 457812 324820 457876
rect 324884 457874 324890 457876
rect 324957 457874 325023 457877
rect 324884 457872 325023 457874
rect 324884 457816 324962 457872
rect 325018 457816 325023 457872
rect 324884 457814 325023 457816
rect 324884 457812 324890 457814
rect 317413 457811 317479 457812
rect 324957 457811 325023 457814
rect 326102 457812 326108 457876
rect 326172 457874 326178 457876
rect 326337 457874 326403 457877
rect 330477 457876 330543 457877
rect 330477 457874 330524 457876
rect 326172 457872 326403 457874
rect 326172 457816 326342 457872
rect 326398 457816 326403 457872
rect 326172 457814 326403 457816
rect 330432 457872 330524 457874
rect 330432 457816 330482 457872
rect 330432 457814 330524 457816
rect 326172 457812 326178 457814
rect 326337 457811 326403 457814
rect 330477 457812 330524 457814
rect 330588 457812 330594 457876
rect 355041 457874 355107 457877
rect 355174 457874 355180 457876
rect 355041 457872 355180 457874
rect 355041 457816 355046 457872
rect 355102 457816 355180 457872
rect 355041 457814 355180 457816
rect 330477 457811 330543 457812
rect 355041 457811 355107 457814
rect 355174 457812 355180 457814
rect 355244 457812 355250 457876
rect 458173 457874 458239 457877
rect 458582 457874 458588 457876
rect 458173 457872 458588 457874
rect 458173 457816 458178 457872
rect 458234 457816 458588 457872
rect 458173 457814 458588 457816
rect 458173 457811 458239 457814
rect 458582 457812 458588 457814
rect 458652 457812 458658 457876
rect 466494 457812 466500 457876
rect 466564 457874 466570 457876
rect 466637 457874 466703 457877
rect 466564 457872 466703 457874
rect 466564 457816 466642 457872
rect 466698 457816 466703 457872
rect 466564 457814 466703 457816
rect 466564 457812 466570 457814
rect 466637 457811 466703 457814
rect 478873 457874 478939 457877
rect 479558 457874 479564 457876
rect 478873 457872 479564 457874
rect 478873 457816 478878 457872
rect 478934 457816 479564 457872
rect 478873 457814 479564 457816
rect 478873 457811 478939 457814
rect 479558 457812 479564 457814
rect 479628 457812 479634 457876
rect 480529 457874 480595 457877
rect 480846 457874 480852 457876
rect 480529 457872 480852 457874
rect 480529 457816 480534 457872
rect 480590 457816 480852 457872
rect 480529 457814 480852 457816
rect 480529 457811 480595 457814
rect 480846 457812 480852 457814
rect 480916 457812 480922 457876
rect 484393 457874 484459 457877
rect 484710 457874 484716 457876
rect 484393 457872 484716 457874
rect 484393 457816 484398 457872
rect 484454 457816 484716 457872
rect 484393 457814 484716 457816
rect 484393 457811 484459 457814
rect 484710 457812 484716 457814
rect 484780 457812 484786 457876
rect 72734 457676 72740 457740
rect 72804 457738 72810 457740
rect 73061 457738 73127 457741
rect 201493 457740 201559 457741
rect 209681 457740 209747 457741
rect 201493 457738 201540 457740
rect 72804 457736 73127 457738
rect 72804 457680 73066 457736
rect 73122 457680 73127 457736
rect 72804 457678 73127 457680
rect 201448 457736 201540 457738
rect 201448 457680 201498 457736
rect 201448 457678 201540 457680
rect 72804 457676 72810 457678
rect 73061 457675 73127 457678
rect 201493 457676 201540 457678
rect 201604 457676 201610 457740
rect 209630 457738 209636 457740
rect 209590 457678 209636 457738
rect 209700 457736 209747 457740
rect 237373 457740 237439 457741
rect 237373 457738 237420 457740
rect 209742 457680 209747 457736
rect 209630 457676 209636 457678
rect 209700 457676 209747 457680
rect 237328 457736 237420 457738
rect 237328 457680 237378 457736
rect 237328 457678 237420 457680
rect 201493 457675 201559 457676
rect 209681 457675 209747 457676
rect 237373 457676 237420 457678
rect 237484 457676 237490 457740
rect 238753 457738 238819 457741
rect 238886 457738 238892 457740
rect 238753 457736 238892 457738
rect 238753 457680 238758 457736
rect 238814 457680 238892 457736
rect 238753 457678 238892 457680
rect 237373 457675 237439 457676
rect 238753 457675 238819 457678
rect 238886 457676 238892 457678
rect 238956 457676 238962 457740
rect 331213 457738 331279 457741
rect 331990 457738 331996 457740
rect 331213 457736 331996 457738
rect 331213 457680 331218 457736
rect 331274 457680 331996 457736
rect 331213 457678 331996 457680
rect 331213 457675 331279 457678
rect 331990 457676 331996 457678
rect 332060 457676 332066 457740
rect 343725 457738 343791 457741
rect 357433 457740 357499 457741
rect 344870 457738 344876 457740
rect 343725 457736 344876 457738
rect 343725 457680 343730 457736
rect 343786 457680 344876 457736
rect 343725 457678 344876 457680
rect 343725 457675 343791 457678
rect 344870 457676 344876 457678
rect 344940 457676 344946 457740
rect 357382 457676 357388 457740
rect 357452 457738 357499 457740
rect 460381 457738 460447 457741
rect 481633 457740 481699 457741
rect 460790 457738 460796 457740
rect 357452 457736 357544 457738
rect 357494 457680 357544 457736
rect 357452 457678 357544 457680
rect 460381 457736 460796 457738
rect 460381 457680 460386 457736
rect 460442 457680 460796 457736
rect 460381 457678 460796 457680
rect 357452 457676 357499 457678
rect 357433 457675 357499 457676
rect 460381 457675 460447 457678
rect 460790 457676 460796 457678
rect 460860 457676 460866 457740
rect 481582 457676 481588 457740
rect 481652 457738 481699 457740
rect 485773 457738 485839 457741
rect 488533 457740 488599 457741
rect 485998 457738 486004 457740
rect 481652 457736 481744 457738
rect 481694 457680 481744 457736
rect 481652 457678 481744 457680
rect 485773 457736 486004 457738
rect 485773 457680 485778 457736
rect 485834 457680 486004 457736
rect 485773 457678 486004 457680
rect 481652 457676 481699 457678
rect 481633 457675 481699 457676
rect 485773 457675 485839 457678
rect 485998 457676 486004 457678
rect 486068 457676 486074 457740
rect 488533 457738 488580 457740
rect 488488 457736 488580 457738
rect 488488 457680 488538 457736
rect 488488 457678 488580 457680
rect 488533 457676 488580 457678
rect 488644 457676 488650 457740
rect 488533 457675 488599 457676
rect 63677 457604 63743 457605
rect 63677 457600 63724 457604
rect 63788 457602 63794 457604
rect 63677 457544 63682 457600
rect 63677 457540 63724 457544
rect 63788 457542 63834 457602
rect 63788 457540 63794 457542
rect 75862 457540 75868 457604
rect 75932 457602 75938 457604
rect 77201 457602 77267 457605
rect 75932 457600 77267 457602
rect 75932 457544 77206 457600
rect 77262 457544 77267 457600
rect 75932 457542 77267 457544
rect 75932 457540 75938 457542
rect 63677 457539 63743 457540
rect 77201 457539 77267 457542
rect 195973 457602 196039 457605
rect 196750 457602 196756 457604
rect 195973 457600 196756 457602
rect 195973 457544 195978 457600
rect 196034 457544 196756 457600
rect 195973 457542 196756 457544
rect 195973 457539 196039 457542
rect 196750 457540 196756 457542
rect 196820 457540 196826 457604
rect 230473 457602 230539 457605
rect 230606 457602 230612 457604
rect 230473 457600 230612 457602
rect 230473 457544 230478 457600
rect 230534 457544 230612 457600
rect 230473 457542 230612 457544
rect 230473 457539 230539 457542
rect 230606 457540 230612 457542
rect 230676 457540 230682 457604
rect 456793 457602 456859 457605
rect 457478 457602 457484 457604
rect 456793 457600 457484 457602
rect 456793 457544 456798 457600
rect 456854 457544 457484 457600
rect 456793 457542 457484 457544
rect 456793 457539 456859 457542
rect 457478 457540 457484 457542
rect 457548 457540 457554 457604
rect 459553 457602 459619 457605
rect 459686 457602 459692 457604
rect 459553 457600 459692 457602
rect 459553 457544 459558 457600
rect 459614 457544 459692 457600
rect 459553 457542 459692 457544
rect 459553 457539 459619 457542
rect 459686 457540 459692 457542
rect 459756 457540 459762 457604
rect 487153 457602 487219 457605
rect 487838 457602 487844 457604
rect 487153 457600 487844 457602
rect 487153 457544 487158 457600
rect 487214 457544 487844 457600
rect 487153 457542 487844 457544
rect 487153 457539 487219 457542
rect 487838 457540 487844 457542
rect 487908 457540 487914 457604
rect 73153 457466 73219 457469
rect 74206 457466 74212 457468
rect 73153 457464 74212 457466
rect 73153 457408 73158 457464
rect 73214 457408 74212 457464
rect 73153 457406 74212 457408
rect 73153 457403 73219 457406
rect 74206 457404 74212 457406
rect 74276 457404 74282 457468
rect 75913 457466 75979 457469
rect 76230 457466 76236 457468
rect 75913 457464 76236 457466
rect 75913 457408 75918 457464
rect 75974 457408 76236 457464
rect 75913 457406 76236 457408
rect 75913 457403 75979 457406
rect 76230 457404 76236 457406
rect 76300 457404 76306 457468
rect 208526 457404 208532 457468
rect 208596 457466 208602 457468
rect 209037 457466 209103 457469
rect 208596 457464 209103 457466
rect 208596 457408 209042 457464
rect 209098 457408 209103 457464
rect 208596 457406 209103 457408
rect 208596 457404 208602 457406
rect 209037 457403 209103 457406
rect 216254 457404 216260 457468
rect 216324 457466 216330 457468
rect 216581 457466 216647 457469
rect 216324 457464 216647 457466
rect 216324 457408 216586 457464
rect 216642 457408 216647 457464
rect 216324 457406 216647 457408
rect 216324 457404 216330 457406
rect 216581 457403 216647 457406
rect 452653 457466 452719 457469
rect 453798 457466 453804 457468
rect 452653 457464 453804 457466
rect 452653 457408 452658 457464
rect 452714 457408 453804 457464
rect 452653 457406 453804 457408
rect 452653 457403 452719 457406
rect 453798 457404 453804 457406
rect 453868 457404 453874 457468
rect 454033 457466 454099 457469
rect 455086 457466 455092 457468
rect 454033 457464 455092 457466
rect 454033 457408 454038 457464
rect 454094 457408 455092 457464
rect 454033 457406 455092 457408
rect 454033 457403 454099 457406
rect 455086 457404 455092 457406
rect 455156 457404 455162 457468
rect 483013 457466 483079 457469
rect 483606 457466 483612 457468
rect 483013 457464 483612 457466
rect 483013 457408 483018 457464
rect 483074 457408 483612 457464
rect 483013 457406 483612 457408
rect 483013 457403 483079 457406
rect 483606 457404 483612 457406
rect 483676 457404 483682 457468
rect 485773 457466 485839 457469
rect 486550 457466 486556 457468
rect 485773 457464 486556 457466
rect 485773 457408 485778 457464
rect 485834 457408 486556 457464
rect 485773 457406 486556 457408
rect 485773 457403 485839 457406
rect 486550 457404 486556 457406
rect 486620 457404 486626 457468
rect 488533 457466 488599 457469
rect 488942 457466 488948 457468
rect 488533 457464 488948 457466
rect 488533 457408 488538 457464
rect 488594 457408 488948 457464
rect 488533 457406 488948 457408
rect 488533 457403 488599 457406
rect 488942 457404 488948 457406
rect 489012 457404 489018 457468
rect 206134 457268 206140 457332
rect 206204 457330 206210 457332
rect 206277 457330 206343 457333
rect 206829 457330 206895 457333
rect 329833 457332 329899 457333
rect 206204 457328 206895 457330
rect 206204 457272 206282 457328
rect 206338 457272 206834 457328
rect 206890 457272 206895 457328
rect 206204 457270 206895 457272
rect 206204 457268 206210 457270
rect 206277 457267 206343 457270
rect 206829 457267 206895 457270
rect 329782 457268 329788 457332
rect 329852 457330 329899 457332
rect 476113 457330 476179 457333
rect 477166 457330 477172 457332
rect 329852 457328 329944 457330
rect 329894 457272 329944 457328
rect 329852 457270 329944 457272
rect 476113 457328 477172 457330
rect 476113 457272 476118 457328
rect 476174 457272 477172 457328
rect 476113 457270 477172 457272
rect 329852 457268 329899 457270
rect 329833 457267 329899 457268
rect 476113 457267 476179 457270
rect 477166 457268 477172 457270
rect 477236 457268 477242 457332
rect 477493 457330 477559 457333
rect 478454 457330 478460 457332
rect 477493 457328 478460 457330
rect 477493 457272 477498 457328
rect 477554 457272 478460 457328
rect 477493 457270 478460 457272
rect 477493 457267 477559 457270
rect 478454 457268 478460 457270
rect 478524 457268 478530 457332
rect 71773 457194 71839 457197
rect 77293 457196 77359 457197
rect 72918 457194 72924 457196
rect 71773 457192 72924 457194
rect 71773 457136 71778 457192
rect 71834 457136 72924 457192
rect 71773 457134 72924 457136
rect 71773 457131 71839 457134
rect 72918 457132 72924 457134
rect 72988 457132 72994 457196
rect 77293 457194 77340 457196
rect 77248 457192 77340 457194
rect 77248 457136 77298 457192
rect 77248 457134 77340 457136
rect 77293 457132 77340 457134
rect 77404 457132 77410 457196
rect 94998 457132 95004 457196
rect 95068 457194 95074 457196
rect 95141 457194 95207 457197
rect 95068 457192 95207 457194
rect 95068 457136 95146 457192
rect 95202 457136 95207 457192
rect 95068 457134 95207 457136
rect 95068 457132 95074 457134
rect 77293 457131 77359 457132
rect 95141 457131 95207 457134
rect 98494 457132 98500 457196
rect 98564 457194 98570 457196
rect 99281 457194 99347 457197
rect 98564 457192 99347 457194
rect 98564 457136 99286 457192
rect 99342 457136 99347 457192
rect 98564 457134 99347 457136
rect 98564 457132 98570 457134
rect 99281 457131 99347 457134
rect 202137 457194 202203 457197
rect 202454 457194 202460 457196
rect 202137 457192 202460 457194
rect 202137 457136 202142 457192
rect 202198 457136 202460 457192
rect 202137 457134 202460 457136
rect 202137 457131 202203 457134
rect 202454 457132 202460 457134
rect 202524 457132 202530 457196
rect 202638 457132 202644 457196
rect 202708 457194 202714 457196
rect 202781 457194 202847 457197
rect 202708 457192 202847 457194
rect 202708 457136 202786 457192
rect 202842 457136 202847 457192
rect 202708 457134 202847 457136
rect 202708 457132 202714 457134
rect 202781 457131 202847 457134
rect 206318 457132 206324 457196
rect 206388 457194 206394 457196
rect 206921 457194 206987 457197
rect 206388 457192 206987 457194
rect 206388 457136 206926 457192
rect 206982 457136 206987 457192
rect 206388 457134 206987 457136
rect 206388 457132 206394 457134
rect 206921 457131 206987 457134
rect 209814 457132 209820 457196
rect 209884 457194 209890 457196
rect 210969 457194 211035 457197
rect 209884 457192 211035 457194
rect 209884 457136 210974 457192
rect 211030 457136 211035 457192
rect 209884 457134 211035 457136
rect 209884 457132 209890 457134
rect 210969 457131 211035 457134
rect 214414 457132 214420 457196
rect 214484 457194 214490 457196
rect 215201 457194 215267 457197
rect 214484 457192 215267 457194
rect 214484 457136 215206 457192
rect 215262 457136 215267 457192
rect 214484 457134 215267 457136
rect 214484 457132 214490 457134
rect 215201 457131 215267 457134
rect 216806 457132 216812 457196
rect 216876 457194 216882 457196
rect 217961 457194 218027 457197
rect 216876 457192 218027 457194
rect 216876 457136 217966 457192
rect 218022 457136 218027 457192
rect 216876 457134 218027 457136
rect 216876 457132 216882 457134
rect 217961 457131 218027 457134
rect 220302 457132 220308 457196
rect 220372 457194 220378 457196
rect 220721 457194 220787 457197
rect 220372 457192 220787 457194
rect 220372 457136 220726 457192
rect 220782 457136 220787 457192
rect 220372 457134 220787 457136
rect 220372 457132 220378 457134
rect 220721 457131 220787 457134
rect 324313 457194 324379 457197
rect 328453 457196 328519 457197
rect 324998 457194 325004 457196
rect 324313 457192 325004 457194
rect 324313 457136 324318 457192
rect 324374 457136 325004 457192
rect 324313 457134 325004 457136
rect 324313 457131 324379 457134
rect 324998 457132 325004 457134
rect 325068 457132 325074 457196
rect 328453 457194 328500 457196
rect 328408 457192 328500 457194
rect 328408 457136 328458 457192
rect 328408 457134 328500 457136
rect 328453 457132 328500 457134
rect 328564 457132 328570 457196
rect 335353 457194 335419 457197
rect 335486 457194 335492 457196
rect 335353 457192 335492 457194
rect 335353 457136 335358 457192
rect 335414 457136 335492 457192
rect 335353 457134 335492 457136
rect 328453 457131 328519 457132
rect 335353 457131 335419 457134
rect 335486 457132 335492 457134
rect 335556 457132 335562 457196
rect 340873 457194 340939 457197
rect 341374 457194 341380 457196
rect 340873 457192 341380 457194
rect 340873 457136 340878 457192
rect 340934 457136 341380 457192
rect 340873 457134 341380 457136
rect 340873 457131 340939 457134
rect 341374 457132 341380 457134
rect 341444 457132 341450 457196
rect 353293 457194 353359 457197
rect 354254 457194 354260 457196
rect 353293 457192 354260 457194
rect 353293 457136 353298 457192
rect 353354 457136 354260 457192
rect 353293 457134 354260 457136
rect 353293 457131 353359 457134
rect 354254 457132 354260 457134
rect 354324 457132 354330 457196
rect 450537 457194 450603 457197
rect 454677 457196 454743 457197
rect 451406 457194 451412 457196
rect 450537 457192 451412 457194
rect 450537 457136 450542 457192
rect 450598 457136 451412 457192
rect 450537 457134 451412 457136
rect 450537 457131 450603 457134
rect 451406 457132 451412 457134
rect 451476 457132 451482 457196
rect 454677 457192 454724 457196
rect 454788 457194 454794 457196
rect 454677 457136 454682 457192
rect 454677 457132 454724 457136
rect 454788 457134 454834 457194
rect 454788 457132 454794 457134
rect 458214 457132 458220 457196
rect 458284 457194 458290 457196
rect 458817 457194 458883 457197
rect 459369 457194 459435 457197
rect 458284 457192 459435 457194
rect 458284 457136 458822 457192
rect 458878 457136 459374 457192
rect 459430 457136 459435 457192
rect 458284 457134 459435 457136
rect 458284 457132 458290 457134
rect 454677 457131 454743 457132
rect 458817 457131 458883 457134
rect 459369 457131 459435 457134
rect 461025 457194 461091 457197
rect 462078 457194 462084 457196
rect 461025 457192 462084 457194
rect 461025 457136 461030 457192
rect 461086 457136 462084 457192
rect 461025 457134 462084 457136
rect 461025 457131 461091 457134
rect 462078 457132 462084 457134
rect 462148 457132 462154 457196
rect 467925 457194 467991 457197
rect 469070 457194 469076 457196
rect 467925 457192 469076 457194
rect 467925 457136 467930 457192
rect 467986 457136 469076 457192
rect 467925 457134 469076 457136
rect 467925 457131 467991 457134
rect 469070 457132 469076 457134
rect 469140 457132 469146 457196
rect 471973 457194 472039 457197
rect 472566 457194 472572 457196
rect 471973 457192 472572 457194
rect 471973 457136 471978 457192
rect 472034 457136 472572 457192
rect 471973 457134 472572 457136
rect 471973 457131 472039 457134
rect 472566 457132 472572 457134
rect 472636 457132 472642 457196
rect 476062 457132 476068 457196
rect 476132 457194 476138 457196
rect 476205 457194 476271 457197
rect 476132 457192 476271 457194
rect 476132 457136 476210 457192
rect 476266 457136 476271 457192
rect 476132 457134 476271 457136
rect 476132 457132 476138 457134
rect 476205 457131 476271 457134
rect 481633 457194 481699 457197
rect 481950 457194 481956 457196
rect 481633 457192 481956 457194
rect 481633 457136 481638 457192
rect 481694 457136 481956 457192
rect 481633 457134 481956 457136
rect 481633 457131 481699 457134
rect 481950 457132 481956 457134
rect 482020 457132 482026 457196
rect 70209 457060 70275 457061
rect 70158 456996 70164 457060
rect 70228 457058 70275 457060
rect 74717 457058 74783 457061
rect 75126 457058 75132 457060
rect 70228 457056 70320 457058
rect 70270 457000 70320 457056
rect 70228 456998 70320 457000
rect 74717 457056 75132 457058
rect 74717 457000 74722 457056
rect 74778 457000 75132 457056
rect 74717 456998 75132 457000
rect 70228 456996 70275 456998
rect 70209 456995 70275 456996
rect 74717 456995 74783 456998
rect 75126 456996 75132 456998
rect 75196 456996 75202 457060
rect 78622 456996 78628 457060
rect 78692 457058 78698 457060
rect 78765 457058 78831 457061
rect 78692 457056 78831 457058
rect 78692 457000 78770 457056
rect 78826 457000 78831 457056
rect 78692 456998 78831 457000
rect 78692 456996 78698 456998
rect 78765 456995 78831 456998
rect 93158 456996 93164 457060
rect 93228 457058 93234 457060
rect 93761 457058 93827 457061
rect 93228 457056 93827 457058
rect 93228 457000 93766 457056
rect 93822 457000 93827 457056
rect 93228 456998 93827 457000
rect 93228 456996 93234 456998
rect 93761 456995 93827 456998
rect 204897 457058 204963 457061
rect 205030 457058 205036 457060
rect 204897 457056 205036 457058
rect 204897 457000 204902 457056
rect 204958 457000 205036 457056
rect 204897 456998 205036 457000
rect 204897 456995 204963 456998
rect 205030 456996 205036 456998
rect 205100 457058 205106 457060
rect 205449 457058 205515 457061
rect 205100 457056 205515 457058
rect 205100 457000 205454 457056
rect 205510 457000 205515 457056
rect 205100 456998 205515 457000
rect 205100 456996 205106 456998
rect 205449 456995 205515 456998
rect 225638 456996 225644 457060
rect 225708 457058 225714 457060
rect 226241 457058 226307 457061
rect 225708 457056 226307 457058
rect 225708 457000 226246 457056
rect 226302 457000 226307 457056
rect 225708 456998 226307 457000
rect 225708 456996 225714 456998
rect 226241 456995 226307 456998
rect 232630 456996 232636 457060
rect 232700 457058 232706 457060
rect 233049 457058 233115 457061
rect 232700 457056 233115 457058
rect 232700 457000 233054 457056
rect 233110 457000 233115 457056
rect 232700 456998 233115 457000
rect 232700 456996 232706 456998
rect 233049 456995 233115 456998
rect 320265 457058 320331 457061
rect 320950 457058 320956 457060
rect 320265 457056 320956 457058
rect 320265 457000 320270 457056
rect 320326 457000 320956 457056
rect 320265 456998 320956 457000
rect 320265 456995 320331 456998
rect 320950 456996 320956 456998
rect 321020 456996 321026 457060
rect 336825 457058 336891 457061
rect 337878 457058 337884 457060
rect 336825 457056 337884 457058
rect 336825 457000 336830 457056
rect 336886 457000 337884 457056
rect 336825 456998 337884 457000
rect 336825 456995 336891 456998
rect 337878 456996 337884 456998
rect 337948 456996 337954 457060
rect 352005 457058 352071 457061
rect 353150 457058 353156 457060
rect 352005 457056 353156 457058
rect 352005 457000 352010 457056
rect 352066 457000 353156 457056
rect 352005 456998 353156 457000
rect 352005 456995 352071 456998
rect 353150 456996 353156 456998
rect 353220 456996 353226 457060
rect 446397 457058 446463 457061
rect 456057 457060 456123 457061
rect 447910 457058 447916 457060
rect 446397 457056 447916 457058
rect 446397 457000 446402 457056
rect 446458 457000 447916 457056
rect 446397 456998 447916 457000
rect 446397 456995 446463 456998
rect 447910 456996 447916 456998
rect 447980 456996 447986 457060
rect 456006 457058 456012 457060
rect 455930 456998 456012 457058
rect 456076 457058 456123 457060
rect 456701 457058 456767 457061
rect 456076 457056 456767 457058
rect 456118 457000 456706 457056
rect 456762 457000 456767 457056
rect 456006 456996 456012 456998
rect 456076 456998 456767 457000
rect 456076 456996 456123 456998
rect 456057 456995 456123 456996
rect 456701 456995 456767 456998
rect 66846 456860 66852 456924
rect 66916 456922 66922 456924
rect 67541 456922 67607 456925
rect 66916 456920 67607 456922
rect 66916 456864 67546 456920
rect 67602 456864 67607 456920
rect 66916 456862 67607 456864
rect 66916 456860 66922 456862
rect 67541 456859 67607 456862
rect 67950 456860 67956 456924
rect 68020 456922 68026 456924
rect 68829 456922 68895 456925
rect 68020 456920 68895 456922
rect 68020 456864 68834 456920
rect 68890 456864 68895 456920
rect 68020 456862 68895 456864
rect 68020 456860 68026 456862
rect 68829 456859 68895 456862
rect 69790 456860 69796 456924
rect 69860 456922 69866 456924
rect 70117 456922 70183 456925
rect 69860 456920 70183 456922
rect 69860 456864 70122 456920
rect 70178 456864 70183 456920
rect 69860 456862 70183 456864
rect 69860 456860 69866 456862
rect 70117 456859 70183 456862
rect 71446 456860 71452 456924
rect 71516 456922 71522 456924
rect 71681 456922 71747 456925
rect 71516 456920 71747 456922
rect 71516 456864 71686 456920
rect 71742 456864 71747 456920
rect 71516 456862 71747 456864
rect 71516 456860 71522 456862
rect 71681 456859 71747 456862
rect 78673 456922 78739 456925
rect 79726 456922 79732 456924
rect 78673 456920 79732 456922
rect 78673 456864 78678 456920
rect 78734 456864 79732 456920
rect 78673 456862 79732 456864
rect 78673 456859 78739 456862
rect 79726 456860 79732 456862
rect 79796 456860 79802 456924
rect 80053 456922 80119 456925
rect 80830 456922 80836 456924
rect 80053 456920 80836 456922
rect 80053 456864 80058 456920
rect 80114 456864 80836 456920
rect 80053 456862 80836 456864
rect 80053 456859 80119 456862
rect 80830 456860 80836 456862
rect 80900 456860 80906 456924
rect 81433 456922 81499 456925
rect 82118 456922 82124 456924
rect 81433 456920 82124 456922
rect 81433 456864 81438 456920
rect 81494 456864 82124 456920
rect 81433 456862 82124 456864
rect 81433 456859 81499 456862
rect 82118 456860 82124 456862
rect 82188 456860 82194 456924
rect 82813 456922 82879 456925
rect 83222 456922 83228 456924
rect 82813 456920 83228 456922
rect 82813 456864 82818 456920
rect 82874 456864 83228 456920
rect 82813 456862 83228 456864
rect 82813 456859 82879 456862
rect 83222 456860 83228 456862
rect 83292 456860 83298 456924
rect 84193 456922 84259 456925
rect 84326 456922 84332 456924
rect 84193 456920 84332 456922
rect 84193 456864 84198 456920
rect 84254 456864 84332 456920
rect 84193 456862 84332 456864
rect 84193 456859 84259 456862
rect 84326 456860 84332 456862
rect 84396 456860 84402 456924
rect 85614 456860 85620 456924
rect 85684 456922 85690 456924
rect 86217 456922 86283 456925
rect 85684 456920 86283 456922
rect 85684 456864 86222 456920
rect 86278 456864 86283 456920
rect 85684 456862 86283 456864
rect 85684 456860 85690 456862
rect 86217 456859 86283 456862
rect 86718 456860 86724 456924
rect 86788 456922 86794 456924
rect 86861 456922 86927 456925
rect 86788 456920 86927 456922
rect 86788 456864 86866 456920
rect 86922 456864 86927 456920
rect 86788 456862 86927 456864
rect 86788 456860 86794 456862
rect 86861 456859 86927 456862
rect 88006 456860 88012 456924
rect 88076 456922 88082 456924
rect 88241 456922 88307 456925
rect 88076 456920 88307 456922
rect 88076 456864 88246 456920
rect 88302 456864 88307 456920
rect 88076 456862 88307 456864
rect 88076 456860 88082 456862
rect 88241 456859 88307 456862
rect 89110 456860 89116 456924
rect 89180 456922 89186 456924
rect 89621 456922 89687 456925
rect 89180 456920 89687 456922
rect 89180 456864 89626 456920
rect 89682 456864 89687 456920
rect 89180 456862 89687 456864
rect 89180 456860 89186 456862
rect 89621 456859 89687 456862
rect 90582 456860 90588 456924
rect 90652 456922 90658 456924
rect 91001 456922 91067 456925
rect 90652 456920 91067 456922
rect 90652 456864 91006 456920
rect 91062 456864 91067 456920
rect 90652 456862 91067 456864
rect 90652 456860 90658 456862
rect 91001 456859 91067 456862
rect 91502 456860 91508 456924
rect 91572 456922 91578 456924
rect 92381 456922 92447 456925
rect 93669 456924 93735 456925
rect 93669 456922 93716 456924
rect 91572 456920 92447 456922
rect 91572 456864 92386 456920
rect 92442 456864 92447 456920
rect 91572 456862 92447 456864
rect 93624 456920 93716 456922
rect 93624 456864 93674 456920
rect 93624 456862 93716 456864
rect 91572 456860 91578 456862
rect 92381 456859 92447 456862
rect 93669 456860 93716 456862
rect 93780 456860 93786 456924
rect 96102 456860 96108 456924
rect 96172 456922 96178 456924
rect 96521 456922 96587 456925
rect 96172 456920 96587 456922
rect 96172 456864 96526 456920
rect 96582 456864 96587 456920
rect 96172 456862 96587 456864
rect 96172 456860 96178 456862
rect 93669 456859 93735 456860
rect 96521 456859 96587 456862
rect 97758 456860 97764 456924
rect 97828 456922 97834 456924
rect 97901 456922 97967 456925
rect 97828 456920 97967 456922
rect 97828 456864 97906 456920
rect 97962 456864 97967 456920
rect 97828 456862 97967 456864
rect 97828 456860 97834 456862
rect 97901 456859 97967 456862
rect 203517 456922 203583 456925
rect 203742 456922 203748 456924
rect 203517 456920 203748 456922
rect 203517 456864 203522 456920
rect 203578 456864 203748 456920
rect 203517 456862 203748 456864
rect 203517 456859 203583 456862
rect 203742 456860 203748 456862
rect 203812 456860 203818 456924
rect 203926 456860 203932 456924
rect 203996 456922 204002 456924
rect 204161 456922 204227 456925
rect 203996 456920 204227 456922
rect 203996 456864 204166 456920
rect 204222 456864 204227 456920
rect 203996 456862 204227 456864
rect 203996 456860 204002 456862
rect 204161 456859 204227 456862
rect 205398 456860 205404 456924
rect 205468 456922 205474 456924
rect 205541 456922 205607 456925
rect 205468 456920 205607 456922
rect 205468 456864 205546 456920
rect 205602 456864 205607 456920
rect 205468 456862 205607 456864
rect 205468 456860 205474 456862
rect 205541 456859 205607 456862
rect 207422 456860 207428 456924
rect 207492 456922 207498 456924
rect 208301 456922 208367 456925
rect 207492 456920 208367 456922
rect 207492 456864 208306 456920
rect 208362 456864 208367 456920
rect 207492 456862 208367 456864
rect 207492 456860 207498 456862
rect 208301 456859 208367 456862
rect 209262 456860 209268 456924
rect 209332 456922 209338 456924
rect 209681 456922 209747 456925
rect 209332 456920 209747 456922
rect 209332 456864 209686 456920
rect 209742 456864 209747 456920
rect 209332 456862 209747 456864
rect 209332 456860 209338 456862
rect 209681 456859 209747 456862
rect 210918 456860 210924 456924
rect 210988 456922 210994 456924
rect 211061 456922 211127 456925
rect 212441 456924 212507 456925
rect 210988 456920 211127 456922
rect 210988 456864 211066 456920
rect 211122 456864 211127 456920
rect 210988 456862 211127 456864
rect 210988 456860 210994 456862
rect 211061 456859 211127 456862
rect 212390 456860 212396 456924
rect 212460 456922 212507 456924
rect 212460 456920 212552 456922
rect 212502 456864 212552 456920
rect 212460 456862 212552 456864
rect 212460 456860 212507 456862
rect 213310 456860 213316 456924
rect 213380 456922 213386 456924
rect 213821 456922 213887 456925
rect 217869 456924 217935 456925
rect 217869 456922 217916 456924
rect 213380 456920 213887 456922
rect 213380 456864 213826 456920
rect 213882 456864 213887 456920
rect 213380 456862 213887 456864
rect 217824 456920 217916 456922
rect 217824 456864 217874 456920
rect 217824 456862 217916 456864
rect 213380 456860 213386 456862
rect 212441 456859 212507 456860
rect 213821 456859 213887 456862
rect 217869 456860 217916 456862
rect 217980 456860 217986 456924
rect 219198 456860 219204 456924
rect 219268 456922 219274 456924
rect 219341 456922 219407 456925
rect 219268 456920 219407 456922
rect 219268 456864 219346 456920
rect 219402 456864 219407 456920
rect 219268 456862 219407 456864
rect 219268 456860 219274 456862
rect 217869 456859 217935 456860
rect 219341 456859 219407 456862
rect 221958 456860 221964 456924
rect 222028 456922 222034 456924
rect 222101 456922 222167 456925
rect 222028 456920 222167 456922
rect 222028 456864 222106 456920
rect 222162 456864 222167 456920
rect 222028 456862 222167 456864
rect 222028 456860 222034 456862
rect 222101 456859 222167 456862
rect 223246 456860 223252 456924
rect 223316 456922 223322 456924
rect 223481 456922 223547 456925
rect 223316 456920 223547 456922
rect 223316 456864 223486 456920
rect 223542 456864 223547 456920
rect 223316 456862 223547 456864
rect 223316 456860 223322 456862
rect 223481 456859 223547 456862
rect 223798 456860 223804 456924
rect 223868 456922 223874 456924
rect 224861 456922 224927 456925
rect 226149 456924 226215 456925
rect 226149 456922 226196 456924
rect 223868 456920 224927 456922
rect 223868 456864 224866 456920
rect 224922 456864 224927 456920
rect 223868 456862 224927 456864
rect 226104 456920 226196 456922
rect 226104 456864 226154 456920
rect 226104 456862 226196 456864
rect 223868 456860 223874 456862
rect 224861 456859 224927 456862
rect 226149 456860 226196 456862
rect 226260 456860 226266 456924
rect 227294 456860 227300 456924
rect 227364 456922 227370 456924
rect 227621 456922 227687 456925
rect 229001 456924 229067 456925
rect 228950 456922 228956 456924
rect 227364 456920 227687 456922
rect 227364 456864 227626 456920
rect 227682 456864 227687 456920
rect 227364 456862 227687 456864
rect 228910 456862 228956 456922
rect 229020 456920 229067 456924
rect 229062 456864 229067 456920
rect 227364 456860 227370 456862
rect 226149 456859 226215 456860
rect 227621 456859 227687 456862
rect 228950 456860 228956 456862
rect 229020 456860 229067 456864
rect 229686 456860 229692 456924
rect 229756 456922 229762 456924
rect 230381 456922 230447 456925
rect 229756 456920 230447 456922
rect 229756 456864 230386 456920
rect 230442 456864 230447 456920
rect 229756 456862 230447 456864
rect 229756 456860 229762 456862
rect 229001 456859 229067 456860
rect 230381 456859 230447 456862
rect 230790 456860 230796 456924
rect 230860 456922 230866 456924
rect 231761 456922 231827 456925
rect 230860 456920 231827 456922
rect 230860 456864 231766 456920
rect 231822 456864 231827 456920
rect 230860 456862 231827 456864
rect 230860 456860 230866 456862
rect 231761 456859 231827 456862
rect 232998 456860 233004 456924
rect 233068 456922 233074 456924
rect 233141 456922 233207 456925
rect 233068 456920 233207 456922
rect 233068 456864 233146 456920
rect 233202 456864 233207 456920
rect 233068 456862 233207 456864
rect 233068 456860 233074 456862
rect 233141 456859 233207 456862
rect 234286 456860 234292 456924
rect 234356 456922 234362 456924
rect 234521 456922 234587 456925
rect 234356 456920 234587 456922
rect 234356 456864 234526 456920
rect 234582 456864 234587 456920
rect 234356 456862 234587 456864
rect 234356 456860 234362 456862
rect 234521 456859 234587 456862
rect 235758 456860 235764 456924
rect 235828 456922 235834 456924
rect 235901 456922 235967 456925
rect 235828 456920 235967 456922
rect 235828 456864 235906 456920
rect 235962 456864 235967 456920
rect 235828 456862 235967 456864
rect 235828 456860 235834 456862
rect 235901 456859 235967 456862
rect 236678 456860 236684 456924
rect 236748 456922 236754 456924
rect 237281 456922 237347 456925
rect 236748 456920 237347 456922
rect 236748 456864 237286 456920
rect 237342 456864 237347 456920
rect 236748 456862 237347 456864
rect 236748 456860 236754 456862
rect 237281 456859 237347 456862
rect 237782 456860 237788 456924
rect 237852 456922 237858 456924
rect 238661 456922 238727 456925
rect 237852 456920 238727 456922
rect 237852 456864 238666 456920
rect 238722 456864 238727 456920
rect 237852 456862 238727 456864
rect 237852 456860 237858 456862
rect 238661 456859 238727 456862
rect 239622 456860 239628 456924
rect 239692 456922 239698 456924
rect 240041 456922 240107 456925
rect 239692 456920 240107 456922
rect 239692 456864 240046 456920
rect 240102 456864 240107 456920
rect 239692 456862 240107 456864
rect 239692 456860 239698 456862
rect 240041 456859 240107 456862
rect 316033 456922 316099 456925
rect 316166 456922 316172 456924
rect 316033 456920 316172 456922
rect 316033 456864 316038 456920
rect 316094 456864 316172 456920
rect 316033 456862 316172 456864
rect 316033 456859 316099 456862
rect 316166 456860 316172 456862
rect 316236 456860 316242 456924
rect 318793 456922 318859 456925
rect 320173 456924 320239 456925
rect 319110 456922 319116 456924
rect 318793 456920 319116 456922
rect 318793 456864 318798 456920
rect 318854 456864 319116 456920
rect 318793 456862 319116 456864
rect 318793 456859 318859 456862
rect 319110 456860 319116 456862
rect 319180 456860 319186 456924
rect 320173 456922 320220 456924
rect 320128 456920 320220 456922
rect 320128 456864 320178 456920
rect 320128 456862 320220 456864
rect 320173 456860 320220 456862
rect 320284 456860 320290 456924
rect 332593 456922 332659 456925
rect 333278 456922 333284 456924
rect 332593 456920 333284 456922
rect 332593 456864 332598 456920
rect 332654 456864 333284 456920
rect 332593 456862 333284 456864
rect 320173 456859 320239 456860
rect 332593 456859 332659 456862
rect 333278 456860 333284 456862
rect 333348 456860 333354 456924
rect 333973 456922 334039 456925
rect 336733 456924 336799 456925
rect 334382 456922 334388 456924
rect 333973 456920 334388 456922
rect 333973 456864 333978 456920
rect 334034 456864 334388 456920
rect 333973 456862 334388 456864
rect 333973 456859 334039 456862
rect 334382 456860 334388 456862
rect 334452 456860 334458 456924
rect 336733 456922 336780 456924
rect 336688 456920 336780 456922
rect 336688 456864 336738 456920
rect 336688 456862 336780 456864
rect 336733 456860 336780 456862
rect 336844 456860 336850 456924
rect 338113 456922 338179 456925
rect 339166 456922 339172 456924
rect 338113 456920 339172 456922
rect 338113 456864 338118 456920
rect 338174 456864 339172 456920
rect 338113 456862 339172 456864
rect 336733 456859 336799 456860
rect 338113 456859 338179 456862
rect 339166 456860 339172 456862
rect 339236 456860 339242 456924
rect 339493 456922 339559 456925
rect 340270 456922 340276 456924
rect 339493 456920 340276 456922
rect 339493 456864 339498 456920
rect 339554 456864 340276 456920
rect 339493 456862 340276 456864
rect 339493 456859 339559 456862
rect 340270 456860 340276 456862
rect 340340 456860 340346 456924
rect 350533 456922 350599 456925
rect 351913 456924 351979 456925
rect 350942 456922 350948 456924
rect 350533 456920 350948 456922
rect 350533 456864 350538 456920
rect 350594 456864 350948 456920
rect 350533 456862 350948 456864
rect 350533 456859 350599 456862
rect 350942 456860 350948 456862
rect 351012 456860 351018 456924
rect 351862 456860 351868 456924
rect 351932 456922 351979 456924
rect 354673 456922 354739 456925
rect 355358 456922 355364 456924
rect 351932 456920 352024 456922
rect 351974 456864 352024 456920
rect 351932 456862 352024 456864
rect 354673 456920 355364 456922
rect 354673 456864 354678 456920
rect 354734 456864 355364 456920
rect 354673 456862 355364 456864
rect 351932 456860 351979 456862
rect 351913 456859 351979 456860
rect 354673 456859 354739 456862
rect 355358 456860 355364 456862
rect 355428 456860 355434 456924
rect 356053 456922 356119 456925
rect 356646 456922 356652 456924
rect 356053 456920 356652 456922
rect 356053 456864 356058 456920
rect 356114 456864 356652 456920
rect 356053 456862 356652 456864
rect 356053 456859 356119 456862
rect 356646 456860 356652 456862
rect 356716 456860 356722 456924
rect 357433 456922 357499 456925
rect 358813 456924 358879 456925
rect 357750 456922 357756 456924
rect 357433 456920 357756 456922
rect 357433 456864 357438 456920
rect 357494 456864 357756 456920
rect 357433 456862 357756 456864
rect 357433 456859 357499 456862
rect 357750 456860 357756 456862
rect 357820 456860 357826 456924
rect 358813 456922 358860 456924
rect 358768 456920 358860 456922
rect 358768 456864 358818 456920
rect 358768 456862 358860 456864
rect 358813 456860 358860 456862
rect 358924 456860 358930 456924
rect 445753 456922 445819 456925
rect 446806 456922 446812 456924
rect 445753 456920 446812 456922
rect 445753 456864 445758 456920
rect 445814 456864 446812 456920
rect 445753 456862 446812 456864
rect 358813 456859 358879 456860
rect 445753 456859 445819 456862
rect 446806 456860 446812 456862
rect 446876 456860 446882 456924
rect 447777 456922 447843 456925
rect 448462 456922 448468 456924
rect 447777 456920 448468 456922
rect 447777 456864 447782 456920
rect 447838 456864 448468 456920
rect 447777 456862 448468 456864
rect 447777 456859 447843 456862
rect 448462 456860 448468 456862
rect 448532 456860 448538 456924
rect 449157 456922 449223 456925
rect 452745 456924 452811 456925
rect 450302 456922 450308 456924
rect 449157 456920 450308 456922
rect 449157 456864 449162 456920
rect 449218 456864 450308 456920
rect 449157 456862 450308 456864
rect 449157 456859 449223 456862
rect 450302 456860 450308 456862
rect 450372 456860 450378 456924
rect 452694 456860 452700 456924
rect 452764 456922 452811 456924
rect 452764 456920 452856 456922
rect 452806 456864 452856 456920
rect 452764 456862 452856 456864
rect 452764 456860 452811 456862
rect 453062 456860 453068 456924
rect 453132 456922 453138 456924
rect 453297 456922 453363 456925
rect 453132 456920 453363 456922
rect 453132 456864 453302 456920
rect 453358 456864 453363 456920
rect 453132 456862 453363 456864
rect 453132 456860 453138 456862
rect 452745 456859 452811 456860
rect 453297 456859 453363 456862
rect 453481 456922 453547 456925
rect 453614 456922 453620 456924
rect 453481 456920 453620 456922
rect 453481 456864 453486 456920
rect 453542 456864 453620 456920
rect 453481 456862 453620 456864
rect 453481 456859 453547 456862
rect 453614 456860 453620 456862
rect 453684 456860 453690 456924
rect 455413 456922 455479 456925
rect 456190 456922 456196 456924
rect 455413 456920 456196 456922
rect 455413 456864 455418 456920
rect 455474 456864 456196 456920
rect 455413 456862 456196 456864
rect 455413 456859 455479 456862
rect 456190 456860 456196 456862
rect 456260 456860 456266 456924
rect 457294 456860 457300 456924
rect 457364 456922 457370 456924
rect 457437 456922 457503 456925
rect 458081 456922 458147 456925
rect 457364 456920 458147 456922
rect 457364 456864 457442 456920
rect 457498 456864 458086 456920
rect 458142 456864 458147 456920
rect 457364 456862 458147 456864
rect 457364 456860 457370 456862
rect 457437 456859 457503 456862
rect 458081 456859 458147 456862
rect 460933 456924 460999 456925
rect 460933 456920 460980 456924
rect 461044 456922 461050 456924
rect 462313 456922 462379 456925
rect 463182 456922 463188 456924
rect 460933 456864 460938 456920
rect 460933 456860 460980 456864
rect 461044 456862 461090 456922
rect 462313 456920 463188 456922
rect 462313 456864 462318 456920
rect 462374 456864 463188 456920
rect 462313 456862 463188 456864
rect 461044 456860 461050 456862
rect 460933 456859 460999 456860
rect 462313 456859 462379 456862
rect 463182 456860 463188 456862
rect 463252 456860 463258 456924
rect 463693 456922 463759 456925
rect 464470 456922 464476 456924
rect 463693 456920 464476 456922
rect 463693 456864 463698 456920
rect 463754 456864 464476 456920
rect 463693 456862 464476 456864
rect 463693 456859 463759 456862
rect 464470 456860 464476 456862
rect 464540 456860 464546 456924
rect 465073 456922 465139 456925
rect 465574 456922 465580 456924
rect 465073 456920 465580 456922
rect 465073 456864 465078 456920
rect 465134 456864 465580 456920
rect 465073 456862 465580 456864
rect 465073 456859 465139 456862
rect 465574 456860 465580 456862
rect 465644 456860 465650 456924
rect 466453 456922 466519 456925
rect 466678 456922 466684 456924
rect 466453 456920 466684 456922
rect 466453 456864 466458 456920
rect 466514 456864 466684 456920
rect 466453 456862 466684 456864
rect 466453 456859 466519 456862
rect 466678 456860 466684 456862
rect 466748 456860 466754 456924
rect 467833 456922 467899 456925
rect 467966 456922 467972 456924
rect 467833 456920 467972 456922
rect 467833 456864 467838 456920
rect 467894 456864 467972 456920
rect 467833 456862 467972 456864
rect 467833 456859 467899 456862
rect 467966 456860 467972 456862
rect 468036 456860 468042 456924
rect 469213 456922 469279 456925
rect 470174 456922 470180 456924
rect 469213 456920 470180 456922
rect 469213 456864 469218 456920
rect 469274 456864 470180 456920
rect 469213 456862 470180 456864
rect 469213 456859 469279 456862
rect 470174 456860 470180 456862
rect 470244 456860 470250 456924
rect 470593 456922 470659 456925
rect 471462 456922 471468 456924
rect 470593 456920 471468 456922
rect 470593 456864 470598 456920
rect 470654 456864 471468 456920
rect 470593 456862 471468 456864
rect 470593 456859 470659 456862
rect 471462 456860 471468 456862
rect 471532 456860 471538 456924
rect 473353 456922 473419 456925
rect 473670 456922 473676 456924
rect 473353 456920 473676 456922
rect 473353 456864 473358 456920
rect 473414 456864 473676 456920
rect 473353 456862 473676 456864
rect 473353 456859 473419 456862
rect 473670 456860 473676 456862
rect 473740 456860 473746 456924
rect 474733 456922 474799 456925
rect 474958 456922 474964 456924
rect 474733 456920 474964 456922
rect 474733 456864 474738 456920
rect 474794 456864 474964 456920
rect 474733 456862 474964 456864
rect 474733 456859 474799 456862
rect 474958 456860 474964 456862
rect 475028 456860 475034 456924
rect 327717 454066 327783 454069
rect 327901 454066 327967 454069
rect 327717 454064 327967 454066
rect 327717 454008 327722 454064
rect 327778 454008 327906 454064
rect 327962 454008 327967 454064
rect 327717 454006 327967 454008
rect 327717 454003 327783 454006
rect 327901 454003 327967 454006
rect -960 452434 480 452524
rect 3969 452434 4035 452437
rect -960 452432 4035 452434
rect -960 452376 3974 452432
rect 4030 452376 4035 452432
rect -960 452374 4035 452376
rect -960 452284 480 452374
rect 3969 452371 4035 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 56869 442506 56935 442509
rect 162945 442506 163011 442509
rect 56869 442504 163011 442506
rect 56869 442448 56874 442504
rect 56930 442448 162950 442504
rect 163006 442448 163011 442504
rect 56869 442446 163011 442448
rect 56869 442443 56935 442446
rect 162945 442443 163011 442446
rect 233141 442506 233207 442509
rect 287513 442506 287579 442509
rect 233141 442504 287579 442506
rect 233141 442448 233146 442504
rect 233202 442448 287518 442504
rect 287574 442448 287579 442504
rect 233141 442446 287579 442448
rect 233141 442443 233207 442446
rect 287513 442443 287579 442446
rect 57421 442370 57487 442373
rect 165245 442370 165311 442373
rect 57421 442368 165311 442370
rect 57421 442312 57426 442368
rect 57482 442312 165250 442368
rect 165306 442312 165311 442368
rect 57421 442310 165311 442312
rect 57421 442307 57487 442310
rect 165245 442307 165311 442310
rect 234521 442370 234587 442373
rect 289721 442370 289787 442373
rect 234521 442368 289787 442370
rect 234521 442312 234526 442368
rect 234582 442312 289726 442368
rect 289782 442312 289787 442368
rect 234521 442310 289787 442312
rect 234521 442307 234587 442310
rect 289721 442307 289787 442310
rect 57513 442234 57579 442237
rect 167453 442234 167519 442237
rect 57513 442232 167519 442234
rect 57513 442176 57518 442232
rect 57574 442176 167458 442232
rect 167514 442176 167519 442232
rect 57513 442174 167519 442176
rect 57513 442171 57579 442174
rect 167453 442171 167519 442174
rect 237281 442234 237347 442237
rect 294321 442234 294387 442237
rect 237281 442232 294387 442234
rect 237281 442176 237286 442232
rect 237342 442176 294326 442232
rect 294382 442176 294387 442232
rect 237281 442174 294387 442176
rect 237281 442171 237347 442174
rect 294321 442171 294387 442174
rect 240041 441690 240107 441693
rect 248689 441690 248755 441693
rect 240041 441688 248755 441690
rect 240041 441632 240046 441688
rect 240102 441632 248694 441688
rect 248750 441632 248755 441688
rect 240041 441630 248755 441632
rect 240041 441627 240107 441630
rect 248689 441627 248755 441630
rect 580073 439922 580139 439925
rect 583520 439922 584960 440012
rect 580073 439920 584960 439922
rect 580073 439864 580078 439920
rect 580134 439864 584960 439920
rect 580073 439862 584960 439864
rect 580073 439859 580139 439862
rect 583520 439772 584960 439862
rect 56910 439588 56916 439652
rect 56980 439650 56986 439652
rect 559097 439650 559163 439653
rect 56980 439648 559163 439650
rect 56980 439592 559102 439648
rect 559158 439592 559163 439648
rect 56980 439590 559163 439592
rect 56980 439588 56986 439590
rect 559097 439587 559163 439590
rect 57094 439452 57100 439516
rect 57164 439514 57170 439516
rect 580441 439514 580507 439517
rect 57164 439512 580507 439514
rect 57164 439456 580446 439512
rect 580502 439456 580507 439512
rect 57164 439454 580507 439456
rect 57164 439452 57170 439454
rect 580441 439451 580507 439454
rect 58157 439378 58223 439381
rect 58750 439378 58756 439380
rect 58157 439376 58756 439378
rect 58157 439320 58162 439376
rect 58218 439320 58756 439376
rect 58157 439318 58756 439320
rect 58157 439315 58223 439318
rect 58750 439316 58756 439318
rect 58820 439316 58826 439380
rect 56593 438970 56659 438973
rect 302969 438970 303035 438973
rect 56593 438968 60076 438970
rect 56593 438912 56598 438968
rect 56654 438912 60076 438968
rect 56593 438910 60076 438912
rect 299828 438968 303035 438970
rect 299828 438912 302974 438968
rect 303030 438912 303035 438968
rect 299828 438910 303035 438912
rect 56593 438907 56659 438910
rect 302969 438907 303035 438910
rect -960 438018 480 438108
rect 3325 438018 3391 438021
rect -960 438016 3391 438018
rect -960 437960 3330 438016
rect 3386 437960 3391 438016
rect -960 437958 3391 437960
rect -960 437868 480 437958
rect 3325 437955 3391 437958
rect 56593 436114 56659 436117
rect 60046 436114 60106 436900
rect 302785 436794 302851 436797
rect 299828 436792 302851 436794
rect 299828 436736 302790 436792
rect 302846 436736 302851 436792
rect 299828 436734 302851 436736
rect 302785 436731 302851 436734
rect 56593 436112 60106 436114
rect 56593 436056 56598 436112
rect 56654 436056 60106 436112
rect 56593 436054 60106 436056
rect 56593 436051 56659 436054
rect 56685 434754 56751 434757
rect 56685 434752 60076 434754
rect 56685 434696 56690 434752
rect 56746 434696 60076 434752
rect 56685 434694 60076 434696
rect 56685 434691 56751 434694
rect 302785 434618 302851 434621
rect 299828 434616 302851 434618
rect 299828 434560 302790 434616
rect 302846 434560 302851 434616
rect 299828 434558 302851 434560
rect 302785 434555 302851 434558
rect 56685 432034 56751 432037
rect 60046 432034 60106 432684
rect 302785 432442 302851 432445
rect 299828 432440 302851 432442
rect 299828 432384 302790 432440
rect 302846 432384 302851 432440
rect 299828 432382 302851 432384
rect 302785 432379 302851 432382
rect 56685 432032 60106 432034
rect 56685 431976 56690 432032
rect 56746 431976 60106 432032
rect 56685 431974 60106 431976
rect 56685 431971 56751 431974
rect 57145 430538 57211 430541
rect 57145 430536 60076 430538
rect 57145 430480 57150 430536
rect 57206 430480 60076 430536
rect 57145 430478 60076 430480
rect 57145 430475 57211 430478
rect 302785 430266 302851 430269
rect 299828 430264 302851 430266
rect 299828 430208 302790 430264
rect 302846 430208 302851 430264
rect 299828 430206 302851 430208
rect 302785 430203 302851 430206
rect 57145 428498 57211 428501
rect 57145 428496 60076 428498
rect 57145 428440 57150 428496
rect 57206 428440 60076 428496
rect 57145 428438 60076 428440
rect 57145 428435 57211 428438
rect 583520 428076 584960 428316
rect 302785 427954 302851 427957
rect 299828 427952 302851 427954
rect 299828 427896 302790 427952
rect 302846 427896 302851 427952
rect 299828 427894 302851 427896
rect 302785 427891 302851 427894
rect 57145 426322 57211 426325
rect 57145 426320 60076 426322
rect 57145 426264 57150 426320
rect 57206 426264 60076 426320
rect 57145 426262 60076 426264
rect 57145 426259 57211 426262
rect 302785 425778 302851 425781
rect 299828 425776 302851 425778
rect 299828 425720 302790 425776
rect 302846 425720 302851 425776
rect 299828 425718 302851 425720
rect 302785 425715 302851 425718
rect 57145 424282 57211 424285
rect 57145 424280 60076 424282
rect 57145 424224 57150 424280
rect 57206 424224 60076 424280
rect 57145 424222 60076 424224
rect 57145 424219 57211 424222
rect -960 423738 480 423828
rect 3141 423738 3207 423741
rect -960 423736 3207 423738
rect -960 423680 3146 423736
rect 3202 423680 3207 423736
rect -960 423678 3207 423680
rect -960 423588 480 423678
rect 3141 423675 3207 423678
rect 302785 423602 302851 423605
rect 299828 423600 302851 423602
rect 299828 423544 302790 423600
rect 302846 423544 302851 423600
rect 299828 423542 302851 423544
rect 302785 423539 302851 423542
rect 57145 422106 57211 422109
rect 57145 422104 60076 422106
rect 57145 422048 57150 422104
rect 57206 422048 60076 422104
rect 57145 422046 60076 422048
rect 57145 422043 57211 422046
rect 302785 421426 302851 421429
rect 299828 421424 302851 421426
rect 299828 421368 302790 421424
rect 302846 421368 302851 421424
rect 299828 421366 302851 421368
rect 302785 421363 302851 421366
rect 57145 420066 57211 420069
rect 57145 420064 60076 420066
rect 57145 420008 57150 420064
rect 57206 420008 60076 420064
rect 57145 420006 60076 420008
rect 57145 420003 57211 420006
rect 302785 419250 302851 419253
rect 299828 419248 302851 419250
rect 299828 419192 302790 419248
rect 302846 419192 302851 419248
rect 299828 419190 302851 419192
rect 302785 419187 302851 419190
rect 57145 417890 57211 417893
rect 57145 417888 60076 417890
rect 57145 417832 57150 417888
rect 57206 417832 60076 417888
rect 57145 417830 60076 417832
rect 57145 417827 57211 417830
rect 302785 416938 302851 416941
rect 299828 416936 302851 416938
rect 299828 416880 302790 416936
rect 302846 416880 302851 416936
rect 299828 416878 302851 416880
rect 302785 416875 302851 416878
rect 580441 416530 580507 416533
rect 583520 416530 584960 416620
rect 580441 416528 584960 416530
rect 580441 416472 580446 416528
rect 580502 416472 584960 416528
rect 580441 416470 584960 416472
rect 580441 416467 580507 416470
rect 583520 416380 584960 416470
rect 57145 415850 57211 415853
rect 57145 415848 60076 415850
rect 57145 415792 57150 415848
rect 57206 415792 60076 415848
rect 57145 415790 60076 415792
rect 57145 415787 57211 415790
rect 302785 414762 302851 414765
rect 299828 414760 302851 414762
rect 299828 414704 302790 414760
rect 302846 414704 302851 414760
rect 299828 414702 302851 414704
rect 302785 414699 302851 414702
rect 57145 413674 57211 413677
rect 57145 413672 60076 413674
rect 57145 413616 57150 413672
rect 57206 413616 60076 413672
rect 57145 413614 60076 413616
rect 57145 413611 57211 413614
rect 302785 412586 302851 412589
rect 299828 412584 302851 412586
rect 299828 412528 302790 412584
rect 302846 412528 302851 412584
rect 299828 412526 302851 412528
rect 302785 412523 302851 412526
rect 57145 411634 57211 411637
rect 57145 411632 60076 411634
rect 57145 411576 57150 411632
rect 57206 411576 60076 411632
rect 57145 411574 60076 411576
rect 57145 411571 57211 411574
rect 302785 410410 302851 410413
rect 299828 410408 302851 410410
rect 299828 410352 302790 410408
rect 302846 410352 302851 410408
rect 299828 410350 302851 410352
rect 302785 410347 302851 410350
rect 57145 409458 57211 409461
rect 57145 409456 60076 409458
rect -960 409172 480 409412
rect 57145 409400 57150 409456
rect 57206 409400 60076 409456
rect 57145 409398 60076 409400
rect 57145 409395 57211 409398
rect 302785 408234 302851 408237
rect 299828 408232 302851 408234
rect 299828 408176 302790 408232
rect 302846 408176 302851 408232
rect 299828 408174 302851 408176
rect 302785 408171 302851 408174
rect 57145 407418 57211 407421
rect 57145 407416 60076 407418
rect 57145 407360 57150 407416
rect 57206 407360 60076 407416
rect 57145 407358 60076 407360
rect 57145 407355 57211 407358
rect 302785 405922 302851 405925
rect 299828 405920 302851 405922
rect 299828 405864 302790 405920
rect 302846 405864 302851 405920
rect 299828 405862 302851 405864
rect 302785 405859 302851 405862
rect 57145 405242 57211 405245
rect 57145 405240 60076 405242
rect 57145 405184 57150 405240
rect 57206 405184 60076 405240
rect 57145 405182 60076 405184
rect 57145 405179 57211 405182
rect 580349 404834 580415 404837
rect 583520 404834 584960 404924
rect 580349 404832 584960 404834
rect 580349 404776 580354 404832
rect 580410 404776 584960 404832
rect 580349 404774 584960 404776
rect 580349 404771 580415 404774
rect 583520 404684 584960 404774
rect 302693 403746 302759 403749
rect 299828 403744 302759 403746
rect 299828 403688 302698 403744
rect 302754 403688 302759 403744
rect 299828 403686 302759 403688
rect 302693 403683 302759 403686
rect 57145 403202 57211 403205
rect 57145 403200 60076 403202
rect 57145 403144 57150 403200
rect 57206 403144 60076 403200
rect 57145 403142 60076 403144
rect 57145 403139 57211 403142
rect 302785 401570 302851 401573
rect 299828 401568 302851 401570
rect 299828 401512 302790 401568
rect 302846 401512 302851 401568
rect 299828 401510 302851 401512
rect 302785 401507 302851 401510
rect 56685 401026 56751 401029
rect 56685 401024 60076 401026
rect 56685 400968 56690 401024
rect 56746 400968 60076 401024
rect 56685 400966 60076 400968
rect 56685 400963 56751 400966
rect 302785 399394 302851 399397
rect 299828 399392 302851 399394
rect 299828 399336 302790 399392
rect 302846 399336 302851 399392
rect 299828 399334 302851 399336
rect 302785 399331 302851 399334
rect 56685 398986 56751 398989
rect 56685 398984 60076 398986
rect 56685 398928 56690 398984
rect 56746 398928 60076 398984
rect 56685 398926 60076 398928
rect 56685 398923 56751 398926
rect 302785 397218 302851 397221
rect 299828 397216 302851 397218
rect 299828 397160 302790 397216
rect 302846 397160 302851 397216
rect 299828 397158 302851 397160
rect 302785 397155 302851 397158
rect 56685 396810 56751 396813
rect 56685 396808 60076 396810
rect 56685 396752 56690 396808
rect 56746 396752 60076 396808
rect 56685 396750 60076 396752
rect 56685 396747 56751 396750
rect -960 395042 480 395132
rect 2773 395042 2839 395045
rect -960 395040 2839 395042
rect -960 394984 2778 395040
rect 2834 394984 2839 395040
rect -960 394982 2839 394984
rect -960 394892 480 394982
rect 2773 394979 2839 394982
rect 302509 394906 302575 394909
rect 299828 394904 302575 394906
rect 299828 394848 302514 394904
rect 302570 394848 302575 394904
rect 299828 394846 302575 394848
rect 302509 394843 302575 394846
rect 56501 394770 56567 394773
rect 56501 394768 60076 394770
rect 56501 394712 56506 394768
rect 56562 394712 60076 394768
rect 56501 394710 60076 394712
rect 56501 394707 56567 394710
rect 580625 393002 580691 393005
rect 583520 393002 584960 393092
rect 580625 393000 584960 393002
rect 580625 392944 580630 393000
rect 580686 392944 584960 393000
rect 580625 392942 584960 392944
rect 580625 392939 580691 392942
rect 583520 392852 584960 392942
rect 302693 392730 302759 392733
rect 299828 392728 302759 392730
rect 299828 392672 302698 392728
rect 302754 392672 302759 392728
rect 299828 392670 302759 392672
rect 302693 392667 302759 392670
rect 56593 392594 56659 392597
rect 56593 392592 60076 392594
rect 56593 392536 56598 392592
rect 56654 392536 60076 392592
rect 56593 392534 60076 392536
rect 56593 392531 56659 392534
rect 56593 390554 56659 390557
rect 302785 390554 302851 390557
rect 56593 390552 60076 390554
rect 56593 390496 56598 390552
rect 56654 390496 60076 390552
rect 56593 390494 60076 390496
rect 299828 390552 302851 390554
rect 299828 390496 302790 390552
rect 302846 390496 302851 390552
rect 299828 390494 302851 390496
rect 56593 390491 56659 390494
rect 302785 390491 302851 390494
rect 302785 388378 302851 388381
rect 299828 388376 302851 388378
rect 56593 387834 56659 387837
rect 56726 387834 56732 387836
rect 56593 387832 56732 387834
rect 56593 387776 56598 387832
rect 56654 387776 56732 387832
rect 56593 387774 56732 387776
rect 56593 387771 56659 387774
rect 56726 387772 56732 387774
rect 56796 387772 56802 387836
rect 60046 387834 60106 388348
rect 299828 388320 302790 388376
rect 302846 388320 302851 388376
rect 299828 388318 302851 388320
rect 302785 388315 302851 388318
rect 56918 387774 60106 387834
rect 56593 387698 56659 387701
rect 56918 387698 56978 387774
rect 56593 387696 56978 387698
rect 56593 387640 56598 387696
rect 56654 387640 56978 387696
rect 56593 387638 56978 387640
rect 56593 387635 56659 387638
rect 56593 386338 56659 386341
rect 56593 386336 60076 386338
rect 56593 386280 56598 386336
rect 56654 386280 60076 386336
rect 56593 386278 60076 386280
rect 56593 386275 56659 386278
rect 302509 386202 302575 386205
rect 299828 386200 302575 386202
rect 299828 386144 302514 386200
rect 302570 386144 302575 386200
rect 299828 386142 302575 386144
rect 302509 386139 302575 386142
rect 38653 384978 38719 384981
rect 42885 384978 42951 384981
rect 38653 384976 42951 384978
rect 38653 384920 38658 384976
rect 38714 384920 42890 384976
rect 42946 384920 42951 384976
rect 38653 384918 42951 384920
rect 38653 384915 38719 384918
rect 42885 384915 42951 384918
rect 19333 384842 19399 384845
rect 22093 384842 22159 384845
rect 19333 384840 22159 384842
rect 19333 384784 19338 384840
rect 19394 384784 22098 384840
rect 22154 384784 22159 384840
rect 19333 384782 22159 384784
rect 19333 384779 19399 384782
rect 22093 384779 22159 384782
rect 56593 384162 56659 384165
rect 56593 384160 60076 384162
rect 56593 384104 56598 384160
rect 56654 384104 60076 384160
rect 56593 384102 60076 384104
rect 56593 384099 56659 384102
rect 302509 383890 302575 383893
rect 299828 383888 302575 383890
rect 299828 383832 302514 383888
rect 302570 383832 302575 383888
rect 299828 383830 302575 383832
rect 302509 383827 302575 383830
rect 56593 382122 56659 382125
rect 56593 382120 60076 382122
rect 56593 382064 56598 382120
rect 56654 382064 60076 382120
rect 56593 382062 60076 382064
rect 56593 382059 56659 382062
rect 302785 381714 302851 381717
rect 299828 381712 302851 381714
rect 299828 381656 302790 381712
rect 302846 381656 302851 381712
rect 299828 381654 302851 381656
rect 302785 381651 302851 381654
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3325 380626 3391 380629
rect -960 380624 3391 380626
rect -960 380568 3330 380624
rect 3386 380568 3391 380624
rect -960 380566 3391 380568
rect -960 380476 480 380566
rect 3325 380563 3391 380566
rect 56593 380082 56659 380085
rect 56593 380080 60076 380082
rect 56593 380024 56598 380080
rect 56654 380024 60076 380080
rect 56593 380022 60076 380024
rect 56593 380019 56659 380022
rect 302601 379538 302667 379541
rect 299828 379536 302667 379538
rect 299828 379480 302606 379536
rect 302662 379480 302667 379536
rect 299828 379478 302667 379480
rect 302601 379475 302667 379478
rect 56593 377906 56659 377909
rect 56593 377904 60076 377906
rect 56593 377848 56598 377904
rect 56654 377848 60076 377904
rect 56593 377846 60076 377848
rect 56593 377843 56659 377846
rect 302785 377362 302851 377365
rect 299828 377360 302851 377362
rect 299828 377304 302790 377360
rect 302846 377304 302851 377360
rect 299828 377302 302851 377304
rect 302785 377299 302851 377302
rect 56593 375866 56659 375869
rect 56593 375864 60076 375866
rect 56593 375808 56598 375864
rect 56654 375808 60076 375864
rect 56593 375806 60076 375808
rect 56593 375803 56659 375806
rect 302785 375186 302851 375189
rect 299828 375184 302851 375186
rect 299828 375128 302790 375184
rect 302846 375128 302851 375184
rect 299828 375126 302851 375128
rect 302785 375123 302851 375126
rect 56593 373690 56659 373693
rect 56593 373688 60076 373690
rect 56593 373632 56598 373688
rect 56654 373632 60076 373688
rect 56593 373630 60076 373632
rect 56593 373627 56659 373630
rect 302785 373010 302851 373013
rect 299828 373008 302851 373010
rect 299828 372952 302790 373008
rect 302846 372952 302851 373008
rect 299828 372950 302851 372952
rect 302785 372947 302851 372950
rect 56593 371650 56659 371653
rect 56593 371648 60076 371650
rect 56593 371592 56598 371648
rect 56654 371592 60076 371648
rect 56593 371590 60076 371592
rect 56593 371587 56659 371590
rect 302325 370698 302391 370701
rect 299828 370696 302391 370698
rect 299828 370640 302330 370696
rect 302386 370640 302391 370696
rect 299828 370638 302391 370640
rect 302325 370635 302391 370638
rect 580257 369610 580323 369613
rect 583520 369610 584960 369700
rect 580257 369608 584960 369610
rect 580257 369552 580262 369608
rect 580318 369552 584960 369608
rect 580257 369550 584960 369552
rect 580257 369547 580323 369550
rect 56593 369474 56659 369477
rect 56593 369472 60076 369474
rect 56593 369416 56598 369472
rect 56654 369416 60076 369472
rect 583520 369460 584960 369550
rect 56593 369414 60076 369416
rect 56593 369411 56659 369414
rect 302601 368522 302667 368525
rect 299828 368520 302667 368522
rect 299828 368464 302606 368520
rect 302662 368464 302667 368520
rect 299828 368462 302667 368464
rect 302601 368459 302667 368462
rect 56593 367434 56659 367437
rect 56593 367432 60076 367434
rect 56593 367376 56598 367432
rect 56654 367376 60076 367432
rect 56593 367374 60076 367376
rect 56593 367371 56659 367374
rect 327809 367026 327875 367029
rect 328085 367026 328151 367029
rect 327809 367024 328151 367026
rect 327809 366968 327814 367024
rect 327870 366968 328090 367024
rect 328146 366968 328151 367024
rect 327809 366966 328151 366968
rect 327809 366963 327875 366966
rect 328085 366963 328151 366966
rect 302785 366346 302851 366349
rect 299828 366344 302851 366346
rect -960 366210 480 366300
rect 299828 366288 302790 366344
rect 302846 366288 302851 366344
rect 299828 366286 302851 366288
rect 302785 366283 302851 366286
rect 3049 366210 3115 366213
rect -960 366208 3115 366210
rect -960 366152 3054 366208
rect 3110 366152 3115 366208
rect -960 366150 3115 366152
rect -960 366060 480 366150
rect 3049 366147 3115 366150
rect 56593 365258 56659 365261
rect 56593 365256 60076 365258
rect 56593 365200 56598 365256
rect 56654 365200 60076 365256
rect 56593 365198 60076 365200
rect 56593 365195 56659 365198
rect 302509 364170 302575 364173
rect 299828 364168 302575 364170
rect 299828 364112 302514 364168
rect 302570 364112 302575 364168
rect 299828 364110 302575 364112
rect 302509 364107 302575 364110
rect 56593 363218 56659 363221
rect 56593 363216 60076 363218
rect 56593 363160 56598 363216
rect 56654 363160 60076 363216
rect 56593 363158 60076 363160
rect 56593 363155 56659 363158
rect 302417 361994 302483 361997
rect 299828 361992 302483 361994
rect 299828 361936 302422 361992
rect 302478 361936 302483 361992
rect 299828 361934 302483 361936
rect 302417 361931 302483 361934
rect 56593 361042 56659 361045
rect 56593 361040 60076 361042
rect 56593 360984 56598 361040
rect 56654 360984 60076 361040
rect 56593 360982 60076 360984
rect 56593 360979 56659 360982
rect 302325 359682 302391 359685
rect 299828 359680 302391 359682
rect 299828 359624 302330 359680
rect 302386 359624 302391 359680
rect 299828 359622 302391 359624
rect 302325 359619 302391 359622
rect 56593 359002 56659 359005
rect 56593 359000 60076 359002
rect 56593 358944 56598 359000
rect 56654 358944 60076 359000
rect 56593 358942 60076 358944
rect 56593 358939 56659 358942
rect 580349 357914 580415 357917
rect 583520 357914 584960 358004
rect 580349 357912 584960 357914
rect 580349 357856 580354 357912
rect 580410 357856 584960 357912
rect 580349 357854 584960 357856
rect 580349 357851 580415 357854
rect 583520 357764 584960 357854
rect 302509 357506 302575 357509
rect 299828 357504 302575 357506
rect 299828 357448 302514 357504
rect 302570 357448 302575 357504
rect 299828 357446 302575 357448
rect 302509 357443 302575 357446
rect 56593 356826 56659 356829
rect 56593 356824 60076 356826
rect 56593 356768 56598 356824
rect 56654 356768 60076 356824
rect 56593 356766 60076 356768
rect 56593 356763 56659 356766
rect 302785 355330 302851 355333
rect 299828 355328 302851 355330
rect 299828 355272 302790 355328
rect 302846 355272 302851 355328
rect 299828 355270 302851 355272
rect 302785 355267 302851 355270
rect 56593 354786 56659 354789
rect 56593 354784 60076 354786
rect 56593 354728 56598 354784
rect 56654 354728 60076 354784
rect 56593 354726 60076 354728
rect 56593 354723 56659 354726
rect 302785 353154 302851 353157
rect 299828 353152 302851 353154
rect 299828 353096 302790 353152
rect 302846 353096 302851 353152
rect 299828 353094 302851 353096
rect 302785 353091 302851 353094
rect 56593 352610 56659 352613
rect 56593 352608 60076 352610
rect 56593 352552 56598 352608
rect 56654 352552 60076 352608
rect 56593 352550 60076 352552
rect 56593 352547 56659 352550
rect -960 351780 480 352020
rect 302417 350978 302483 350981
rect 299828 350976 302483 350978
rect 299828 350920 302422 350976
rect 302478 350920 302483 350976
rect 299828 350918 302483 350920
rect 302417 350915 302483 350918
rect 56593 350570 56659 350573
rect 56593 350568 60076 350570
rect 56593 350512 56598 350568
rect 56654 350512 60076 350568
rect 56593 350510 60076 350512
rect 56593 350507 56659 350510
rect 302693 348666 302759 348669
rect 299828 348664 302759 348666
rect 299828 348608 302698 348664
rect 302754 348608 302759 348664
rect 299828 348606 302759 348608
rect 302693 348603 302759 348606
rect 56593 348394 56659 348397
rect 56593 348392 60076 348394
rect 56593 348336 56598 348392
rect 56654 348336 60076 348392
rect 56593 348334 60076 348336
rect 56593 348331 56659 348334
rect 302509 346490 302575 346493
rect 299828 346488 302575 346490
rect 299828 346432 302514 346488
rect 302570 346432 302575 346488
rect 299828 346430 302575 346432
rect 302509 346427 302575 346430
rect 56593 346354 56659 346357
rect 56593 346352 60076 346354
rect 56593 346296 56598 346352
rect 56654 346296 60076 346352
rect 56593 346294 60076 346296
rect 56593 346291 56659 346294
rect 580441 346082 580507 346085
rect 583520 346082 584960 346172
rect 580441 346080 584960 346082
rect 580441 346024 580446 346080
rect 580502 346024 584960 346080
rect 580441 346022 584960 346024
rect 580441 346019 580507 346022
rect 583520 345932 584960 346022
rect 302785 344314 302851 344317
rect 299828 344312 302851 344314
rect 299828 344256 302790 344312
rect 302846 344256 302851 344312
rect 299828 344254 302851 344256
rect 302785 344251 302851 344254
rect 58433 344178 58499 344181
rect 58433 344176 60076 344178
rect 58433 344120 58438 344176
rect 58494 344120 60076 344176
rect 58433 344118 60076 344120
rect 58433 344115 58499 344118
rect 58525 342138 58591 342141
rect 302785 342138 302851 342141
rect 58525 342136 60076 342138
rect 58525 342080 58530 342136
rect 58586 342080 60076 342136
rect 58525 342078 60076 342080
rect 299828 342136 302851 342138
rect 299828 342080 302790 342136
rect 302846 342080 302851 342136
rect 299828 342078 302851 342080
rect 58525 342075 58591 342078
rect 302785 342075 302851 342078
rect 59537 339962 59603 339965
rect 302417 339962 302483 339965
rect 59537 339960 60076 339962
rect 59537 339904 59542 339960
rect 59598 339904 60076 339960
rect 59537 339902 60076 339904
rect 299828 339960 302483 339962
rect 299828 339904 302422 339960
rect 302478 339904 302483 339960
rect 299828 339902 302483 339904
rect 59537 339899 59603 339902
rect 302417 339899 302483 339902
rect 58617 337922 58683 337925
rect 58617 337920 60076 337922
rect 58617 337864 58622 337920
rect 58678 337864 60076 337920
rect 58617 337862 60076 337864
rect 58617 337859 58683 337862
rect 302693 337650 302759 337653
rect 299828 337648 302759 337650
rect -960 337514 480 337604
rect 299828 337592 302698 337648
rect 302754 337592 302759 337648
rect 299828 337590 302759 337592
rect 302693 337587 302759 337590
rect 3233 337514 3299 337517
rect -960 337512 3299 337514
rect -960 337456 3238 337512
rect 3294 337456 3299 337512
rect -960 337454 3299 337456
rect -960 337364 480 337454
rect 3233 337451 3299 337454
rect 58709 335746 58775 335749
rect 58709 335744 60076 335746
rect 58709 335688 58714 335744
rect 58770 335688 60076 335744
rect 58709 335686 60076 335688
rect 58709 335683 58775 335686
rect 302509 335474 302575 335477
rect 299828 335472 302575 335474
rect 299828 335416 302514 335472
rect 302570 335416 302575 335472
rect 299828 335414 302575 335416
rect 302509 335411 302575 335414
rect 583520 334236 584960 334476
rect 57697 333706 57763 333709
rect 57697 333704 60076 333706
rect 57697 333648 57702 333704
rect 57758 333648 60076 333704
rect 57697 333646 60076 333648
rect 57697 333643 57763 333646
rect 302785 333298 302851 333301
rect 299828 333296 302851 333298
rect 299828 333240 302790 333296
rect 302846 333240 302851 333296
rect 299828 333238 302851 333240
rect 302785 333235 302851 333238
rect 57789 331530 57855 331533
rect 57789 331528 60076 331530
rect 57789 331472 57794 331528
rect 57850 331472 60076 331528
rect 57789 331470 60076 331472
rect 57789 331467 57855 331470
rect 302509 331122 302575 331125
rect 299828 331120 302575 331122
rect 299828 331064 302514 331120
rect 302570 331064 302575 331120
rect 299828 331062 302575 331064
rect 302509 331059 302575 331062
rect 58801 329490 58867 329493
rect 58801 329488 60076 329490
rect 58801 329432 58806 329488
rect 58862 329432 60076 329488
rect 58801 329430 60076 329432
rect 58801 329427 58867 329430
rect 302325 328946 302391 328949
rect 299828 328944 302391 328946
rect 299828 328888 302330 328944
rect 302386 328888 302391 328944
rect 299828 328886 302391 328888
rect 302325 328883 302391 328886
rect 56777 327314 56843 327317
rect 56777 327312 60076 327314
rect 56777 327256 56782 327312
rect 56838 327256 60076 327312
rect 56777 327254 60076 327256
rect 56777 327251 56843 327254
rect 302509 326634 302575 326637
rect 299828 326632 302575 326634
rect 299828 326576 302514 326632
rect 302570 326576 302575 326632
rect 299828 326574 302575 326576
rect 302509 326571 302575 326574
rect 59445 325274 59511 325277
rect 59445 325272 60076 325274
rect 59445 325216 59450 325272
rect 59506 325216 60076 325272
rect 59445 325214 60076 325216
rect 59445 325211 59511 325214
rect 302325 324458 302391 324461
rect 299828 324456 302391 324458
rect 299828 324400 302330 324456
rect 302386 324400 302391 324456
rect 299828 324398 302391 324400
rect 302325 324395 302391 324398
rect -960 323098 480 323188
rect 4061 323098 4127 323101
rect -960 323096 4127 323098
rect -960 323040 4066 323096
rect 4122 323040 4127 323096
rect -960 323038 4127 323040
rect -960 322948 480 323038
rect 4061 323035 4127 323038
rect 58893 323098 58959 323101
rect 58893 323096 60076 323098
rect 58893 323040 58898 323096
rect 58954 323040 60076 323096
rect 58893 323038 60076 323040
rect 58893 323035 58959 323038
rect 580533 322690 580599 322693
rect 583520 322690 584960 322780
rect 580533 322688 584960 322690
rect 580533 322632 580538 322688
rect 580594 322632 584960 322688
rect 580533 322630 584960 322632
rect 580533 322627 580599 322630
rect 583520 322540 584960 322630
rect 302325 322282 302391 322285
rect 299828 322280 302391 322282
rect 299828 322224 302330 322280
rect 302386 322224 302391 322280
rect 299828 322222 302391 322224
rect 302325 322219 302391 322222
rect 56869 321058 56935 321061
rect 56869 321056 60076 321058
rect 56869 321000 56874 321056
rect 56930 321000 60076 321056
rect 56869 320998 60076 321000
rect 56869 320995 56935 320998
rect 302325 320106 302391 320109
rect 299828 320104 302391 320106
rect 299828 320048 302330 320104
rect 302386 320048 302391 320104
rect 299828 320046 302391 320048
rect 302325 320043 302391 320046
rect 57881 319018 57947 319021
rect 57881 319016 60076 319018
rect 57881 318960 57886 319016
rect 57942 318960 60076 319016
rect 57881 318958 60076 318960
rect 57881 318955 57947 318958
rect 302693 317930 302759 317933
rect 299828 317928 302759 317930
rect 299828 317872 302698 317928
rect 302754 317872 302759 317928
rect 299828 317870 302759 317872
rect 302693 317867 302759 317870
rect 58985 316842 59051 316845
rect 58985 316840 60076 316842
rect 58985 316784 58990 316840
rect 59046 316784 60076 316840
rect 58985 316782 60076 316784
rect 58985 316779 59051 316782
rect 302785 315754 302851 315757
rect 299828 315752 302851 315754
rect 299828 315696 302790 315752
rect 302846 315696 302851 315752
rect 299828 315694 302851 315696
rect 302785 315691 302851 315694
rect 56961 314802 57027 314805
rect 56961 314800 60076 314802
rect 56961 314744 56966 314800
rect 57022 314744 60076 314800
rect 56961 314742 60076 314744
rect 56961 314739 57027 314742
rect 302785 313442 302851 313445
rect 299828 313440 302851 313442
rect 299828 313384 302790 313440
rect 302846 313384 302851 313440
rect 299828 313382 302851 313384
rect 302785 313379 302851 313382
rect 59077 312626 59143 312629
rect 59077 312624 60076 312626
rect 59077 312568 59082 312624
rect 59138 312568 60076 312624
rect 59077 312566 60076 312568
rect 59077 312563 59143 312566
rect 302693 311266 302759 311269
rect 299828 311264 302759 311266
rect 299828 311208 302698 311264
rect 302754 311208 302759 311264
rect 299828 311206 302759 311208
rect 302693 311203 302759 311206
rect 580625 310858 580691 310861
rect 583520 310858 584960 310948
rect 580625 310856 584960 310858
rect 580625 310800 580630 310856
rect 580686 310800 584960 310856
rect 580625 310798 584960 310800
rect 580625 310795 580691 310798
rect 583520 310708 584960 310798
rect 59169 310586 59235 310589
rect 59169 310584 60076 310586
rect 59169 310528 59174 310584
rect 59230 310528 60076 310584
rect 59169 310526 60076 310528
rect 59169 310523 59235 310526
rect 302785 309090 302851 309093
rect 299828 309088 302851 309090
rect 299828 309032 302790 309088
rect 302846 309032 302851 309088
rect 299828 309030 302851 309032
rect 302785 309027 302851 309030
rect -960 308818 480 308908
rect 3877 308818 3943 308821
rect -960 308816 3943 308818
rect -960 308760 3882 308816
rect 3938 308760 3943 308816
rect -960 308758 3943 308760
rect -960 308668 480 308758
rect 3877 308755 3943 308758
rect 57053 308410 57119 308413
rect 57053 308408 60076 308410
rect 57053 308352 57058 308408
rect 57114 308352 60076 308408
rect 57053 308350 60076 308352
rect 57053 308347 57119 308350
rect 302785 306914 302851 306917
rect 299828 306912 302851 306914
rect 299828 306856 302790 306912
rect 302846 306856 302851 306912
rect 299828 306854 302851 306856
rect 302785 306851 302851 306854
rect 57462 306308 57468 306372
rect 57532 306370 57538 306372
rect 57532 306310 60076 306370
rect 57532 306308 57538 306310
rect 302785 304738 302851 304741
rect 299828 304736 302851 304738
rect 299828 304680 302790 304736
rect 302846 304680 302851 304736
rect 299828 304678 302851 304680
rect 302785 304675 302851 304678
rect 59261 304194 59327 304197
rect 59261 304192 60076 304194
rect 59261 304136 59266 304192
rect 59322 304136 60076 304192
rect 59261 304134 60076 304136
rect 59261 304131 59327 304134
rect 302785 302426 302851 302429
rect 299828 302424 302851 302426
rect 299828 302368 302790 302424
rect 302846 302368 302851 302424
rect 299828 302366 302851 302368
rect 302785 302363 302851 302366
rect 57646 302092 57652 302156
rect 57716 302154 57722 302156
rect 57716 302094 60076 302154
rect 57716 302092 57722 302094
rect 302693 300250 302759 300253
rect 299828 300248 302759 300250
rect 299828 300192 302698 300248
rect 302754 300192 302759 300248
rect 299828 300190 302759 300192
rect 302693 300187 302759 300190
rect 57830 299916 57836 299980
rect 57900 299978 57906 299980
rect 57900 299918 60076 299978
rect 57900 299916 57906 299918
rect 580717 299162 580783 299165
rect 583520 299162 584960 299252
rect 580717 299160 584960 299162
rect 580717 299104 580722 299160
rect 580778 299104 584960 299160
rect 580717 299102 584960 299104
rect 580717 299099 580783 299102
rect 583520 299012 584960 299102
rect 302785 298074 302851 298077
rect 299828 298072 302851 298074
rect 299828 298016 302790 298072
rect 302846 298016 302851 298072
rect 299828 298014 302851 298016
rect 302785 298011 302851 298014
rect 59118 297876 59124 297940
rect 59188 297938 59194 297940
rect 59188 297878 60076 297938
rect 59188 297876 59194 297878
rect 302601 295898 302667 295901
rect 299828 295896 302667 295898
rect 299828 295840 302606 295896
rect 302662 295840 302667 295896
rect 299828 295838 302667 295840
rect 302601 295835 302667 295838
rect 56910 295700 56916 295764
rect 56980 295762 56986 295764
rect 56980 295702 60076 295762
rect 56980 295700 56986 295702
rect -960 294402 480 294492
rect 3049 294402 3115 294405
rect -960 294400 3115 294402
rect -960 294344 3054 294400
rect 3110 294344 3115 294400
rect -960 294342 3115 294344
rect -960 294252 480 294342
rect 3049 294339 3115 294342
rect 59353 293722 59419 293725
rect 302785 293722 302851 293725
rect 59353 293720 60076 293722
rect 59353 293664 59358 293720
rect 59414 293664 60076 293720
rect 59353 293662 60076 293664
rect 299828 293720 302851 293722
rect 299828 293664 302790 293720
rect 302846 293664 302851 293720
rect 299828 293662 302851 293664
rect 59353 293659 59419 293662
rect 302785 293659 302851 293662
rect 58750 291484 58756 291548
rect 58820 291546 58826 291548
rect 58820 291486 60076 291546
rect 58820 291484 58826 291486
rect 302509 291410 302575 291413
rect 299828 291408 302575 291410
rect 299828 291352 302514 291408
rect 302570 291352 302575 291408
rect 299828 291350 302575 291352
rect 302509 291347 302575 291350
rect 57278 289444 57284 289508
rect 57348 289506 57354 289508
rect 57348 289446 60076 289506
rect 57348 289444 57354 289446
rect 302693 289234 302759 289237
rect 299828 289232 302759 289234
rect 299828 289176 302698 289232
rect 302754 289176 302759 289232
rect 299828 289174 302759 289176
rect 302693 289171 302759 289174
rect 59629 287330 59695 287333
rect 59629 287328 60076 287330
rect 59629 287272 59634 287328
rect 59690 287272 60076 287328
rect 583520 287316 584960 287556
rect 59629 287270 60076 287272
rect 59629 287267 59695 287270
rect 302785 287058 302851 287061
rect 299828 287056 302851 287058
rect 299828 287000 302790 287056
rect 302846 287000 302851 287056
rect 299828 286998 302851 287000
rect 302785 286995 302851 286998
rect 58198 285228 58204 285292
rect 58268 285290 58274 285292
rect 58268 285230 60076 285290
rect 58268 285228 58274 285230
rect 302693 284882 302759 284885
rect 299828 284880 302759 284882
rect 299828 284824 302698 284880
rect 302754 284824 302759 284880
rect 299828 284822 302759 284824
rect 302693 284819 302759 284822
rect 58014 283052 58020 283116
rect 58084 283114 58090 283116
rect 58084 283054 60076 283114
rect 58084 283052 58090 283054
rect 302509 282706 302575 282709
rect 299828 282704 302575 282706
rect 299828 282648 302514 282704
rect 302570 282648 302575 282704
rect 299828 282646 302575 282648
rect 302509 282643 302575 282646
rect 59721 281074 59787 281077
rect 59721 281072 60076 281074
rect 59721 281016 59726 281072
rect 59782 281016 60076 281072
rect 59721 281014 60076 281016
rect 59721 281011 59787 281014
rect 302509 280394 302575 280397
rect 299828 280392 302575 280394
rect 299828 280336 302514 280392
rect 302570 280336 302575 280392
rect 299828 280334 302575 280336
rect 302509 280331 302575 280334
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 58934 278836 58940 278900
rect 59004 278898 59010 278900
rect 59004 278838 60076 278898
rect 59004 278836 59010 278838
rect 302325 278218 302391 278221
rect 299828 278216 302391 278218
rect 299828 278160 302330 278216
rect 302386 278160 302391 278216
rect 299828 278158 302391 278160
rect 302325 278155 302391 278158
rect 58341 276858 58407 276861
rect 58341 276856 60076 276858
rect 58341 276800 58346 276856
rect 58402 276800 60076 276856
rect 58341 276798 60076 276800
rect 58341 276795 58407 276798
rect 302601 276042 302667 276045
rect 299828 276040 302667 276042
rect 299828 275984 302606 276040
rect 302662 275984 302667 276040
rect 299828 275982 302667 275984
rect 302601 275979 302667 275982
rect 580809 275770 580875 275773
rect 583520 275770 584960 275860
rect 580809 275768 584960 275770
rect 580809 275712 580814 275768
rect 580870 275712 584960 275768
rect 580809 275710 584960 275712
rect 580809 275707 580875 275710
rect 583520 275620 584960 275710
rect 56726 274620 56732 274684
rect 56796 274682 56802 274684
rect 56796 274622 60076 274682
rect 56796 274620 56802 274622
rect 302785 273866 302851 273869
rect 299828 273864 302851 273866
rect 299828 273808 302790 273864
rect 302846 273808 302851 273864
rect 299828 273806 302851 273808
rect 302785 273803 302851 273806
rect 58249 272642 58315 272645
rect 58249 272640 60076 272642
rect 58249 272584 58254 272640
rect 58310 272584 60076 272640
rect 58249 272582 60076 272584
rect 58249 272579 58315 272582
rect 302509 271690 302575 271693
rect 299828 271688 302575 271690
rect 299828 271632 302514 271688
rect 302570 271632 302575 271688
rect 299828 271630 302575 271632
rect 302509 271627 302575 271630
rect 57973 270466 58039 270469
rect 57973 270464 60076 270466
rect 57973 270408 57978 270464
rect 58034 270408 60076 270464
rect 57973 270406 60076 270408
rect 57973 270403 58039 270406
rect 302509 269378 302575 269381
rect 299828 269376 302575 269378
rect 299828 269320 302514 269376
rect 302570 269320 302575 269376
rect 299828 269318 302575 269320
rect 302509 269315 302575 269318
rect 57237 268426 57303 268429
rect 57237 268424 60076 268426
rect 57237 268368 57242 268424
rect 57298 268368 60076 268424
rect 57237 268366 60076 268368
rect 57237 268363 57303 268366
rect 302325 267202 302391 267205
rect 299828 267200 302391 267202
rect 299828 267144 302330 267200
rect 302386 267144 302391 267200
rect 299828 267142 302391 267144
rect 302325 267139 302391 267142
rect 57094 266188 57100 266252
rect 57164 266250 57170 266252
rect 57164 266190 60076 266250
rect 57164 266188 57170 266190
rect -960 265706 480 265796
rect 2773 265706 2839 265709
rect -960 265704 2839 265706
rect -960 265648 2778 265704
rect 2834 265648 2839 265704
rect -960 265646 2839 265648
rect -960 265556 480 265646
rect 2773 265643 2839 265646
rect 302601 265026 302667 265029
rect 299828 265024 302667 265026
rect 299828 264968 302606 265024
rect 302662 264968 302667 265024
rect 299828 264966 302667 264968
rect 302601 264963 302667 264966
rect 58065 264210 58131 264213
rect 58065 264208 60076 264210
rect 58065 264152 58070 264208
rect 58126 264152 60076 264208
rect 58065 264150 60076 264152
rect 58065 264147 58131 264150
rect 580901 263938 580967 263941
rect 583520 263938 584960 264028
rect 580901 263936 584960 263938
rect 580901 263880 580906 263936
rect 580962 263880 584960 263936
rect 580901 263878 584960 263880
rect 580901 263875 580967 263878
rect 583520 263788 584960 263878
rect 302785 262850 302851 262853
rect 299828 262848 302851 262850
rect 299828 262792 302790 262848
rect 302846 262792 302851 262848
rect 299828 262790 302851 262792
rect 302785 262787 302851 262790
rect 57605 262034 57671 262037
rect 57605 262032 60076 262034
rect 57605 261976 57610 262032
rect 57666 261976 60076 262032
rect 57605 261974 60076 261976
rect 57605 261971 57671 261974
rect 302509 260674 302575 260677
rect 299828 260672 302575 260674
rect 299828 260616 302514 260672
rect 302570 260616 302575 260672
rect 299828 260614 302575 260616
rect 302509 260611 302575 260614
rect 57329 259994 57395 259997
rect 57329 259992 60076 259994
rect 57329 259936 57334 259992
rect 57390 259936 60076 259992
rect 57329 259934 60076 259936
rect 57329 259931 57395 259934
rect 302417 258498 302483 258501
rect 299828 258496 302483 258498
rect 299828 258440 302422 258496
rect 302478 258440 302483 258496
rect 299828 258438 302483 258440
rect 302417 258435 302483 258438
rect 58157 257954 58223 257957
rect 58157 257952 60076 257954
rect 58157 257896 58162 257952
rect 58218 257896 60076 257952
rect 58157 257894 60076 257896
rect 58157 257891 58223 257894
rect 302325 256186 302391 256189
rect 299828 256184 302391 256186
rect 299828 256128 302330 256184
rect 302386 256128 302391 256184
rect 299828 256126 302391 256128
rect 302325 256123 302391 256126
rect 57789 255778 57855 255781
rect 57789 255776 60076 255778
rect 57789 255720 57794 255776
rect 57850 255720 60076 255776
rect 57789 255718 60076 255720
rect 57789 255715 57855 255718
rect 302509 254010 302575 254013
rect 299828 254008 302575 254010
rect 299828 253952 302514 254008
rect 302570 253952 302575 254008
rect 299828 253950 302575 253952
rect 302509 253947 302575 253950
rect 57421 253738 57487 253741
rect 57421 253736 60076 253738
rect 57421 253680 57426 253736
rect 57482 253680 60076 253736
rect 57421 253678 60076 253680
rect 57421 253675 57487 253678
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect 302785 251834 302851 251837
rect 299828 251832 302851 251834
rect 299828 251776 302790 251832
rect 302846 251776 302851 251832
rect 299828 251774 302851 251776
rect 302785 251771 302851 251774
rect 57513 251562 57579 251565
rect 57513 251560 60076 251562
rect 57513 251504 57518 251560
rect 57574 251504 60076 251560
rect 57513 251502 60076 251504
rect 57513 251499 57579 251502
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 302785 249658 302851 249661
rect 299828 249656 302851 249658
rect 299828 249600 302790 249656
rect 302846 249600 302851 249656
rect 299828 249598 302851 249600
rect 302785 249595 302851 249598
rect 57646 249460 57652 249524
rect 57716 249522 57722 249524
rect 57716 249462 60076 249522
rect 57716 249460 57722 249462
rect 302417 247482 302483 247485
rect 299828 247480 302483 247482
rect 299828 247424 302422 247480
rect 302478 247424 302483 247480
rect 299828 247422 302483 247424
rect 302417 247419 302483 247422
rect 57830 247284 57836 247348
rect 57900 247346 57906 247348
rect 57900 247286 60076 247346
rect 57900 247284 57906 247286
rect 57881 245306 57947 245309
rect 57881 245304 60076 245306
rect 57881 245248 57886 245304
rect 57942 245248 60076 245304
rect 57881 245246 60076 245248
rect 57881 245243 57947 245246
rect 302693 245170 302759 245173
rect 299828 245168 302759 245170
rect 299828 245112 302698 245168
rect 302754 245112 302759 245168
rect 299828 245110 302759 245112
rect 302693 245107 302759 245110
rect 56869 243130 56935 243133
rect 56869 243128 60076 243130
rect 56869 243072 56874 243128
rect 56930 243072 60076 243128
rect 56869 243070 60076 243072
rect 56869 243067 56935 243070
rect 302509 242994 302575 242997
rect 299828 242992 302575 242994
rect 299828 242936 302514 242992
rect 302570 242936 302575 242992
rect 299828 242934 302575 242936
rect 302509 242931 302575 242934
rect 57697 241090 57763 241093
rect 57697 241088 60076 241090
rect 57697 241032 57702 241088
rect 57758 241032 60076 241088
rect 57697 241030 60076 241032
rect 57697 241027 57763 241030
rect 302785 240818 302851 240821
rect 299828 240816 302851 240818
rect 299828 240760 302790 240816
rect 302846 240760 302851 240816
rect 299828 240758 302851 240760
rect 302785 240755 302851 240758
rect 583520 240396 584960 240636
rect 57237 238914 57303 238917
rect 57237 238912 60076 238914
rect 57237 238856 57242 238912
rect 57298 238856 60076 238912
rect 57237 238854 60076 238856
rect 57237 238851 57303 238854
rect 302785 238642 302851 238645
rect 299828 238640 302851 238642
rect 299828 238584 302790 238640
rect 302846 238584 302851 238640
rect 299828 238582 302851 238584
rect 302785 238579 302851 238582
rect -960 237010 480 237100
rect 3417 237010 3483 237013
rect -960 237008 3483 237010
rect -960 236952 3422 237008
rect 3478 236952 3483 237008
rect -960 236950 3483 236952
rect -960 236860 480 236950
rect 3417 236947 3483 236950
rect 57605 236874 57671 236877
rect 57605 236872 60076 236874
rect 57605 236816 57610 236872
rect 57666 236816 60076 236872
rect 57605 236814 60076 236816
rect 57605 236811 57671 236814
rect 302417 236466 302483 236469
rect 299828 236464 302483 236466
rect 299828 236408 302422 236464
rect 302478 236408 302483 236464
rect 299828 236406 302483 236408
rect 302417 236403 302483 236406
rect 57145 234698 57211 234701
rect 57145 234696 60076 234698
rect 57145 234640 57150 234696
rect 57206 234640 60076 234696
rect 57145 234638 60076 234640
rect 57145 234635 57211 234638
rect 302693 234154 302759 234157
rect 299828 234152 302759 234154
rect 299828 234096 302698 234152
rect 302754 234096 302759 234152
rect 299828 234094 302759 234096
rect 302693 234091 302759 234094
rect 56961 232658 57027 232661
rect 56961 232656 60076 232658
rect 56961 232600 56966 232656
rect 57022 232600 60076 232656
rect 56961 232598 60076 232600
rect 56961 232595 57027 232598
rect 302509 231978 302575 231981
rect 299828 231976 302575 231978
rect 299828 231920 302514 231976
rect 302570 231920 302575 231976
rect 299828 231918 302575 231920
rect 302509 231915 302575 231918
rect 57053 230482 57119 230485
rect 57053 230480 60076 230482
rect 57053 230424 57058 230480
rect 57114 230424 60076 230480
rect 57053 230422 60076 230424
rect 57053 230419 57119 230422
rect 302785 229802 302851 229805
rect 299828 229800 302851 229802
rect 299828 229744 302790 229800
rect 302846 229744 302851 229800
rect 299828 229742 302851 229744
rect 302785 229739 302851 229742
rect 580073 228850 580139 228853
rect 583520 228850 584960 228940
rect 580073 228848 584960 228850
rect 580073 228792 580078 228848
rect 580134 228792 584960 228848
rect 580073 228790 584960 228792
rect 580073 228787 580139 228790
rect 583520 228700 584960 228790
rect 57789 228442 57855 228445
rect 57789 228440 60076 228442
rect 57789 228384 57794 228440
rect 57850 228384 60076 228440
rect 57789 228382 60076 228384
rect 57789 228379 57855 228382
rect 302785 227626 302851 227629
rect 299828 227624 302851 227626
rect 299828 227568 302790 227624
rect 302846 227568 302851 227624
rect 299828 227566 302851 227568
rect 302785 227563 302851 227566
rect 57513 226266 57579 226269
rect 57513 226264 60076 226266
rect 57513 226208 57518 226264
rect 57574 226208 60076 226264
rect 57513 226206 60076 226208
rect 57513 226203 57579 226206
rect 302785 225450 302851 225453
rect 299828 225448 302851 225450
rect 299828 225392 302790 225448
rect 302846 225392 302851 225448
rect 299828 225390 302851 225392
rect 302785 225387 302851 225390
rect 57421 224226 57487 224229
rect 57421 224224 60076 224226
rect 57421 224168 57426 224224
rect 57482 224168 60076 224224
rect 57421 224166 60076 224168
rect 57421 224163 57487 224166
rect 302693 223138 302759 223141
rect 299828 223136 302759 223138
rect 299828 223080 302698 223136
rect 302754 223080 302759 223136
rect 299828 223078 302759 223080
rect 302693 223075 302759 223078
rect -960 222594 480 222684
rect 2773 222594 2839 222597
rect -960 222592 2839 222594
rect -960 222536 2778 222592
rect 2834 222536 2839 222592
rect -960 222534 2839 222536
rect -960 222444 480 222534
rect 2773 222531 2839 222534
rect 57329 222050 57395 222053
rect 57329 222048 60076 222050
rect 57329 221992 57334 222048
rect 57390 221992 60076 222048
rect 57329 221990 60076 221992
rect 57329 221987 57395 221990
rect 302785 220962 302851 220965
rect 299828 220960 302851 220962
rect 299828 220904 302790 220960
rect 302846 220904 302851 220960
rect 299828 220902 302851 220904
rect 302785 220899 302851 220902
rect 56777 220010 56843 220013
rect 56777 220008 60076 220010
rect 56777 219952 56782 220008
rect 56838 219952 60076 220008
rect 56777 219950 60076 219952
rect 56777 219947 56843 219950
rect 302785 218786 302851 218789
rect 299828 218784 302851 218786
rect 299828 218728 302790 218784
rect 302846 218728 302851 218784
rect 299828 218726 302851 218728
rect 302785 218723 302851 218726
rect 56685 217834 56751 217837
rect 56685 217832 60076 217834
rect 56685 217776 56690 217832
rect 56746 217776 60076 217832
rect 56685 217774 60076 217776
rect 56685 217771 56751 217774
rect 579981 217018 580047 217021
rect 583520 217018 584960 217108
rect 579981 217016 584960 217018
rect 579981 216960 579986 217016
rect 580042 216960 584960 217016
rect 579981 216958 584960 216960
rect 579981 216955 580047 216958
rect 583520 216868 584960 216958
rect 302785 216610 302851 216613
rect 299828 216608 302851 216610
rect 299828 216552 302790 216608
rect 302846 216552 302851 216608
rect 299828 216550 302851 216552
rect 302785 216547 302851 216550
rect 56593 215794 56659 215797
rect 56593 215792 60076 215794
rect 56593 215736 56598 215792
rect 56654 215736 60076 215792
rect 56593 215734 60076 215736
rect 56593 215731 56659 215734
rect 302785 214434 302851 214437
rect 299828 214432 302851 214434
rect 299828 214376 302790 214432
rect 302846 214376 302851 214432
rect 299828 214374 302851 214376
rect 302785 214371 302851 214374
rect 56910 213556 56916 213620
rect 56980 213618 56986 213620
rect 56980 213558 60076 213618
rect 56980 213556 56986 213558
rect 302601 212122 302667 212125
rect 299828 212120 302667 212122
rect 299828 212064 302606 212120
rect 302662 212064 302667 212120
rect 299828 212062 302667 212064
rect 302601 212059 302667 212062
rect 57278 211516 57284 211580
rect 57348 211578 57354 211580
rect 57348 211518 60076 211578
rect 57348 211516 57354 211518
rect 302785 209946 302851 209949
rect 299828 209944 302851 209946
rect 299828 209888 302790 209944
rect 302846 209888 302851 209944
rect 299828 209886 302851 209888
rect 302785 209883 302851 209886
rect 57094 209340 57100 209404
rect 57164 209402 57170 209404
rect 57164 209342 60076 209402
rect 57164 209340 57170 209342
rect -960 208178 480 208268
rect 3509 208178 3575 208181
rect -960 208176 3575 208178
rect -960 208120 3514 208176
rect 3570 208120 3575 208176
rect -960 208118 3575 208120
rect -960 208028 480 208118
rect 3509 208115 3575 208118
rect 302785 207770 302851 207773
rect 299828 207768 302851 207770
rect 299828 207712 302790 207768
rect 302846 207712 302851 207768
rect 299828 207710 302851 207712
rect 302785 207707 302851 207710
rect 57462 207300 57468 207364
rect 57532 207362 57538 207364
rect 57532 207302 60076 207362
rect 57532 207300 57538 207302
rect 302785 205594 302851 205597
rect 299828 205592 302851 205594
rect 299828 205536 302790 205592
rect 302846 205536 302851 205592
rect 299828 205534 302851 205536
rect 302785 205531 302851 205534
rect 580165 205322 580231 205325
rect 583520 205322 584960 205412
rect 580165 205320 584960 205322
rect 580165 205264 580170 205320
rect 580226 205264 584960 205320
rect 580165 205262 584960 205264
rect 580165 205259 580231 205262
rect 56726 205124 56732 205188
rect 56796 205186 56802 205188
rect 56796 205126 60076 205186
rect 583520 205172 584960 205262
rect 56796 205124 56802 205126
rect 57646 204988 57652 205052
rect 57716 205050 57722 205052
rect 59813 205050 59879 205053
rect 57716 205048 59879 205050
rect 57716 204992 59818 205048
rect 59874 204992 59879 205048
rect 57716 204990 59879 204992
rect 57716 204988 57722 204990
rect 59813 204987 59879 204990
rect 302233 203418 302299 203421
rect 299828 203416 302299 203418
rect 299828 203360 302238 203416
rect 302294 203360 302299 203416
rect 299828 203358 302299 203360
rect 302233 203355 302299 203358
rect 57646 203084 57652 203148
rect 57716 203146 57722 203148
rect 57716 203086 60076 203146
rect 57716 203084 57722 203086
rect 302877 201242 302943 201245
rect 299828 201240 302943 201242
rect 299828 201184 302882 201240
rect 302938 201184 302943 201240
rect 299828 201182 302943 201184
rect 302877 201179 302943 201182
rect 57789 201106 57855 201109
rect 57789 201104 60076 201106
rect 57789 201048 57794 201104
rect 57850 201048 60076 201104
rect 57789 201046 60076 201048
rect 57789 201043 57855 201046
rect 57830 200636 57836 200700
rect 57900 200698 57906 200700
rect 580257 200698 580323 200701
rect 57900 200696 580323 200698
rect 57900 200640 580262 200696
rect 580318 200640 580323 200696
rect 57900 200638 580323 200640
rect 57900 200636 57906 200638
rect 580257 200635 580323 200638
rect 115841 198114 115907 198117
rect 264881 198114 264947 198117
rect 115841 198112 264947 198114
rect 115841 198056 115846 198112
rect 115902 198056 264886 198112
rect 264942 198056 264947 198112
rect 115841 198054 264947 198056
rect 115841 198051 115907 198054
rect 264881 198051 264947 198054
rect 117221 197978 117287 197981
rect 269113 197978 269179 197981
rect 117221 197976 269179 197978
rect 117221 197920 117226 197976
rect 117282 197920 269118 197976
rect 269174 197920 269179 197976
rect 117221 197918 269179 197920
rect 117221 197915 117287 197918
rect 269113 197915 269179 197918
rect -960 193898 480 193988
rect 3141 193898 3207 193901
rect -960 193896 3207 193898
rect -960 193840 3146 193896
rect 3202 193840 3207 193896
rect -960 193838 3207 193840
rect -960 193748 480 193838
rect 3141 193835 3207 193838
rect 583520 193476 584960 193716
rect 92197 193218 92263 193221
rect 92381 193218 92447 193221
rect 92197 193216 92447 193218
rect 92197 193160 92202 193216
rect 92258 193160 92386 193216
rect 92442 193160 92447 193216
rect 92197 193158 92447 193160
rect 92197 193155 92263 193158
rect 92381 193155 92447 193158
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 92197 173906 92263 173909
rect 92381 173906 92447 173909
rect 92197 173904 92447 173906
rect 92197 173848 92202 173904
rect 92258 173848 92386 173904
rect 92442 173848 92447 173904
rect 92197 173846 92447 173848
rect 92197 173843 92263 173846
rect 92381 173843 92447 173846
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 2773 165066 2839 165069
rect -960 165064 2839 165066
rect -960 165008 2778 165064
rect 2834 165008 2839 165064
rect -960 165006 2839 165008
rect -960 164916 480 165006
rect 2773 165003 2839 165006
rect 92197 164250 92263 164253
rect 92381 164250 92447 164253
rect 92197 164248 92447 164250
rect 92197 164192 92202 164248
rect 92258 164192 92386 164248
rect 92442 164192 92447 164248
rect 92197 164190 92447 164192
rect 92197 164187 92263 164190
rect 92381 164187 92447 164190
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 583520 146556 584960 146796
rect 92197 144938 92263 144941
rect 92381 144938 92447 144941
rect 92197 144936 92447 144938
rect 92197 144880 92202 144936
rect 92258 144880 92386 144936
rect 92442 144880 92447 144936
rect 92197 144878 92447 144880
rect 92197 144875 92263 144878
rect 92381 144875 92447 144878
rect -960 136370 480 136460
rect 3233 136370 3299 136373
rect -960 136368 3299 136370
rect -960 136312 3238 136368
rect 3294 136312 3299 136368
rect -960 136310 3299 136312
rect -960 136220 480 136310
rect 3233 136307 3299 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 92105 125626 92171 125629
rect 92381 125626 92447 125629
rect 92105 125624 92447 125626
rect 92105 125568 92110 125624
rect 92166 125568 92386 125624
rect 92442 125568 92447 125624
rect 92105 125566 92447 125568
rect 92105 125563 92171 125566
rect 92381 125563 92447 125566
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 2773 122090 2839 122093
rect -960 122088 2839 122090
rect -960 122032 2778 122088
rect 2834 122032 2839 122088
rect -960 122030 2839 122032
rect -960 121940 480 122030
rect 2773 122027 2839 122030
rect 583520 111482 584960 111572
rect 583342 111422 584960 111482
rect 125542 111012 125548 111076
rect 125612 111074 125618 111076
rect 135161 111074 135227 111077
rect 125612 111072 135227 111074
rect 125612 111016 135166 111072
rect 135222 111016 135227 111072
rect 125612 111014 135227 111016
rect 125612 111012 125618 111014
rect 135161 111011 135227 111014
rect 115790 110938 115796 110940
rect 108806 110878 115796 110938
rect 56910 110740 56916 110804
rect 56980 110802 56986 110804
rect 89621 110802 89687 110805
rect 56980 110742 64890 110802
rect 56980 110740 56986 110742
rect 64830 110666 64890 110742
rect 74582 110800 89687 110802
rect 74582 110744 89626 110800
rect 89682 110744 89687 110800
rect 74582 110742 89687 110744
rect 64830 110606 74458 110666
rect 74398 110530 74458 110606
rect 74582 110530 74642 110742
rect 89621 110739 89687 110742
rect 96521 110802 96587 110805
rect 96521 110800 99298 110802
rect 96521 110744 96526 110800
rect 96582 110744 99298 110800
rect 96521 110742 99298 110744
rect 96521 110739 96587 110742
rect 74398 110470 74642 110530
rect 99238 110530 99298 110742
rect 108806 110666 108866 110878
rect 115790 110876 115796 110878
rect 115860 110876 115866 110940
rect 140037 110938 140103 110941
rect 135302 110936 140103 110938
rect 135302 110880 140042 110936
rect 140098 110880 140103 110936
rect 135302 110878 140103 110880
rect 118785 110802 118851 110805
rect 125542 110802 125548 110804
rect 118785 110800 125548 110802
rect 118785 110744 118790 110800
rect 118846 110744 125548 110800
rect 118785 110742 125548 110744
rect 118785 110739 118851 110742
rect 125542 110740 125548 110742
rect 125612 110740 125618 110804
rect 99422 110606 108866 110666
rect 135161 110666 135227 110669
rect 135302 110666 135362 110878
rect 140037 110875 140103 110878
rect 154481 110802 154547 110805
rect 154481 110800 161490 110802
rect 154481 110744 154486 110800
rect 154542 110744 161490 110800
rect 154481 110742 161490 110744
rect 154481 110739 154547 110742
rect 147581 110666 147647 110669
rect 135161 110664 135362 110666
rect 135161 110608 135166 110664
rect 135222 110608 135362 110664
rect 135161 110606 135362 110608
rect 144870 110664 147647 110666
rect 144870 110608 147586 110664
rect 147642 110608 147647 110664
rect 144870 110606 147647 110608
rect 161430 110666 161490 110742
rect 171182 110742 180810 110802
rect 161430 110606 171058 110666
rect 99422 110530 99482 110606
rect 135161 110603 135227 110606
rect 99238 110470 99482 110530
rect 115790 110468 115796 110532
rect 115860 110530 115866 110532
rect 116025 110530 116091 110533
rect 115860 110528 116091 110530
rect 115860 110472 116030 110528
rect 116086 110472 116091 110528
rect 115860 110470 116091 110472
rect 115860 110468 115866 110470
rect 116025 110467 116091 110470
rect 140037 110530 140103 110533
rect 144870 110530 144930 110606
rect 147581 110603 147647 110606
rect 140037 110528 144930 110530
rect 140037 110472 140042 110528
rect 140098 110472 144930 110528
rect 140037 110470 144930 110472
rect 170998 110530 171058 110606
rect 171182 110530 171242 110742
rect 180750 110666 180810 110742
rect 190502 110742 200130 110802
rect 180750 110606 190378 110666
rect 170998 110470 171242 110530
rect 190318 110530 190378 110606
rect 190502 110530 190562 110742
rect 200070 110666 200130 110742
rect 209822 110742 219450 110802
rect 200070 110606 209698 110666
rect 190318 110470 190562 110530
rect 209638 110530 209698 110606
rect 209822 110530 209882 110742
rect 219390 110666 219450 110742
rect 229142 110742 238770 110802
rect 219390 110606 229018 110666
rect 209638 110470 209882 110530
rect 228958 110530 229018 110606
rect 229142 110530 229202 110742
rect 238710 110666 238770 110742
rect 248462 110742 258090 110802
rect 238710 110606 248338 110666
rect 228958 110470 229202 110530
rect 248278 110530 248338 110606
rect 248462 110530 248522 110742
rect 258030 110666 258090 110742
rect 267782 110742 277410 110802
rect 258030 110606 267658 110666
rect 248278 110470 248522 110530
rect 267598 110530 267658 110606
rect 267782 110530 267842 110742
rect 277350 110666 277410 110742
rect 287102 110742 296730 110802
rect 277350 110606 286978 110666
rect 267598 110470 267842 110530
rect 286918 110530 286978 110606
rect 287102 110530 287162 110742
rect 296670 110666 296730 110742
rect 306422 110742 316050 110802
rect 296670 110606 306298 110666
rect 286918 110470 287162 110530
rect 306238 110530 306298 110606
rect 306422 110530 306482 110742
rect 315990 110666 316050 110742
rect 325742 110742 335370 110802
rect 315990 110606 325618 110666
rect 306238 110470 306482 110530
rect 325558 110530 325618 110606
rect 325742 110530 325802 110742
rect 335310 110666 335370 110742
rect 345062 110742 354690 110802
rect 335310 110606 344938 110666
rect 325558 110470 325802 110530
rect 344878 110530 344938 110606
rect 345062 110530 345122 110742
rect 354630 110666 354690 110742
rect 364382 110742 374010 110802
rect 354630 110606 364258 110666
rect 344878 110470 345122 110530
rect 364198 110530 364258 110606
rect 364382 110530 364442 110742
rect 373950 110666 374010 110742
rect 383702 110742 393330 110802
rect 373950 110606 383578 110666
rect 364198 110470 364442 110530
rect 383518 110530 383578 110606
rect 383702 110530 383762 110742
rect 393270 110666 393330 110742
rect 403022 110742 412650 110802
rect 393270 110606 402898 110666
rect 383518 110470 383762 110530
rect 402838 110530 402898 110606
rect 403022 110530 403082 110742
rect 412590 110666 412650 110742
rect 422342 110742 431970 110802
rect 412590 110606 422218 110666
rect 402838 110470 403082 110530
rect 422158 110530 422218 110606
rect 422342 110530 422402 110742
rect 431910 110666 431970 110742
rect 441662 110742 451290 110802
rect 431910 110606 441538 110666
rect 422158 110470 422402 110530
rect 441478 110530 441538 110606
rect 441662 110530 441722 110742
rect 451230 110666 451290 110742
rect 460982 110742 470610 110802
rect 451230 110606 460858 110666
rect 441478 110470 441722 110530
rect 460798 110530 460858 110606
rect 460982 110530 461042 110742
rect 470550 110666 470610 110742
rect 480302 110742 489930 110802
rect 470550 110606 480178 110666
rect 460798 110470 461042 110530
rect 480118 110530 480178 110606
rect 480302 110530 480362 110742
rect 489870 110666 489930 110742
rect 499622 110742 509250 110802
rect 489870 110606 499498 110666
rect 480118 110470 480362 110530
rect 499438 110530 499498 110606
rect 499622 110530 499682 110742
rect 509190 110666 509250 110742
rect 518942 110742 528570 110802
rect 509190 110606 518818 110666
rect 499438 110470 499682 110530
rect 518758 110530 518818 110606
rect 518942 110530 519002 110742
rect 528510 110666 528570 110742
rect 538262 110742 547890 110802
rect 528510 110606 538138 110666
rect 518758 110470 519002 110530
rect 538078 110530 538138 110606
rect 538262 110530 538322 110742
rect 547830 110666 547890 110742
rect 557582 110742 567210 110802
rect 547830 110606 557458 110666
rect 538078 110470 538322 110530
rect 557398 110530 557458 110606
rect 557582 110530 557642 110742
rect 567150 110666 567210 110742
rect 583342 110666 583402 111422
rect 583520 111332 584960 111422
rect 567150 110606 576778 110666
rect 557398 110470 557642 110530
rect 576718 110530 576778 110606
rect 576902 110606 583402 110666
rect 576902 110530 576962 110606
rect 576718 110470 576962 110530
rect 140037 110467 140103 110470
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 115790 87410 115796 87412
rect 108806 87350 115796 87410
rect 57094 87212 57100 87276
rect 57164 87274 57170 87276
rect 89621 87274 89687 87277
rect 57164 87214 64890 87274
rect 57164 87212 57170 87214
rect 64830 87138 64890 87214
rect 74582 87272 89687 87274
rect 74582 87216 89626 87272
rect 89682 87216 89687 87272
rect 74582 87214 89687 87216
rect 64830 87078 74458 87138
rect 74398 87002 74458 87078
rect 74582 87002 74642 87214
rect 89621 87211 89687 87214
rect 96521 87274 96587 87277
rect 96521 87272 99298 87274
rect 96521 87216 96526 87272
rect 96582 87216 99298 87272
rect 96521 87214 99298 87216
rect 96521 87211 96587 87214
rect 74398 86942 74642 87002
rect 99238 87002 99298 87214
rect 108806 87138 108866 87350
rect 115790 87348 115796 87350
rect 115860 87348 115866 87412
rect 133822 87348 133828 87412
rect 133892 87410 133898 87412
rect 143441 87410 143507 87413
rect 133892 87408 143507 87410
rect 133892 87352 143446 87408
rect 143502 87352 143507 87408
rect 133892 87350 143507 87352
rect 133892 87348 133898 87350
rect 143441 87347 143507 87350
rect 120809 87274 120875 87277
rect 128169 87274 128235 87277
rect 120809 87272 128235 87274
rect 120809 87216 120814 87272
rect 120870 87216 128174 87272
rect 128230 87216 128235 87272
rect 120809 87214 128235 87216
rect 120809 87211 120875 87214
rect 128169 87211 128235 87214
rect 128353 87274 128419 87277
rect 154481 87274 154547 87277
rect 128353 87272 130394 87274
rect 128353 87216 128358 87272
rect 128414 87216 130394 87272
rect 128353 87214 130394 87216
rect 128353 87211 128419 87214
rect 99422 87078 108866 87138
rect 130334 87138 130394 87214
rect 154481 87272 161490 87274
rect 154481 87216 154486 87272
rect 154542 87216 161490 87272
rect 154481 87214 161490 87216
rect 154481 87211 154547 87214
rect 133822 87138 133828 87140
rect 130334 87078 133828 87138
rect 99422 87002 99482 87078
rect 133822 87076 133828 87078
rect 133892 87076 133898 87140
rect 161430 87138 161490 87214
rect 171182 87214 180810 87274
rect 161430 87078 171058 87138
rect 99238 86942 99482 87002
rect 115790 86940 115796 87004
rect 115860 87002 115866 87004
rect 116025 87002 116091 87005
rect 115860 87000 116091 87002
rect 115860 86944 116030 87000
rect 116086 86944 116091 87000
rect 115860 86942 116091 86944
rect 115860 86940 115866 86942
rect 116025 86939 116091 86942
rect 143441 87002 143507 87005
rect 145557 87002 145623 87005
rect 143441 87000 145623 87002
rect 143441 86944 143446 87000
rect 143502 86944 145562 87000
rect 145618 86944 145623 87000
rect 143441 86942 145623 86944
rect 170998 87002 171058 87078
rect 171182 87002 171242 87214
rect 180750 87138 180810 87214
rect 190502 87214 200130 87274
rect 180750 87078 190378 87138
rect 170998 86942 171242 87002
rect 190318 87002 190378 87078
rect 190502 87002 190562 87214
rect 200070 87138 200130 87214
rect 209822 87214 219450 87274
rect 200070 87078 209698 87138
rect 190318 86942 190562 87002
rect 209638 87002 209698 87078
rect 209822 87002 209882 87214
rect 219390 87138 219450 87214
rect 229142 87214 238770 87274
rect 219390 87078 229018 87138
rect 209638 86942 209882 87002
rect 228958 87002 229018 87078
rect 229142 87002 229202 87214
rect 238710 87138 238770 87214
rect 248462 87214 258090 87274
rect 238710 87078 248338 87138
rect 228958 86942 229202 87002
rect 248278 87002 248338 87078
rect 248462 87002 248522 87214
rect 258030 87138 258090 87214
rect 267782 87214 277410 87274
rect 258030 87078 267658 87138
rect 248278 86942 248522 87002
rect 267598 87002 267658 87078
rect 267782 87002 267842 87214
rect 277350 87138 277410 87214
rect 287102 87214 296730 87274
rect 277350 87078 286978 87138
rect 267598 86942 267842 87002
rect 286918 87002 286978 87078
rect 287102 87002 287162 87214
rect 296670 87138 296730 87214
rect 306422 87214 316050 87274
rect 296670 87078 306298 87138
rect 286918 86942 287162 87002
rect 306238 87002 306298 87078
rect 306422 87002 306482 87214
rect 315990 87138 316050 87214
rect 325742 87214 335370 87274
rect 315990 87078 325618 87138
rect 306238 86942 306482 87002
rect 325558 87002 325618 87078
rect 325742 87002 325802 87214
rect 335310 87138 335370 87214
rect 345062 87214 354690 87274
rect 335310 87078 344938 87138
rect 325558 86942 325802 87002
rect 344878 87002 344938 87078
rect 345062 87002 345122 87214
rect 354630 87138 354690 87214
rect 364382 87214 374010 87274
rect 354630 87078 364258 87138
rect 344878 86942 345122 87002
rect 364198 87002 364258 87078
rect 364382 87002 364442 87214
rect 373950 87138 374010 87214
rect 383702 87214 393330 87274
rect 373950 87078 383578 87138
rect 364198 86942 364442 87002
rect 383518 87002 383578 87078
rect 383702 87002 383762 87214
rect 393270 87138 393330 87214
rect 403022 87214 412650 87274
rect 393270 87078 402898 87138
rect 383518 86942 383762 87002
rect 402838 87002 402898 87078
rect 403022 87002 403082 87214
rect 412590 87138 412650 87214
rect 422342 87214 431970 87274
rect 412590 87078 422218 87138
rect 402838 86942 403082 87002
rect 422158 87002 422218 87078
rect 422342 87002 422402 87214
rect 431910 87138 431970 87214
rect 441662 87214 451290 87274
rect 431910 87078 441538 87138
rect 422158 86942 422402 87002
rect 441478 87002 441538 87078
rect 441662 87002 441722 87214
rect 451230 87138 451290 87214
rect 460982 87214 470610 87274
rect 451230 87078 460858 87138
rect 441478 86942 441722 87002
rect 460798 87002 460858 87078
rect 460982 87002 461042 87214
rect 470550 87138 470610 87214
rect 480302 87214 489930 87274
rect 470550 87078 480178 87138
rect 460798 86942 461042 87002
rect 480118 87002 480178 87078
rect 480302 87002 480362 87214
rect 489870 87138 489930 87214
rect 499622 87214 509250 87274
rect 489870 87078 499498 87138
rect 480118 86942 480362 87002
rect 499438 87002 499498 87078
rect 499622 87002 499682 87214
rect 509190 87138 509250 87214
rect 518942 87214 528570 87274
rect 509190 87078 518818 87138
rect 499438 86942 499682 87002
rect 518758 87002 518818 87078
rect 518942 87002 519002 87214
rect 528510 87138 528570 87214
rect 538262 87214 547890 87274
rect 528510 87078 538138 87138
rect 518758 86942 519002 87002
rect 538078 87002 538138 87078
rect 538262 87002 538322 87214
rect 547830 87138 547890 87214
rect 557582 87214 567210 87274
rect 547830 87078 557458 87138
rect 538078 86942 538322 87002
rect 557398 87002 557458 87078
rect 557582 87002 557642 87214
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 557398 86942 557642 87002
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 143441 86939 143507 86942
rect 145557 86939 145623 86942
rect -960 78978 480 79068
rect 3417 78978 3483 78981
rect -960 78976 3483 78978
rect -960 78920 3422 78976
rect 3478 78920 3483 78976
rect -960 78918 3483 78920
rect -960 78828 480 78918
rect 3417 78915 3483 78918
rect 125542 76468 125548 76532
rect 125612 76530 125618 76532
rect 135161 76530 135227 76533
rect 125612 76528 135227 76530
rect 125612 76472 135166 76528
rect 135222 76472 135227 76528
rect 125612 76470 135227 76472
rect 125612 76468 125618 76470
rect 135161 76467 135227 76470
rect 115790 76394 115796 76396
rect 108806 76334 115796 76394
rect 57278 76196 57284 76260
rect 57348 76258 57354 76260
rect 89621 76258 89687 76261
rect 57348 76198 64890 76258
rect 57348 76196 57354 76198
rect 64830 76122 64890 76198
rect 74582 76256 89687 76258
rect 74582 76200 89626 76256
rect 89682 76200 89687 76256
rect 74582 76198 89687 76200
rect 64830 76062 74458 76122
rect 74398 75986 74458 76062
rect 74582 75986 74642 76198
rect 89621 76195 89687 76198
rect 96521 76258 96587 76261
rect 96521 76256 99298 76258
rect 96521 76200 96526 76256
rect 96582 76200 99298 76256
rect 96521 76198 99298 76200
rect 96521 76195 96587 76198
rect 74398 75926 74642 75986
rect 99238 75986 99298 76198
rect 108806 76122 108866 76334
rect 115790 76332 115796 76334
rect 115860 76332 115866 76396
rect 140037 76394 140103 76397
rect 135302 76392 140103 76394
rect 135302 76336 140042 76392
rect 140098 76336 140103 76392
rect 135302 76334 140103 76336
rect 118785 76258 118851 76261
rect 125542 76258 125548 76260
rect 118785 76256 125548 76258
rect 118785 76200 118790 76256
rect 118846 76200 125548 76256
rect 118785 76198 125548 76200
rect 118785 76195 118851 76198
rect 125542 76196 125548 76198
rect 125612 76196 125618 76260
rect 99422 76062 108866 76122
rect 135161 76122 135227 76125
rect 135302 76122 135362 76334
rect 140037 76331 140103 76334
rect 154481 76258 154547 76261
rect 583520 76258 584960 76348
rect 154481 76256 161490 76258
rect 154481 76200 154486 76256
rect 154542 76200 161490 76256
rect 154481 76198 161490 76200
rect 154481 76195 154547 76198
rect 147581 76122 147647 76125
rect 135161 76120 135362 76122
rect 135161 76064 135166 76120
rect 135222 76064 135362 76120
rect 135161 76062 135362 76064
rect 144870 76120 147647 76122
rect 144870 76064 147586 76120
rect 147642 76064 147647 76120
rect 144870 76062 147647 76064
rect 161430 76122 161490 76198
rect 171182 76198 180810 76258
rect 161430 76062 171058 76122
rect 99422 75986 99482 76062
rect 135161 76059 135227 76062
rect 99238 75926 99482 75986
rect 115790 75924 115796 75988
rect 115860 75986 115866 75988
rect 116025 75986 116091 75989
rect 115860 75984 116091 75986
rect 115860 75928 116030 75984
rect 116086 75928 116091 75984
rect 115860 75926 116091 75928
rect 115860 75924 115866 75926
rect 116025 75923 116091 75926
rect 140037 75986 140103 75989
rect 144870 75986 144930 76062
rect 147581 76059 147647 76062
rect 140037 75984 144930 75986
rect 140037 75928 140042 75984
rect 140098 75928 144930 75984
rect 140037 75926 144930 75928
rect 170998 75986 171058 76062
rect 171182 75986 171242 76198
rect 180750 76122 180810 76198
rect 190502 76198 200130 76258
rect 180750 76062 190378 76122
rect 170998 75926 171242 75986
rect 190318 75986 190378 76062
rect 190502 75986 190562 76198
rect 200070 76122 200130 76198
rect 209822 76198 219450 76258
rect 200070 76062 209698 76122
rect 190318 75926 190562 75986
rect 209638 75986 209698 76062
rect 209822 75986 209882 76198
rect 219390 76122 219450 76198
rect 229142 76198 238770 76258
rect 219390 76062 229018 76122
rect 209638 75926 209882 75986
rect 228958 75986 229018 76062
rect 229142 75986 229202 76198
rect 238710 76122 238770 76198
rect 248462 76198 258090 76258
rect 238710 76062 248338 76122
rect 228958 75926 229202 75986
rect 248278 75986 248338 76062
rect 248462 75986 248522 76198
rect 258030 76122 258090 76198
rect 267782 76198 277410 76258
rect 258030 76062 267658 76122
rect 248278 75926 248522 75986
rect 267598 75986 267658 76062
rect 267782 75986 267842 76198
rect 277350 76122 277410 76198
rect 287102 76198 296730 76258
rect 277350 76062 286978 76122
rect 267598 75926 267842 75986
rect 286918 75986 286978 76062
rect 287102 75986 287162 76198
rect 296670 76122 296730 76198
rect 306422 76198 316050 76258
rect 296670 76062 306298 76122
rect 286918 75926 287162 75986
rect 306238 75986 306298 76062
rect 306422 75986 306482 76198
rect 315990 76122 316050 76198
rect 325742 76198 335370 76258
rect 315990 76062 325618 76122
rect 306238 75926 306482 75986
rect 325558 75986 325618 76062
rect 325742 75986 325802 76198
rect 335310 76122 335370 76198
rect 345062 76198 354690 76258
rect 335310 76062 344938 76122
rect 325558 75926 325802 75986
rect 344878 75986 344938 76062
rect 345062 75986 345122 76198
rect 354630 76122 354690 76198
rect 364382 76198 374010 76258
rect 354630 76062 364258 76122
rect 344878 75926 345122 75986
rect 364198 75986 364258 76062
rect 364382 75986 364442 76198
rect 373950 76122 374010 76198
rect 383702 76198 393330 76258
rect 373950 76062 383578 76122
rect 364198 75926 364442 75986
rect 383518 75986 383578 76062
rect 383702 75986 383762 76198
rect 393270 76122 393330 76198
rect 403022 76198 412650 76258
rect 393270 76062 402898 76122
rect 383518 75926 383762 75986
rect 402838 75986 402898 76062
rect 403022 75986 403082 76198
rect 412590 76122 412650 76198
rect 422342 76198 431970 76258
rect 412590 76062 422218 76122
rect 402838 75926 403082 75986
rect 422158 75986 422218 76062
rect 422342 75986 422402 76198
rect 431910 76122 431970 76198
rect 441662 76198 451290 76258
rect 431910 76062 441538 76122
rect 422158 75926 422402 75986
rect 441478 75986 441538 76062
rect 441662 75986 441722 76198
rect 451230 76122 451290 76198
rect 460982 76198 470610 76258
rect 451230 76062 460858 76122
rect 441478 75926 441722 75986
rect 460798 75986 460858 76062
rect 460982 75986 461042 76198
rect 470550 76122 470610 76198
rect 480302 76198 489930 76258
rect 470550 76062 480178 76122
rect 460798 75926 461042 75986
rect 480118 75986 480178 76062
rect 480302 75986 480362 76198
rect 489870 76122 489930 76198
rect 499622 76198 509250 76258
rect 489870 76062 499498 76122
rect 480118 75926 480362 75986
rect 499438 75986 499498 76062
rect 499622 75986 499682 76198
rect 509190 76122 509250 76198
rect 518942 76198 528570 76258
rect 509190 76062 518818 76122
rect 499438 75926 499682 75986
rect 518758 75986 518818 76062
rect 518942 75986 519002 76198
rect 528510 76122 528570 76198
rect 538262 76198 547890 76258
rect 528510 76062 538138 76122
rect 518758 75926 519002 75986
rect 538078 75986 538138 76062
rect 538262 75986 538322 76198
rect 547830 76122 547890 76198
rect 557582 76198 567210 76258
rect 547830 76062 557458 76122
rect 538078 75926 538322 75986
rect 557398 75986 557458 76062
rect 557582 75986 557642 76198
rect 567150 76122 567210 76198
rect 583342 76198 584960 76258
rect 583342 76122 583402 76198
rect 567150 76062 576778 76122
rect 557398 75926 557642 75986
rect 576718 75986 576778 76062
rect 576902 76062 583402 76122
rect 583520 76108 584960 76198
rect 576902 75986 576962 76062
rect 576718 75926 576962 75986
rect 140037 75923 140103 75926
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect 583520 64562 584960 64652
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 583342 64502 584960 64562
rect 125542 64092 125548 64156
rect 125612 64154 125618 64156
rect 135161 64154 135227 64157
rect 125612 64152 135227 64154
rect 125612 64096 135166 64152
rect 135222 64096 135227 64152
rect 125612 64094 135227 64096
rect 125612 64092 125618 64094
rect 135161 64091 135227 64094
rect 115790 64018 115796 64020
rect 108806 63958 115796 64018
rect 57462 63820 57468 63884
rect 57532 63882 57538 63884
rect 88885 63882 88951 63885
rect 57532 63822 64890 63882
rect 57532 63820 57538 63822
rect 64830 63746 64890 63822
rect 74582 63880 88951 63882
rect 74582 63824 88890 63880
rect 88946 63824 88951 63880
rect 74582 63822 88951 63824
rect 64830 63686 74458 63746
rect 74398 63610 74458 63686
rect 74582 63610 74642 63822
rect 88885 63819 88951 63822
rect 96521 63882 96587 63885
rect 96521 63880 99298 63882
rect 96521 63824 96526 63880
rect 96582 63824 99298 63880
rect 96521 63822 99298 63824
rect 96521 63819 96587 63822
rect 74398 63550 74642 63610
rect 99238 63610 99298 63822
rect 108806 63746 108866 63958
rect 115790 63956 115796 63958
rect 115860 63956 115866 64020
rect 140037 64018 140103 64021
rect 135302 64016 140103 64018
rect 135302 63960 140042 64016
rect 140098 63960 140103 64016
rect 135302 63958 140103 63960
rect 118785 63882 118851 63885
rect 125542 63882 125548 63884
rect 118785 63880 125548 63882
rect 118785 63824 118790 63880
rect 118846 63824 125548 63880
rect 118785 63822 125548 63824
rect 118785 63819 118851 63822
rect 125542 63820 125548 63822
rect 125612 63820 125618 63884
rect 99422 63686 108866 63746
rect 135161 63746 135227 63749
rect 135302 63746 135362 63958
rect 140037 63955 140103 63958
rect 154481 63882 154547 63885
rect 154481 63880 161490 63882
rect 154481 63824 154486 63880
rect 154542 63824 161490 63880
rect 154481 63822 161490 63824
rect 154481 63819 154547 63822
rect 147581 63746 147647 63749
rect 135161 63744 135362 63746
rect 135161 63688 135166 63744
rect 135222 63688 135362 63744
rect 135161 63686 135362 63688
rect 144870 63744 147647 63746
rect 144870 63688 147586 63744
rect 147642 63688 147647 63744
rect 144870 63686 147647 63688
rect 161430 63746 161490 63822
rect 171182 63822 180810 63882
rect 161430 63686 171058 63746
rect 99422 63610 99482 63686
rect 135161 63683 135227 63686
rect 99238 63550 99482 63610
rect 115790 63548 115796 63612
rect 115860 63610 115866 63612
rect 116025 63610 116091 63613
rect 115860 63608 116091 63610
rect 115860 63552 116030 63608
rect 116086 63552 116091 63608
rect 115860 63550 116091 63552
rect 115860 63548 115866 63550
rect 116025 63547 116091 63550
rect 140037 63610 140103 63613
rect 144870 63610 144930 63686
rect 147581 63683 147647 63686
rect 140037 63608 144930 63610
rect 140037 63552 140042 63608
rect 140098 63552 144930 63608
rect 140037 63550 144930 63552
rect 170998 63610 171058 63686
rect 171182 63610 171242 63822
rect 180750 63746 180810 63822
rect 190502 63822 200130 63882
rect 180750 63686 190378 63746
rect 170998 63550 171242 63610
rect 190318 63610 190378 63686
rect 190502 63610 190562 63822
rect 200070 63746 200130 63822
rect 209822 63822 219450 63882
rect 200070 63686 209698 63746
rect 190318 63550 190562 63610
rect 209638 63610 209698 63686
rect 209822 63610 209882 63822
rect 219390 63746 219450 63822
rect 229142 63822 238770 63882
rect 219390 63686 229018 63746
rect 209638 63550 209882 63610
rect 228958 63610 229018 63686
rect 229142 63610 229202 63822
rect 238710 63746 238770 63822
rect 248462 63822 258090 63882
rect 238710 63686 248338 63746
rect 228958 63550 229202 63610
rect 248278 63610 248338 63686
rect 248462 63610 248522 63822
rect 258030 63746 258090 63822
rect 267782 63822 277410 63882
rect 258030 63686 267658 63746
rect 248278 63550 248522 63610
rect 267598 63610 267658 63686
rect 267782 63610 267842 63822
rect 277350 63746 277410 63822
rect 287102 63822 296730 63882
rect 277350 63686 286978 63746
rect 267598 63550 267842 63610
rect 286918 63610 286978 63686
rect 287102 63610 287162 63822
rect 296670 63746 296730 63822
rect 306422 63822 316050 63882
rect 296670 63686 306298 63746
rect 286918 63550 287162 63610
rect 306238 63610 306298 63686
rect 306422 63610 306482 63822
rect 315990 63746 316050 63822
rect 325742 63822 335370 63882
rect 315990 63686 325618 63746
rect 306238 63550 306482 63610
rect 325558 63610 325618 63686
rect 325742 63610 325802 63822
rect 335310 63746 335370 63822
rect 345062 63822 354690 63882
rect 335310 63686 344938 63746
rect 325558 63550 325802 63610
rect 344878 63610 344938 63686
rect 345062 63610 345122 63822
rect 354630 63746 354690 63822
rect 364382 63822 374010 63882
rect 354630 63686 364258 63746
rect 344878 63550 345122 63610
rect 364198 63610 364258 63686
rect 364382 63610 364442 63822
rect 373950 63746 374010 63822
rect 383702 63822 393330 63882
rect 373950 63686 383578 63746
rect 364198 63550 364442 63610
rect 383518 63610 383578 63686
rect 383702 63610 383762 63822
rect 393270 63746 393330 63822
rect 403022 63822 412650 63882
rect 393270 63686 402898 63746
rect 383518 63550 383762 63610
rect 402838 63610 402898 63686
rect 403022 63610 403082 63822
rect 412590 63746 412650 63822
rect 422342 63822 431970 63882
rect 412590 63686 422218 63746
rect 402838 63550 403082 63610
rect 422158 63610 422218 63686
rect 422342 63610 422402 63822
rect 431910 63746 431970 63822
rect 441662 63822 451290 63882
rect 431910 63686 441538 63746
rect 422158 63550 422402 63610
rect 441478 63610 441538 63686
rect 441662 63610 441722 63822
rect 451230 63746 451290 63822
rect 460982 63822 470610 63882
rect 451230 63686 460858 63746
rect 441478 63550 441722 63610
rect 460798 63610 460858 63686
rect 460982 63610 461042 63822
rect 470550 63746 470610 63822
rect 480302 63822 489930 63882
rect 470550 63686 480178 63746
rect 460798 63550 461042 63610
rect 480118 63610 480178 63686
rect 480302 63610 480362 63822
rect 489870 63746 489930 63822
rect 499622 63822 509250 63882
rect 489870 63686 499498 63746
rect 480118 63550 480362 63610
rect 499438 63610 499498 63686
rect 499622 63610 499682 63822
rect 509190 63746 509250 63822
rect 518942 63822 528570 63882
rect 509190 63686 518818 63746
rect 499438 63550 499682 63610
rect 518758 63610 518818 63686
rect 518942 63610 519002 63822
rect 528510 63746 528570 63822
rect 538262 63822 547890 63882
rect 528510 63686 538138 63746
rect 518758 63550 519002 63610
rect 538078 63610 538138 63686
rect 538262 63610 538322 63822
rect 547830 63746 547890 63822
rect 557582 63822 567210 63882
rect 547830 63686 557458 63746
rect 538078 63550 538322 63610
rect 557398 63610 557458 63686
rect 557582 63610 557642 63822
rect 567150 63746 567210 63822
rect 583342 63746 583402 64502
rect 583520 64412 584960 64502
rect 567150 63686 576778 63746
rect 557398 63550 557642 63610
rect 576718 63610 576778 63686
rect 576902 63686 583402 63746
rect 576902 63610 576962 63686
rect 576718 63550 576962 63610
rect 140037 63547 140103 63550
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 125542 40564 125548 40628
rect 125612 40626 125618 40628
rect 135161 40626 135227 40629
rect 125612 40624 135227 40626
rect 125612 40568 135166 40624
rect 135222 40568 135227 40624
rect 125612 40566 135227 40568
rect 125612 40564 125618 40566
rect 135161 40563 135227 40566
rect 115790 40490 115796 40492
rect 108806 40430 115796 40490
rect 57646 40292 57652 40356
rect 57716 40354 57722 40356
rect 88885 40354 88951 40357
rect 57716 40294 64890 40354
rect 57716 40292 57722 40294
rect 64830 40218 64890 40294
rect 74582 40352 88951 40354
rect 74582 40296 88890 40352
rect 88946 40296 88951 40352
rect 74582 40294 88951 40296
rect 64830 40158 74458 40218
rect 74398 40082 74458 40158
rect 74582 40082 74642 40294
rect 88885 40291 88951 40294
rect 96521 40354 96587 40357
rect 96521 40352 99298 40354
rect 96521 40296 96526 40352
rect 96582 40296 99298 40352
rect 96521 40294 99298 40296
rect 96521 40291 96587 40294
rect 74398 40022 74642 40082
rect 99238 40082 99298 40294
rect 108806 40218 108866 40430
rect 115790 40428 115796 40430
rect 115860 40428 115866 40492
rect 140037 40490 140103 40493
rect 135302 40488 140103 40490
rect 135302 40432 140042 40488
rect 140098 40432 140103 40488
rect 135302 40430 140103 40432
rect 118785 40354 118851 40357
rect 125542 40354 125548 40356
rect 118785 40352 125548 40354
rect 118785 40296 118790 40352
rect 118846 40296 125548 40352
rect 118785 40294 125548 40296
rect 118785 40291 118851 40294
rect 125542 40292 125548 40294
rect 125612 40292 125618 40356
rect 99422 40158 108866 40218
rect 135161 40218 135227 40221
rect 135302 40218 135362 40430
rect 140037 40427 140103 40430
rect 154481 40354 154547 40357
rect 154481 40352 161490 40354
rect 154481 40296 154486 40352
rect 154542 40296 161490 40352
rect 154481 40294 161490 40296
rect 154481 40291 154547 40294
rect 147581 40218 147647 40221
rect 135161 40216 135362 40218
rect 135161 40160 135166 40216
rect 135222 40160 135362 40216
rect 135161 40158 135362 40160
rect 144870 40216 147647 40218
rect 144870 40160 147586 40216
rect 147642 40160 147647 40216
rect 144870 40158 147647 40160
rect 161430 40218 161490 40294
rect 171182 40294 180810 40354
rect 161430 40158 171058 40218
rect 99422 40082 99482 40158
rect 135161 40155 135227 40158
rect 99238 40022 99482 40082
rect 115790 40020 115796 40084
rect 115860 40082 115866 40084
rect 116025 40082 116091 40085
rect 115860 40080 116091 40082
rect 115860 40024 116030 40080
rect 116086 40024 116091 40080
rect 115860 40022 116091 40024
rect 115860 40020 115866 40022
rect 116025 40019 116091 40022
rect 140037 40082 140103 40085
rect 144870 40082 144930 40158
rect 147581 40155 147647 40158
rect 140037 40080 144930 40082
rect 140037 40024 140042 40080
rect 140098 40024 144930 40080
rect 140037 40022 144930 40024
rect 170998 40082 171058 40158
rect 171182 40082 171242 40294
rect 180750 40218 180810 40294
rect 190502 40294 200130 40354
rect 180750 40158 190378 40218
rect 170998 40022 171242 40082
rect 190318 40082 190378 40158
rect 190502 40082 190562 40294
rect 200070 40218 200130 40294
rect 209822 40294 219450 40354
rect 200070 40158 209698 40218
rect 190318 40022 190562 40082
rect 209638 40082 209698 40158
rect 209822 40082 209882 40294
rect 219390 40218 219450 40294
rect 229142 40294 238770 40354
rect 219390 40158 229018 40218
rect 209638 40022 209882 40082
rect 228958 40082 229018 40158
rect 229142 40082 229202 40294
rect 238710 40218 238770 40294
rect 248462 40294 258090 40354
rect 238710 40158 248338 40218
rect 228958 40022 229202 40082
rect 248278 40082 248338 40158
rect 248462 40082 248522 40294
rect 258030 40218 258090 40294
rect 267782 40294 277410 40354
rect 258030 40158 267658 40218
rect 248278 40022 248522 40082
rect 267598 40082 267658 40158
rect 267782 40082 267842 40294
rect 277350 40218 277410 40294
rect 287102 40294 296730 40354
rect 277350 40158 286978 40218
rect 267598 40022 267842 40082
rect 286918 40082 286978 40158
rect 287102 40082 287162 40294
rect 296670 40218 296730 40294
rect 306422 40294 316050 40354
rect 296670 40158 306298 40218
rect 286918 40022 287162 40082
rect 306238 40082 306298 40158
rect 306422 40082 306482 40294
rect 315990 40218 316050 40294
rect 325742 40294 335370 40354
rect 315990 40158 325618 40218
rect 306238 40022 306482 40082
rect 325558 40082 325618 40158
rect 325742 40082 325802 40294
rect 335310 40218 335370 40294
rect 345062 40294 354690 40354
rect 335310 40158 344938 40218
rect 325558 40022 325802 40082
rect 344878 40082 344938 40158
rect 345062 40082 345122 40294
rect 354630 40218 354690 40294
rect 364382 40294 374010 40354
rect 354630 40158 364258 40218
rect 344878 40022 345122 40082
rect 364198 40082 364258 40158
rect 364382 40082 364442 40294
rect 373950 40218 374010 40294
rect 383702 40294 393330 40354
rect 373950 40158 383578 40218
rect 364198 40022 364442 40082
rect 383518 40082 383578 40158
rect 383702 40082 383762 40294
rect 393270 40218 393330 40294
rect 403022 40294 412650 40354
rect 393270 40158 402898 40218
rect 383518 40022 383762 40082
rect 402838 40082 402898 40158
rect 403022 40082 403082 40294
rect 412590 40218 412650 40294
rect 422342 40294 431970 40354
rect 412590 40158 422218 40218
rect 402838 40022 403082 40082
rect 422158 40082 422218 40158
rect 422342 40082 422402 40294
rect 431910 40218 431970 40294
rect 441662 40294 451290 40354
rect 431910 40158 441538 40218
rect 422158 40022 422402 40082
rect 441478 40082 441538 40158
rect 441662 40082 441722 40294
rect 451230 40218 451290 40294
rect 460982 40294 470610 40354
rect 451230 40158 460858 40218
rect 441478 40022 441722 40082
rect 460798 40082 460858 40158
rect 460982 40082 461042 40294
rect 470550 40218 470610 40294
rect 480302 40294 489930 40354
rect 470550 40158 480178 40218
rect 460798 40022 461042 40082
rect 480118 40082 480178 40158
rect 480302 40082 480362 40294
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 480118 40022 480362 40082
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576902 40158 583402 40218
rect 576902 40082 576962 40158
rect 576718 40022 576962 40082
rect 140037 40019 140103 40022
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 115790 29474 115796 29476
rect 108806 29414 115796 29474
rect 56726 29276 56732 29340
rect 56796 29338 56802 29340
rect 89621 29338 89687 29341
rect 56796 29278 64890 29338
rect 56796 29276 56802 29278
rect 64830 29202 64890 29278
rect 74582 29336 89687 29338
rect 74582 29280 89626 29336
rect 89682 29280 89687 29336
rect 74582 29278 89687 29280
rect 64830 29142 74458 29202
rect 74398 29066 74458 29142
rect 74582 29066 74642 29278
rect 89621 29275 89687 29278
rect 96521 29338 96587 29341
rect 96521 29336 99298 29338
rect 96521 29280 96526 29336
rect 96582 29280 99298 29336
rect 96521 29278 99298 29280
rect 96521 29275 96587 29278
rect 74398 29006 74642 29066
rect 99238 29066 99298 29278
rect 108806 29202 108866 29414
rect 115790 29412 115796 29414
rect 115860 29412 115866 29476
rect 133822 29412 133828 29476
rect 133892 29474 133898 29476
rect 143441 29474 143507 29477
rect 133892 29472 143507 29474
rect 133892 29416 143446 29472
rect 143502 29416 143507 29472
rect 133892 29414 143507 29416
rect 133892 29412 133898 29414
rect 143441 29411 143507 29414
rect 120809 29338 120875 29341
rect 128169 29338 128235 29341
rect 120809 29336 128235 29338
rect 120809 29280 120814 29336
rect 120870 29280 128174 29336
rect 128230 29280 128235 29336
rect 120809 29278 128235 29280
rect 120809 29275 120875 29278
rect 128169 29275 128235 29278
rect 128353 29338 128419 29341
rect 154481 29338 154547 29341
rect 583520 29338 584960 29428
rect 128353 29336 130394 29338
rect 128353 29280 128358 29336
rect 128414 29280 130394 29336
rect 128353 29278 130394 29280
rect 128353 29275 128419 29278
rect 99422 29142 108866 29202
rect 130334 29202 130394 29278
rect 154481 29336 161490 29338
rect 154481 29280 154486 29336
rect 154542 29280 161490 29336
rect 154481 29278 161490 29280
rect 154481 29275 154547 29278
rect 133822 29202 133828 29204
rect 130334 29142 133828 29202
rect 99422 29066 99482 29142
rect 133822 29140 133828 29142
rect 133892 29140 133898 29204
rect 161430 29202 161490 29278
rect 171182 29278 180810 29338
rect 161430 29142 171058 29202
rect 99238 29006 99482 29066
rect 115790 29004 115796 29068
rect 115860 29066 115866 29068
rect 116025 29066 116091 29069
rect 115860 29064 116091 29066
rect 115860 29008 116030 29064
rect 116086 29008 116091 29064
rect 115860 29006 116091 29008
rect 115860 29004 115866 29006
rect 116025 29003 116091 29006
rect 143441 29066 143507 29069
rect 145005 29066 145071 29069
rect 143441 29064 145071 29066
rect 143441 29008 143446 29064
rect 143502 29008 145010 29064
rect 145066 29008 145071 29064
rect 143441 29006 145071 29008
rect 170998 29066 171058 29142
rect 171182 29066 171242 29278
rect 180750 29202 180810 29278
rect 190502 29278 200130 29338
rect 180750 29142 190378 29202
rect 170998 29006 171242 29066
rect 190318 29066 190378 29142
rect 190502 29066 190562 29278
rect 200070 29202 200130 29278
rect 209822 29278 219450 29338
rect 200070 29142 209698 29202
rect 190318 29006 190562 29066
rect 209638 29066 209698 29142
rect 209822 29066 209882 29278
rect 219390 29202 219450 29278
rect 229142 29278 238770 29338
rect 219390 29142 229018 29202
rect 209638 29006 209882 29066
rect 228958 29066 229018 29142
rect 229142 29066 229202 29278
rect 238710 29202 238770 29278
rect 248462 29278 258090 29338
rect 238710 29142 248338 29202
rect 228958 29006 229202 29066
rect 248278 29066 248338 29142
rect 248462 29066 248522 29278
rect 258030 29202 258090 29278
rect 267782 29278 277410 29338
rect 258030 29142 267658 29202
rect 248278 29006 248522 29066
rect 267598 29066 267658 29142
rect 267782 29066 267842 29278
rect 277350 29202 277410 29278
rect 287102 29278 296730 29338
rect 277350 29142 286978 29202
rect 267598 29006 267842 29066
rect 286918 29066 286978 29142
rect 287102 29066 287162 29278
rect 296670 29202 296730 29278
rect 306422 29278 316050 29338
rect 296670 29142 306298 29202
rect 286918 29006 287162 29066
rect 306238 29066 306298 29142
rect 306422 29066 306482 29278
rect 315990 29202 316050 29278
rect 325742 29278 335370 29338
rect 315990 29142 325618 29202
rect 306238 29006 306482 29066
rect 325558 29066 325618 29142
rect 325742 29066 325802 29278
rect 335310 29202 335370 29278
rect 345062 29278 354690 29338
rect 335310 29142 344938 29202
rect 325558 29006 325802 29066
rect 344878 29066 344938 29142
rect 345062 29066 345122 29278
rect 354630 29202 354690 29278
rect 364382 29278 374010 29338
rect 354630 29142 364258 29202
rect 344878 29006 345122 29066
rect 364198 29066 364258 29142
rect 364382 29066 364442 29278
rect 373950 29202 374010 29278
rect 383702 29278 393330 29338
rect 373950 29142 383578 29202
rect 364198 29006 364442 29066
rect 383518 29066 383578 29142
rect 383702 29066 383762 29278
rect 393270 29202 393330 29278
rect 403022 29278 412650 29338
rect 393270 29142 402898 29202
rect 383518 29006 383762 29066
rect 402838 29066 402898 29142
rect 403022 29066 403082 29278
rect 412590 29202 412650 29278
rect 422342 29278 431970 29338
rect 412590 29142 422218 29202
rect 402838 29006 403082 29066
rect 422158 29066 422218 29142
rect 422342 29066 422402 29278
rect 431910 29202 431970 29278
rect 441662 29278 451290 29338
rect 431910 29142 441538 29202
rect 422158 29006 422402 29066
rect 441478 29066 441538 29142
rect 441662 29066 441722 29278
rect 451230 29202 451290 29278
rect 460982 29278 470610 29338
rect 451230 29142 460858 29202
rect 441478 29006 441722 29066
rect 460798 29066 460858 29142
rect 460982 29066 461042 29278
rect 470550 29202 470610 29278
rect 480302 29278 489930 29338
rect 470550 29142 480178 29202
rect 460798 29006 461042 29066
rect 480118 29066 480178 29142
rect 480302 29066 480362 29278
rect 489870 29202 489930 29278
rect 499622 29278 509250 29338
rect 489870 29142 499498 29202
rect 480118 29006 480362 29066
rect 499438 29066 499498 29142
rect 499622 29066 499682 29278
rect 509190 29202 509250 29278
rect 518942 29278 528570 29338
rect 509190 29142 518818 29202
rect 499438 29006 499682 29066
rect 518758 29066 518818 29142
rect 518942 29066 519002 29278
rect 528510 29202 528570 29278
rect 538262 29278 547890 29338
rect 528510 29142 538138 29202
rect 518758 29006 519002 29066
rect 538078 29066 538138 29142
rect 538262 29066 538322 29278
rect 547830 29202 547890 29278
rect 557582 29278 567210 29338
rect 547830 29142 557458 29202
rect 538078 29006 538322 29066
rect 557398 29066 557458 29142
rect 557582 29066 557642 29278
rect 567150 29202 567210 29278
rect 583342 29278 584960 29338
rect 583342 29202 583402 29278
rect 567150 29142 576778 29202
rect 557398 29006 557642 29066
rect 576718 29066 576778 29142
rect 576902 29142 583402 29202
rect 583520 29188 584960 29278
rect 576902 29066 576962 29142
rect 576718 29006 576962 29066
rect 143441 29003 143507 29006
rect 145005 29003 145071 29006
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
rect 80237 5266 80303 5269
rect 202873 5266 202939 5269
rect 80237 5264 202939 5266
rect 80237 5208 80242 5264
rect 80298 5208 202878 5264
rect 202934 5208 202939 5264
rect 80237 5206 202939 5208
rect 80237 5203 80303 5206
rect 202873 5203 202939 5206
rect 87321 5130 87387 5133
rect 215293 5130 215359 5133
rect 87321 5128 215359 5130
rect 87321 5072 87326 5128
rect 87382 5072 215298 5128
rect 215354 5072 215359 5128
rect 87321 5070 215359 5072
rect 87321 5067 87387 5070
rect 215293 5067 215359 5070
rect 94497 4994 94563 4997
rect 227713 4994 227779 4997
rect 94497 4992 227779 4994
rect 94497 4936 94502 4992
rect 94558 4936 227718 4992
rect 227774 4936 227779 4992
rect 94497 4934 227779 4936
rect 94497 4931 94563 4934
rect 227713 4931 227779 4934
rect 105169 4858 105235 4861
rect 247033 4858 247099 4861
rect 105169 4856 247099 4858
rect 105169 4800 105174 4856
rect 105230 4800 247038 4856
rect 247094 4800 247099 4856
rect 105169 4798 247099 4800
rect 105169 4795 105235 4798
rect 247033 4795 247099 4798
rect 106273 4042 106339 4045
rect 115657 4042 115723 4045
rect 106273 4040 115723 4042
rect 106273 3984 106278 4040
rect 106334 3984 115662 4040
rect 115718 3984 115723 4040
rect 106273 3982 115723 3984
rect 106273 3979 106339 3982
rect 115657 3979 115723 3982
rect 114645 3906 114711 3909
rect 117313 3906 117379 3909
rect 114645 3904 117379 3906
rect 114645 3848 114650 3904
rect 114706 3848 117318 3904
rect 117374 3848 117379 3904
rect 114645 3846 117379 3848
rect 114645 3843 114711 3846
rect 117313 3843 117379 3846
rect 89713 3770 89779 3773
rect 219433 3770 219499 3773
rect 89713 3768 219499 3770
rect 89713 3712 89718 3768
rect 89774 3712 219438 3768
rect 219494 3712 219499 3768
rect 89713 3710 219499 3712
rect 89713 3707 89779 3710
rect 219433 3707 219499 3710
rect 96889 3634 96955 3637
rect 231853 3634 231919 3637
rect 96889 3632 231919 3634
rect 96889 3576 96894 3632
rect 96950 3576 231858 3632
rect 231914 3576 231919 3632
rect 96889 3574 231919 3576
rect 96889 3571 96955 3574
rect 231853 3571 231919 3574
rect 111149 3498 111215 3501
rect 258073 3498 258139 3501
rect 111149 3496 258139 3498
rect 111149 3440 111154 3496
rect 111210 3440 258078 3496
rect 258134 3440 258139 3496
rect 111149 3438 258139 3440
rect 111149 3435 111215 3438
rect 258073 3435 258139 3438
rect 125409 3362 125475 3365
rect 282913 3362 282979 3365
rect 125409 3360 282979 3362
rect 125409 3304 125414 3360
rect 125470 3304 282918 3360
rect 282974 3304 282979 3360
rect 125409 3302 282979 3304
rect 125409 3299 125475 3302
rect 282913 3299 282979 3302
<< via3 >>
rect 57468 700708 57532 700772
rect 57652 700572 57716 700636
rect 59124 700436 59188 700500
rect 57836 700300 57900 700364
rect 550588 673916 550652 673980
rect 57284 673780 57348 673844
rect 299428 673780 299492 673844
rect 299428 673508 299492 673572
rect 550588 673508 550652 673572
rect 550588 650388 550652 650452
rect 58204 650252 58268 650316
rect 299428 650252 299492 650316
rect 299428 649980 299492 650044
rect 550588 649980 550652 650044
rect 550588 626996 550652 627060
rect 58020 626860 58084 626924
rect 299428 626860 299492 626924
rect 299428 626588 299492 626652
rect 434668 626860 434732 626924
rect 434668 626588 434732 626652
rect 550588 626588 550652 626652
rect 299428 603332 299492 603396
rect 299428 603060 299492 603124
rect 434668 603196 434732 603260
rect 434668 602924 434732 602988
rect 59492 596124 59556 596188
rect 59308 581572 59372 581636
rect 59860 581572 59924 581636
rect 59860 579592 59924 579596
rect 59860 579536 59874 579592
rect 59874 579536 59924 579592
rect 59860 579532 59924 579536
rect 59676 570012 59740 570076
rect 59676 563212 59740 563276
rect 59492 562940 59556 563004
rect 133644 553480 133708 553484
rect 133644 553424 133694 553480
rect 133694 553424 133708 553480
rect 133644 553420 133708 553424
rect 259132 553480 259196 553484
rect 259132 553424 259182 553480
rect 259182 553424 259196 553480
rect 259132 553420 259196 553424
rect 263732 553480 263796 553484
rect 263732 553424 263782 553480
rect 263782 553424 263796 553480
rect 263732 553420 263796 553424
rect 378548 553480 378612 553484
rect 378548 553424 378562 553480
rect 378562 553424 378612 553480
rect 378548 553420 378612 553424
rect 382964 553480 383028 553484
rect 382964 553424 382978 553480
rect 382978 553424 383028 553480
rect 382964 553420 383028 553424
rect 507900 553480 507964 553484
rect 507900 553424 507914 553480
rect 507914 553424 507964 553480
rect 507900 553420 507964 553424
rect 513420 553480 513484 553484
rect 513420 553424 513434 553480
rect 513434 553424 513484 553480
rect 513420 553420 513484 553424
rect 129228 551108 129292 551172
rect 132908 551108 132972 551172
rect 514156 550700 514220 550764
rect 351840 459640 351904 459644
rect 351840 459584 351882 459640
rect 351882 459584 351904 459640
rect 351840 459580 351904 459584
rect 77312 459504 77376 459508
rect 77312 459448 77354 459504
rect 77354 459448 77376 459504
rect 77312 459444 77376 459448
rect 327312 459444 327376 459508
rect 328480 459444 328544 459508
rect 328868 459444 328932 459508
rect 358848 459504 358912 459508
rect 358848 459448 358874 459504
rect 358874 459448 358912 459504
rect 358848 459444 358912 459448
rect 452640 459444 452704 459508
rect 453068 459444 453132 459508
rect 483008 459504 483072 459508
rect 483008 459448 483018 459504
rect 483018 459448 483072 459504
rect 483008 459444 483072 459448
rect 73844 458084 73908 458148
rect 74948 458084 75012 458148
rect 79364 458084 79428 458148
rect 81940 458144 82004 458148
rect 81940 458088 81954 458144
rect 81954 458088 82004 458144
rect 81940 458084 82004 458088
rect 82860 458144 82924 458148
rect 82860 458088 82874 458144
rect 82874 458088 82924 458144
rect 82860 458084 82924 458088
rect 84148 458144 84212 458148
rect 84148 458088 84198 458144
rect 84198 458088 84212 458144
rect 84148 458084 84212 458088
rect 85436 458144 85500 458148
rect 85436 458088 85486 458144
rect 85486 458088 85500 458144
rect 85436 458084 85500 458088
rect 86356 458144 86420 458148
rect 86356 458088 86370 458144
rect 86370 458088 86420 458144
rect 86356 458084 86420 458088
rect 87828 458144 87892 458148
rect 87828 458088 87878 458144
rect 87878 458088 87892 458144
rect 87828 458084 87892 458088
rect 88932 458084 88996 458148
rect 90220 458144 90284 458148
rect 90220 458088 90234 458144
rect 90234 458088 90284 458144
rect 90220 458084 90284 458088
rect 91324 458084 91388 458148
rect 92428 458144 92492 458148
rect 92428 458088 92478 458144
rect 92478 458088 92492 458144
rect 92428 458084 92492 458088
rect 93532 458144 93596 458148
rect 93532 458088 93582 458144
rect 93582 458088 93596 458144
rect 93532 458084 93596 458088
rect 94820 458144 94884 458148
rect 94820 458088 94834 458144
rect 94834 458088 94884 458144
rect 94820 458084 94884 458088
rect 95740 458144 95804 458148
rect 95740 458088 95790 458144
rect 95790 458088 95804 458144
rect 95740 458084 95804 458088
rect 97212 458144 97276 458148
rect 97212 458088 97226 458144
rect 97226 458088 97276 458144
rect 97212 458084 97276 458088
rect 98316 458084 98380 458148
rect 99420 458144 99484 458148
rect 99420 458088 99470 458144
rect 99470 458088 99484 458144
rect 99420 458084 99484 458088
rect 100156 458084 100220 458148
rect 101996 458144 102060 458148
rect 101996 458088 102010 458144
rect 102010 458088 102060 458144
rect 101996 458084 102060 458088
rect 102732 458144 102796 458148
rect 102732 458088 102782 458144
rect 102782 458088 102796 458144
rect 102732 458084 102796 458088
rect 103100 458084 103164 458148
rect 104204 458144 104268 458148
rect 104204 458088 104254 458144
rect 104254 458088 104268 458144
rect 104204 458084 104268 458088
rect 104756 458144 104820 458148
rect 104756 458088 104806 458144
rect 104806 458088 104820 458144
rect 104756 458084 104820 458088
rect 105308 458144 105372 458148
rect 105308 458088 105358 458144
rect 105358 458088 105372 458144
rect 105308 458084 105372 458088
rect 105492 458084 105556 458148
rect 107148 458084 107212 458148
rect 108804 458144 108868 458148
rect 108804 458088 108818 458144
rect 108818 458088 108868 458144
rect 108804 458084 108868 458088
rect 108988 458084 109052 458148
rect 193812 458144 193876 458148
rect 193812 458088 193862 458144
rect 193862 458088 193876 458144
rect 193812 458084 193876 458088
rect 200252 458144 200316 458148
rect 200252 458088 200266 458144
rect 200266 458088 200316 458144
rect 200252 458084 200316 458088
rect 210556 458144 210620 458148
rect 210556 458088 210570 458144
rect 210570 458088 210620 458144
rect 210556 458084 210620 458088
rect 212028 458084 212092 458148
rect 213132 458144 213196 458148
rect 213132 458088 213146 458144
rect 213146 458088 213196 458144
rect 213132 458084 213196 458088
rect 214052 458144 214116 458148
rect 214052 458088 214066 458144
rect 214066 458088 214116 458144
rect 214052 458084 214116 458088
rect 215340 458144 215404 458148
rect 215340 458088 215354 458144
rect 215354 458088 215404 458144
rect 215340 458084 215404 458088
rect 216628 458144 216692 458148
rect 216628 458088 216678 458144
rect 216678 458088 216692 458144
rect 216628 458084 216692 458088
rect 217548 458144 217612 458148
rect 217548 458088 217598 458144
rect 217598 458088 217612 458144
rect 217548 458084 217612 458088
rect 218836 458144 218900 458148
rect 218836 458088 218886 458144
rect 218886 458088 218900 458144
rect 218836 458084 218900 458088
rect 220124 458144 220188 458148
rect 220124 458088 220174 458144
rect 220174 458088 220188 458144
rect 220124 458084 220188 458088
rect 221412 458144 221476 458148
rect 221412 458088 221426 458144
rect 221426 458088 221476 458144
rect 221412 458084 221476 458088
rect 222516 458144 222580 458148
rect 222516 458088 222566 458144
rect 222566 458088 222580 458144
rect 222516 458084 222580 458088
rect 223620 458144 223684 458148
rect 223620 458088 223670 458144
rect 223670 458088 223684 458144
rect 223620 458084 223684 458088
rect 224356 458144 224420 458148
rect 224356 458088 224370 458144
rect 224370 458088 224420 458144
rect 224356 458084 224420 458088
rect 225828 458144 225892 458148
rect 225828 458088 225878 458144
rect 225878 458088 225892 458144
rect 225828 458084 225892 458088
rect 227116 458144 227180 458148
rect 227116 458088 227166 458144
rect 227166 458088 227180 458144
rect 227116 458084 227180 458088
rect 228404 458144 228468 458148
rect 228404 458088 228418 458144
rect 228418 458088 228468 458144
rect 228404 458084 228468 458088
rect 229508 458144 229572 458148
rect 229508 458088 229558 458144
rect 229558 458088 229572 458144
rect 229508 458084 229572 458088
rect 232820 458084 232884 458148
rect 233556 458084 233620 458148
rect 313780 458144 313844 458148
rect 313780 458088 313794 458144
rect 313794 458088 313844 458144
rect 313780 458084 313844 458088
rect 322796 458084 322860 458148
rect 323900 458084 323964 458148
rect 326292 458084 326356 458148
rect 327396 458084 327460 458148
rect 328868 458084 328932 458148
rect 330892 458084 330956 458148
rect 331812 458144 331876 458148
rect 331812 458088 331862 458144
rect 331862 458088 331876 458144
rect 331812 458084 331876 458088
rect 333100 458144 333164 458148
rect 333100 458088 333150 458144
rect 333150 458088 333164 458144
rect 333100 458084 333164 458088
rect 334020 458144 334084 458148
rect 334020 458088 334070 458144
rect 334070 458088 334084 458144
rect 334020 458084 334084 458088
rect 335308 458144 335372 458148
rect 335308 458088 335358 458144
rect 335358 458088 335372 458144
rect 335308 458084 335372 458088
rect 336596 458144 336660 458148
rect 336596 458088 336610 458144
rect 336610 458088 336660 458144
rect 336596 458084 336660 458088
rect 337700 458084 337764 458148
rect 338988 458144 339052 458148
rect 338988 458088 339038 458144
rect 339038 458088 339052 458144
rect 338988 458084 339052 458088
rect 339908 458144 339972 458148
rect 339908 458088 339922 458144
rect 339922 458088 339972 458144
rect 339908 458084 339972 458088
rect 341196 458144 341260 458148
rect 341196 458088 341246 458144
rect 341246 458088 341260 458144
rect 341196 458084 341260 458088
rect 342668 458084 342732 458148
rect 343956 458084 344020 458148
rect 344692 458144 344756 458148
rect 344692 458088 344742 458144
rect 344742 458088 344756 458144
rect 344692 458084 344756 458088
rect 346164 458084 346228 458148
rect 347268 458084 347332 458148
rect 348372 458084 348436 458148
rect 349660 458084 349724 458148
rect 352972 458084 353036 458148
rect 353524 458084 353588 458148
rect 461716 458144 461780 458148
rect 461716 458088 461766 458144
rect 461766 458088 461780 458144
rect 461716 458084 461780 458088
rect 463004 458144 463068 458148
rect 463004 458088 463054 458144
rect 463054 458088 463068 458144
rect 463004 458084 463068 458088
rect 464292 458084 464356 458148
rect 465212 458144 465276 458148
rect 465212 458088 465226 458144
rect 465226 458088 465276 458144
rect 465212 458084 465276 458088
rect 468708 458144 468772 458148
rect 468708 458088 468758 458144
rect 468758 458088 468772 458144
rect 468708 458084 468772 458088
rect 469996 458144 470060 458148
rect 469996 458088 470010 458144
rect 470010 458088 470060 458144
rect 469996 458084 470060 458088
rect 471284 458084 471348 458148
rect 472204 458144 472268 458148
rect 472204 458088 472254 458144
rect 472254 458088 472268 458144
rect 472204 458084 472268 458088
rect 473492 458144 473556 458148
rect 473492 458088 473506 458144
rect 473506 458088 473556 458144
rect 473492 458084 473556 458088
rect 474780 458144 474844 458148
rect 474780 458088 474830 458144
rect 474830 458088 474844 458144
rect 474780 458084 474844 458088
rect 475516 458144 475580 458148
rect 475516 458088 475530 458144
rect 475530 458088 475580 458144
rect 475516 458084 475580 458088
rect 476988 458144 477052 458148
rect 476988 458088 477002 458144
rect 477002 458088 477052 458144
rect 476988 458084 477052 458088
rect 478276 458144 478340 458148
rect 478276 458088 478326 458144
rect 478326 458088 478340 458144
rect 478276 458084 478340 458088
rect 479380 458144 479444 458148
rect 479380 458088 479430 458144
rect 479430 458088 479444 458144
rect 479380 458084 479444 458088
rect 483060 458144 483124 458148
rect 483060 458088 483074 458144
rect 483074 458088 483124 458144
rect 483060 458084 483124 458088
rect 484164 458084 484228 458148
rect 485452 458084 485516 458148
rect 80652 457948 80716 458012
rect 100524 458008 100588 458012
rect 100524 457952 100574 458008
rect 100574 457952 100588 458008
rect 100524 457948 100588 457952
rect 101444 457948 101508 458012
rect 106412 457948 106476 458012
rect 107700 458008 107764 458012
rect 107700 457952 107714 458008
rect 107714 457952 107764 458008
rect 107700 457948 107764 457952
rect 108436 457948 108500 458012
rect 197492 457948 197556 458012
rect 199148 457948 199212 458012
rect 207060 457948 207124 458012
rect 234660 458008 234724 458012
rect 234660 457952 234674 458008
rect 234674 457952 234724 458008
rect 234660 457948 234724 457952
rect 322612 457948 322676 458012
rect 323532 458008 323596 458012
rect 323532 457952 323582 458008
rect 323582 457952 323596 458008
rect 323532 457948 323596 457952
rect 329604 457948 329668 458012
rect 342484 458008 342548 458012
rect 342484 457952 342534 458008
rect 342534 457952 342548 458008
rect 342484 457948 342548 457952
rect 343588 457948 343652 458012
rect 345980 458008 346044 458012
rect 345980 457952 345994 458008
rect 345994 457952 346044 458008
rect 345980 457948 346044 457952
rect 346900 458008 346964 458012
rect 346900 457952 346914 458008
rect 346914 457952 346964 458008
rect 346900 457948 346964 457952
rect 348188 458008 348252 458012
rect 348188 457952 348238 458008
rect 348238 457952 348252 458008
rect 348188 457948 348252 457952
rect 349476 457948 349540 458012
rect 350580 458008 350644 458012
rect 350580 457952 350594 458008
rect 350594 457952 350644 458008
rect 350580 457948 350644 457952
rect 356468 457948 356532 458012
rect 443132 457948 443196 458012
rect 459508 457948 459572 458012
rect 467788 457948 467852 458012
rect 480668 457948 480732 458012
rect 487660 457948 487724 458012
rect 78444 457812 78508 457876
rect 101812 457872 101876 457876
rect 101812 457816 101862 457872
rect 101862 457816 101876 457872
rect 101812 457812 101876 457816
rect 231900 457872 231964 457876
rect 231900 457816 231914 457872
rect 231914 457816 231964 457872
rect 231900 457812 231964 457816
rect 236500 457812 236564 457876
rect 317460 457872 317524 457876
rect 317460 457816 317474 457872
rect 317474 457816 317524 457872
rect 317460 457812 317524 457816
rect 324820 457812 324884 457876
rect 326108 457812 326172 457876
rect 330524 457872 330588 457876
rect 330524 457816 330538 457872
rect 330538 457816 330588 457872
rect 330524 457812 330588 457816
rect 355180 457812 355244 457876
rect 458588 457812 458652 457876
rect 466500 457812 466564 457876
rect 479564 457812 479628 457876
rect 480852 457812 480916 457876
rect 484716 457812 484780 457876
rect 72740 457676 72804 457740
rect 201540 457736 201604 457740
rect 201540 457680 201554 457736
rect 201554 457680 201604 457736
rect 201540 457676 201604 457680
rect 209636 457736 209700 457740
rect 209636 457680 209686 457736
rect 209686 457680 209700 457736
rect 209636 457676 209700 457680
rect 237420 457736 237484 457740
rect 237420 457680 237434 457736
rect 237434 457680 237484 457736
rect 237420 457676 237484 457680
rect 238892 457676 238956 457740
rect 331996 457676 332060 457740
rect 344876 457676 344940 457740
rect 357388 457736 357452 457740
rect 357388 457680 357438 457736
rect 357438 457680 357452 457736
rect 357388 457676 357452 457680
rect 460796 457676 460860 457740
rect 481588 457736 481652 457740
rect 481588 457680 481638 457736
rect 481638 457680 481652 457736
rect 481588 457676 481652 457680
rect 486004 457676 486068 457740
rect 488580 457736 488644 457740
rect 488580 457680 488594 457736
rect 488594 457680 488644 457736
rect 488580 457676 488644 457680
rect 63724 457600 63788 457604
rect 63724 457544 63738 457600
rect 63738 457544 63788 457600
rect 63724 457540 63788 457544
rect 75868 457540 75932 457604
rect 196756 457540 196820 457604
rect 230612 457540 230676 457604
rect 457484 457540 457548 457604
rect 459692 457540 459756 457604
rect 487844 457540 487908 457604
rect 74212 457404 74276 457468
rect 76236 457404 76300 457468
rect 208532 457404 208596 457468
rect 216260 457404 216324 457468
rect 453804 457404 453868 457468
rect 455092 457404 455156 457468
rect 483612 457404 483676 457468
rect 486556 457404 486620 457468
rect 488948 457404 489012 457468
rect 206140 457268 206204 457332
rect 329788 457328 329852 457332
rect 329788 457272 329838 457328
rect 329838 457272 329852 457328
rect 329788 457268 329852 457272
rect 477172 457268 477236 457332
rect 478460 457268 478524 457332
rect 72924 457132 72988 457196
rect 77340 457192 77404 457196
rect 77340 457136 77354 457192
rect 77354 457136 77404 457192
rect 77340 457132 77404 457136
rect 95004 457132 95068 457196
rect 98500 457132 98564 457196
rect 202460 457132 202524 457196
rect 202644 457132 202708 457196
rect 206324 457132 206388 457196
rect 209820 457132 209884 457196
rect 214420 457132 214484 457196
rect 216812 457132 216876 457196
rect 220308 457132 220372 457196
rect 325004 457132 325068 457196
rect 328500 457192 328564 457196
rect 328500 457136 328514 457192
rect 328514 457136 328564 457192
rect 328500 457132 328564 457136
rect 335492 457132 335556 457196
rect 341380 457132 341444 457196
rect 354260 457132 354324 457196
rect 451412 457132 451476 457196
rect 454724 457192 454788 457196
rect 454724 457136 454738 457192
rect 454738 457136 454788 457192
rect 454724 457132 454788 457136
rect 458220 457132 458284 457196
rect 462084 457132 462148 457196
rect 469076 457132 469140 457196
rect 472572 457132 472636 457196
rect 476068 457132 476132 457196
rect 481956 457132 482020 457196
rect 70164 457056 70228 457060
rect 70164 457000 70214 457056
rect 70214 457000 70228 457056
rect 70164 456996 70228 457000
rect 75132 456996 75196 457060
rect 78628 456996 78692 457060
rect 93164 456996 93228 457060
rect 205036 456996 205100 457060
rect 225644 456996 225708 457060
rect 232636 456996 232700 457060
rect 320956 456996 321020 457060
rect 337884 456996 337948 457060
rect 353156 456996 353220 457060
rect 447916 456996 447980 457060
rect 456012 457056 456076 457060
rect 456012 457000 456062 457056
rect 456062 457000 456076 457056
rect 456012 456996 456076 457000
rect 66852 456860 66916 456924
rect 67956 456860 68020 456924
rect 69796 456860 69860 456924
rect 71452 456860 71516 456924
rect 79732 456860 79796 456924
rect 80836 456860 80900 456924
rect 82124 456860 82188 456924
rect 83228 456860 83292 456924
rect 84332 456860 84396 456924
rect 85620 456860 85684 456924
rect 86724 456860 86788 456924
rect 88012 456860 88076 456924
rect 89116 456860 89180 456924
rect 90588 456860 90652 456924
rect 91508 456860 91572 456924
rect 93716 456920 93780 456924
rect 93716 456864 93730 456920
rect 93730 456864 93780 456920
rect 93716 456860 93780 456864
rect 96108 456860 96172 456924
rect 97764 456860 97828 456924
rect 203748 456860 203812 456924
rect 203932 456860 203996 456924
rect 205404 456860 205468 456924
rect 207428 456860 207492 456924
rect 209268 456860 209332 456924
rect 210924 456860 210988 456924
rect 212396 456920 212460 456924
rect 212396 456864 212446 456920
rect 212446 456864 212460 456920
rect 212396 456860 212460 456864
rect 213316 456860 213380 456924
rect 217916 456920 217980 456924
rect 217916 456864 217930 456920
rect 217930 456864 217980 456920
rect 217916 456860 217980 456864
rect 219204 456860 219268 456924
rect 221964 456860 222028 456924
rect 223252 456860 223316 456924
rect 223804 456860 223868 456924
rect 226196 456920 226260 456924
rect 226196 456864 226210 456920
rect 226210 456864 226260 456920
rect 226196 456860 226260 456864
rect 227300 456860 227364 456924
rect 228956 456920 229020 456924
rect 228956 456864 229006 456920
rect 229006 456864 229020 456920
rect 228956 456860 229020 456864
rect 229692 456860 229756 456924
rect 230796 456860 230860 456924
rect 233004 456860 233068 456924
rect 234292 456860 234356 456924
rect 235764 456860 235828 456924
rect 236684 456860 236748 456924
rect 237788 456860 237852 456924
rect 239628 456860 239692 456924
rect 316172 456860 316236 456924
rect 319116 456860 319180 456924
rect 320220 456920 320284 456924
rect 320220 456864 320234 456920
rect 320234 456864 320284 456920
rect 320220 456860 320284 456864
rect 333284 456860 333348 456924
rect 334388 456860 334452 456924
rect 336780 456920 336844 456924
rect 336780 456864 336794 456920
rect 336794 456864 336844 456920
rect 336780 456860 336844 456864
rect 339172 456860 339236 456924
rect 340276 456860 340340 456924
rect 350948 456860 351012 456924
rect 351868 456920 351932 456924
rect 351868 456864 351918 456920
rect 351918 456864 351932 456920
rect 351868 456860 351932 456864
rect 355364 456860 355428 456924
rect 356652 456860 356716 456924
rect 357756 456860 357820 456924
rect 358860 456920 358924 456924
rect 358860 456864 358874 456920
rect 358874 456864 358924 456920
rect 358860 456860 358924 456864
rect 446812 456860 446876 456924
rect 448468 456860 448532 456924
rect 450308 456860 450372 456924
rect 452700 456920 452764 456924
rect 452700 456864 452750 456920
rect 452750 456864 452764 456920
rect 452700 456860 452764 456864
rect 453068 456860 453132 456924
rect 453620 456860 453684 456924
rect 456196 456860 456260 456924
rect 457300 456860 457364 456924
rect 460980 456920 461044 456924
rect 460980 456864 460994 456920
rect 460994 456864 461044 456920
rect 460980 456860 461044 456864
rect 463188 456860 463252 456924
rect 464476 456860 464540 456924
rect 465580 456860 465644 456924
rect 466684 456860 466748 456924
rect 467972 456860 468036 456924
rect 470180 456860 470244 456924
rect 471468 456860 471532 456924
rect 473676 456860 473740 456924
rect 474964 456860 475028 456924
rect 56916 439588 56980 439652
rect 57100 439452 57164 439516
rect 58756 439316 58820 439380
rect 56732 387772 56796 387836
rect 57468 306308 57532 306372
rect 57652 302092 57716 302156
rect 57836 299916 57900 299980
rect 59124 297876 59188 297940
rect 56916 295700 56980 295764
rect 58756 291484 58820 291548
rect 57284 289444 57348 289508
rect 58204 285228 58268 285292
rect 58020 283052 58084 283116
rect 58940 278836 59004 278900
rect 56732 274620 56796 274684
rect 57100 266188 57164 266252
rect 57652 249460 57716 249524
rect 57836 247284 57900 247348
rect 56916 213556 56980 213620
rect 57284 211516 57348 211580
rect 57100 209340 57164 209404
rect 57468 207300 57532 207364
rect 56732 205124 56796 205188
rect 57652 204988 57716 205052
rect 57652 203084 57716 203148
rect 57836 200636 57900 200700
rect 125548 111012 125612 111076
rect 56916 110740 56980 110804
rect 115796 110876 115860 110940
rect 125548 110740 125612 110804
rect 115796 110468 115860 110532
rect 57100 87212 57164 87276
rect 115796 87348 115860 87412
rect 133828 87348 133892 87412
rect 133828 87076 133892 87140
rect 115796 86940 115860 87004
rect 125548 76468 125612 76532
rect 57284 76196 57348 76260
rect 115796 76332 115860 76396
rect 125548 76196 125612 76260
rect 115796 75924 115860 75988
rect 125548 64092 125612 64156
rect 57468 63820 57532 63884
rect 115796 63956 115860 64020
rect 125548 63820 125612 63884
rect 115796 63548 115860 63612
rect 125548 40564 125612 40628
rect 57652 40292 57716 40356
rect 115796 40428 115860 40492
rect 125548 40292 125612 40356
rect 115796 40020 115860 40084
rect 56732 29276 56796 29340
rect 115796 29412 115860 29476
rect 133828 29412 133892 29476
rect 133828 29140 133892 29204
rect 115796 29004 115860 29068
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 57467 700772 57533 700773
rect 57467 700708 57468 700772
rect 57532 700708 57533 700772
rect 57467 700707 57533 700708
rect 57283 673844 57349 673845
rect 57283 673780 57284 673844
rect 57348 673780 57349 673844
rect 57283 673779 57349 673780
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 56915 439652 56981 439653
rect 56915 439588 56916 439652
rect 56980 439588 56981 439652
rect 56915 439587 56981 439588
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 56731 387836 56797 387837
rect 56731 387772 56732 387836
rect 56796 387772 56797 387836
rect 56731 387771 56797 387772
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 56734 274685 56794 387771
rect 56918 295765 56978 439587
rect 57099 439516 57165 439517
rect 57099 439452 57100 439516
rect 57164 439452 57165 439516
rect 57099 439451 57165 439452
rect 56915 295764 56981 295765
rect 56915 295700 56916 295764
rect 56980 295700 56981 295764
rect 56915 295699 56981 295700
rect 56731 274684 56797 274685
rect 56731 274620 56732 274684
rect 56796 274620 56797 274684
rect 56731 274619 56797 274620
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 57102 266253 57162 439451
rect 57286 289509 57346 673779
rect 57470 306373 57530 700707
rect 57651 700636 57717 700637
rect 57651 700572 57652 700636
rect 57716 700572 57717 700636
rect 57651 700571 57717 700572
rect 57467 306372 57533 306373
rect 57467 306308 57468 306372
rect 57532 306308 57533 306372
rect 57467 306307 57533 306308
rect 57654 302157 57714 700571
rect 57835 700364 57901 700365
rect 57835 700300 57836 700364
rect 57900 700300 57901 700364
rect 57835 700299 57901 700300
rect 57651 302156 57717 302157
rect 57651 302092 57652 302156
rect 57716 302092 57717 302156
rect 57651 302091 57717 302092
rect 57838 299981 57898 700299
rect 58404 672054 59004 707102
rect 59123 700500 59189 700501
rect 59123 700436 59124 700500
rect 59188 700436 59189 700500
rect 59123 700435 59189 700436
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58203 650316 58269 650317
rect 58203 650252 58204 650316
rect 58268 650252 58269 650316
rect 58203 650251 58269 650252
rect 58019 626924 58085 626925
rect 58019 626860 58020 626924
rect 58084 626860 58085 626924
rect 58019 626859 58085 626860
rect 57835 299980 57901 299981
rect 57835 299916 57836 299980
rect 57900 299916 57901 299980
rect 57835 299915 57901 299916
rect 57283 289508 57349 289509
rect 57283 289444 57284 289508
rect 57348 289444 57349 289508
rect 57283 289443 57349 289444
rect 58022 283117 58082 626859
rect 58206 285293 58266 650251
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 59126 596730 59186 700435
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 59126 596670 59370 596730
rect 59310 581637 59370 596670
rect 59491 596188 59557 596189
rect 59491 596124 59492 596188
rect 59556 596124 59557 596188
rect 59491 596123 59557 596124
rect 59307 581636 59373 581637
rect 59307 581572 59308 581636
rect 59372 581572 59373 581636
rect 59307 581571 59373 581572
rect 59494 577690 59554 596123
rect 59859 581636 59925 581637
rect 59859 581572 59860 581636
rect 59924 581572 59925 581636
rect 59859 581571 59925 581572
rect 59862 579597 59922 581571
rect 59859 579596 59925 579597
rect 59859 579532 59860 579596
rect 59924 579532 59925 579596
rect 59859 579531 59925 579532
rect 59310 577630 59554 577690
rect 59310 572930 59370 577630
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 554247 59004 563498
rect 59126 572870 59370 572930
rect 59126 553210 59186 572870
rect 59675 570076 59741 570077
rect 59675 570012 59676 570076
rect 59740 570012 59741 570076
rect 59675 570011 59741 570012
rect 59678 563277 59738 570011
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 59675 563276 59741 563277
rect 59675 563212 59676 563276
rect 59740 563212 59741 563276
rect 59675 563211 59741 563212
rect 59491 563004 59557 563005
rect 59491 562940 59492 563004
rect 59556 562940 59557 563004
rect 59491 562939 59557 562940
rect 59494 553210 59554 562939
rect 62004 554247 62604 567098
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 554247 66204 570698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 554247 73404 577898
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 554247 77004 581498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 554247 80604 585098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 554247 84204 588698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 554247 91404 559898
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 554247 95004 563498
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 554247 98604 567098
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 554247 102204 570698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 554247 109404 577898
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 554247 113004 581498
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 554247 116604 585098
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 554247 120204 588698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 554247 127404 559898
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 554247 131004 563498
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 554247 134604 567098
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 554247 138204 570698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 133643 553484 133709 553485
rect 133643 553420 133644 553484
rect 133708 553420 133709 553484
rect 133643 553419 133709 553420
rect 58942 553150 59186 553210
rect 59310 553150 59554 553210
rect 58942 457330 59002 553150
rect 59310 552530 59370 553150
rect 59126 552470 59370 552530
rect 59126 458010 59186 552470
rect 133646 551850 133706 553419
rect 133573 551790 133706 551850
rect 129227 551172 129293 551173
rect 129227 551170 129228 551172
rect 128608 551110 129228 551170
rect 129227 551108 129228 551110
rect 129292 551108 129293 551172
rect 129227 551107 129293 551108
rect 132907 551172 132973 551173
rect 132907 551108 132908 551172
rect 132972 551170 132973 551172
rect 133573 551170 133633 551790
rect 132972 551140 133633 551170
rect 132972 551110 133603 551140
rect 132972 551108 132973 551110
rect 132907 551107 132973 551108
rect 136494 546054 136814 546076
rect 136494 545818 136536 546054
rect 136772 545818 136814 546054
rect 136494 545734 136814 545818
rect 136494 545498 136536 545734
rect 136772 545498 136814 545734
rect 136494 545476 136814 545498
rect 136494 542454 136814 542476
rect 136494 542218 136536 542454
rect 136772 542218 136814 542454
rect 136494 542134 136814 542218
rect 136494 541898 136536 542134
rect 136772 541898 136814 542134
rect 136494 541876 136814 541898
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 136938 535254 137262 535276
rect 136938 535018 136982 535254
rect 137218 535018 137262 535254
rect 136938 534934 137262 535018
rect 136938 534698 136982 534934
rect 137218 534698 137262 534934
rect 136938 534676 137262 534698
rect 136938 531654 137262 531676
rect 136938 531418 136982 531654
rect 137218 531418 137262 531654
rect 136938 531334 137262 531418
rect 136938 531098 136982 531334
rect 137218 531098 137262 531334
rect 136938 531076 137262 531098
rect 136938 528054 137262 528076
rect 136938 527818 136982 528054
rect 137218 527818 137262 528054
rect 136938 527734 137262 527818
rect 136938 527498 136982 527734
rect 137218 527498 137262 527734
rect 136938 527476 137262 527498
rect 136938 524454 137262 524476
rect 136938 524218 136982 524454
rect 137218 524218 137262 524454
rect 136938 524134 137262 524218
rect 136938 523898 136982 524134
rect 137218 523898 137262 524134
rect 136938 523876 137262 523898
rect 136494 517254 136814 517276
rect 136494 517018 136536 517254
rect 136772 517018 136814 517254
rect 136494 516934 136814 517018
rect 136494 516698 136536 516934
rect 136772 516698 136814 516934
rect 136494 516676 136814 516698
rect 136494 513654 136814 513676
rect 136494 513418 136536 513654
rect 136772 513418 136814 513654
rect 136494 513334 136814 513418
rect 136494 513098 136536 513334
rect 136772 513098 136814 513334
rect 136494 513076 136814 513098
rect 136494 510054 136814 510076
rect 136494 509818 136536 510054
rect 136772 509818 136814 510054
rect 136494 509734 136814 509818
rect 136494 509498 136536 509734
rect 136772 509498 136814 509734
rect 136494 509476 136814 509498
rect 136494 506454 136814 506476
rect 136494 506218 136536 506454
rect 136772 506218 136814 506454
rect 136494 506134 136814 506218
rect 136494 505898 136536 506134
rect 136772 505898 136814 506134
rect 136494 505876 136814 505898
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 136938 499254 137262 499276
rect 136938 499018 136982 499254
rect 137218 499018 137262 499254
rect 136938 498934 137262 499018
rect 136938 498698 136982 498934
rect 137218 498698 137262 498934
rect 136938 498676 137262 498698
rect 136938 495654 137262 495676
rect 136938 495418 136982 495654
rect 137218 495418 137262 495654
rect 136938 495334 137262 495418
rect 136938 495098 136982 495334
rect 137218 495098 137262 495334
rect 136938 495076 137262 495098
rect 136938 492054 137262 492076
rect 136938 491818 136982 492054
rect 137218 491818 137262 492054
rect 136938 491734 137262 491818
rect 136938 491498 136982 491734
rect 137218 491498 137262 491734
rect 136938 491476 137262 491498
rect 136938 488454 137262 488476
rect 136938 488218 136982 488454
rect 137218 488218 137262 488454
rect 136938 488134 137262 488218
rect 136938 487898 136982 488134
rect 137218 487898 137262 488134
rect 136938 487876 137262 487898
rect 136494 481254 136814 481276
rect 136494 481018 136536 481254
rect 136772 481018 136814 481254
rect 136494 480934 136814 481018
rect 136494 480698 136536 480934
rect 136772 480698 136814 480934
rect 136494 480676 136814 480698
rect 136494 477654 136814 477676
rect 136494 477418 136536 477654
rect 136772 477418 136814 477654
rect 136494 477334 136814 477418
rect 136494 477098 136536 477334
rect 136772 477098 136814 477334
rect 136494 477076 136814 477098
rect 136494 474054 136814 474076
rect 136494 473818 136536 474054
rect 136772 473818 136814 474054
rect 136494 473734 136814 473818
rect 136494 473498 136536 473734
rect 136772 473498 136814 473734
rect 136494 473476 136814 473498
rect 136494 470454 136814 470476
rect 136494 470218 136536 470454
rect 136772 470218 136814 470454
rect 136494 470134 136814 470218
rect 136494 469898 136536 470134
rect 136772 469898 136814 470134
rect 136494 469876 136814 469898
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 136938 463254 137262 463276
rect 136938 463018 136982 463254
rect 137218 463018 137262 463254
rect 136938 462934 137262 463018
rect 136938 462698 136982 462934
rect 137218 462698 137262 462934
rect 136938 462676 137262 462698
rect 73964 460670 74274 460730
rect 69168 460330 69858 460390
rect 63803 459370 63863 460020
rect 63726 459310 63863 459370
rect 66802 459370 66862 460020
rect 67970 459370 68030 460020
rect 66802 459310 66914 459370
rect 59126 457950 59370 458010
rect 58942 457270 59186 457330
rect 58404 456054 59004 457000
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 443000 59004 455498
rect 59126 439650 59186 457270
rect 58942 439590 59186 439650
rect 58755 439380 58821 439381
rect 58755 439316 58756 439380
rect 58820 439316 58821 439380
rect 58755 439315 58821 439316
rect 58758 291549 58818 439315
rect 58755 291548 58821 291549
rect 58755 291484 58756 291548
rect 58820 291484 58821 291548
rect 58755 291483 58821 291484
rect 58203 285292 58269 285293
rect 58203 285228 58204 285292
rect 58268 285228 58269 285292
rect 58203 285227 58269 285228
rect 58019 283116 58085 283117
rect 58019 283052 58020 283116
rect 58084 283052 58085 283116
rect 58019 283051 58085 283052
rect 58942 278901 59002 439590
rect 59310 438970 59370 457950
rect 63726 457605 63786 459310
rect 63723 457604 63789 457605
rect 63723 457540 63724 457604
rect 63788 457540 63789 457604
rect 63723 457539 63789 457540
rect 62004 443000 62604 457000
rect 65604 443000 66204 457000
rect 66854 456925 66914 459310
rect 67958 459310 68030 459370
rect 67958 456925 68018 459310
rect 69798 456925 69858 460330
rect 70166 460330 70336 460390
rect 72796 460330 72986 460390
rect 70166 457061 70226 460330
rect 71474 459370 71534 460020
rect 71454 459310 71534 459370
rect 72642 459370 72702 460020
rect 72642 459310 72802 459370
rect 70163 457060 70229 457061
rect 70163 456996 70164 457060
rect 70228 456996 70229 457060
rect 70163 456995 70229 456996
rect 71454 456925 71514 459310
rect 72742 457741 72802 459310
rect 72739 457740 72805 457741
rect 72739 457676 72740 457740
rect 72804 457676 72805 457740
rect 72739 457675 72805 457676
rect 72926 457197 72986 460330
rect 73810 459370 73870 460020
rect 73810 459310 73906 459370
rect 73846 458149 73906 459310
rect 73843 458148 73909 458149
rect 73843 458084 73844 458148
rect 73908 458084 73909 458148
rect 73843 458083 73909 458084
rect 74214 457469 74274 460670
rect 75870 460670 76176 460730
rect 79366 460670 79680 460730
rect 82862 460670 83184 460730
rect 86358 460670 86688 460730
rect 95742 460670 96032 460730
rect 102734 460670 103040 460730
rect 74978 459370 75038 460020
rect 74950 459310 75038 459370
rect 75102 459370 75162 460020
rect 75102 459310 75194 459370
rect 74950 458149 75010 459310
rect 74947 458148 75013 458149
rect 74947 458084 74948 458148
rect 75012 458084 75013 458148
rect 74947 458083 75013 458084
rect 74211 457468 74277 457469
rect 74211 457404 74212 457468
rect 74276 457404 74277 457468
rect 74211 457403 74277 457404
rect 72923 457196 72989 457197
rect 72923 457132 72924 457196
rect 72988 457132 72989 457196
rect 72923 457131 72989 457132
rect 75134 457061 75194 459310
rect 75870 457605 75930 460670
rect 76270 459370 76330 460020
rect 77314 459509 77374 460020
rect 77311 459508 77377 459509
rect 77311 459444 77312 459508
rect 77376 459444 77377 459508
rect 77311 459443 77377 459444
rect 77438 459370 77498 460020
rect 78482 459370 78542 460020
rect 76238 459310 76330 459370
rect 77342 459310 77498 459370
rect 78446 459310 78542 459370
rect 75867 457604 75933 457605
rect 75867 457540 75868 457604
rect 75932 457540 75933 457604
rect 75867 457539 75933 457540
rect 76238 457469 76298 459310
rect 76235 457468 76301 457469
rect 76235 457404 76236 457468
rect 76300 457404 76301 457468
rect 76235 457403 76301 457404
rect 77342 457197 77402 459310
rect 78446 457877 78506 459310
rect 78443 457876 78509 457877
rect 78443 457812 78444 457876
rect 78508 457812 78509 457876
rect 78443 457811 78509 457812
rect 77339 457196 77405 457197
rect 77339 457132 77340 457196
rect 77404 457132 77405 457196
rect 77339 457131 77405 457132
rect 78630 457061 78690 460390
rect 79366 458149 79426 460670
rect 80654 460330 80848 460390
rect 79774 459370 79834 460020
rect 79734 459310 79834 459370
rect 79363 458148 79429 458149
rect 79363 458084 79364 458148
rect 79428 458084 79429 458148
rect 79363 458083 79429 458084
rect 75131 457060 75197 457061
rect 66851 456924 66917 456925
rect 66851 456860 66852 456924
rect 66916 456860 66917 456924
rect 66851 456859 66917 456860
rect 67955 456924 68021 456925
rect 67955 456860 67956 456924
rect 68020 456860 68021 456924
rect 67955 456859 68021 456860
rect 69795 456924 69861 456925
rect 69795 456860 69796 456924
rect 69860 456860 69861 456924
rect 69795 456859 69861 456860
rect 71451 456924 71517 456925
rect 71451 456860 71452 456924
rect 71516 456860 71517 456924
rect 71451 456859 71517 456860
rect 72804 443000 73404 457000
rect 75131 456996 75132 457060
rect 75196 456996 75197 457060
rect 78627 457060 78693 457061
rect 75131 456995 75197 456996
rect 76404 443000 77004 457000
rect 78627 456996 78628 457060
rect 78692 456996 78693 457060
rect 78627 456995 78693 456996
rect 79734 456925 79794 459310
rect 80654 458013 80714 460330
rect 80942 459370 81002 460020
rect 81986 459370 82046 460020
rect 80838 459310 81002 459370
rect 81942 459310 82046 459370
rect 82110 459370 82170 460020
rect 82110 459310 82186 459370
rect 80651 458012 80717 458013
rect 80651 457948 80652 458012
rect 80716 457948 80717 458012
rect 80651 457947 80717 457948
rect 79731 456924 79797 456925
rect 79731 456860 79732 456924
rect 79796 456860 79797 456924
rect 79731 456859 79797 456860
rect 80004 443000 80604 457000
rect 80838 456925 80898 459310
rect 81942 458149 82002 459310
rect 81939 458148 82005 458149
rect 81939 458084 81940 458148
rect 82004 458084 82005 458148
rect 81939 458083 82005 458084
rect 82126 456925 82186 459310
rect 82862 458149 82922 460670
rect 84150 460330 84352 460390
rect 83278 459370 83338 460020
rect 83230 459310 83338 459370
rect 82859 458148 82925 458149
rect 82859 458084 82860 458148
rect 82924 458084 82925 458148
rect 82859 458083 82925 458084
rect 83230 456925 83290 459310
rect 84150 458149 84210 460330
rect 84446 459370 84506 460020
rect 85490 459370 85550 460020
rect 84334 459310 84506 459370
rect 85438 459310 85550 459370
rect 85614 459370 85674 460020
rect 85614 459310 85682 459370
rect 84147 458148 84213 458149
rect 84147 458084 84148 458148
rect 84212 458084 84213 458148
rect 84147 458083 84213 458084
rect 80835 456924 80901 456925
rect 80835 456860 80836 456924
rect 80900 456860 80901 456924
rect 80835 456859 80901 456860
rect 82123 456924 82189 456925
rect 82123 456860 82124 456924
rect 82188 456860 82189 456924
rect 82123 456859 82189 456860
rect 83227 456924 83293 456925
rect 83227 456860 83228 456924
rect 83292 456860 83293 456924
rect 83227 456859 83293 456860
rect 83604 445254 84204 457000
rect 84334 456925 84394 459310
rect 85438 458149 85498 459310
rect 85435 458148 85501 458149
rect 85435 458084 85436 458148
rect 85500 458084 85501 458148
rect 85435 458083 85501 458084
rect 85622 456925 85682 459310
rect 86358 458149 86418 460670
rect 90316 460330 90650 460390
rect 92652 460330 93226 460390
rect 86782 459370 86842 460020
rect 86726 459310 86842 459370
rect 87826 459370 87886 460020
rect 87950 459370 88010 460020
rect 88994 459370 89054 460020
rect 87826 459310 87890 459370
rect 87950 459310 88074 459370
rect 86355 458148 86421 458149
rect 86355 458084 86356 458148
rect 86420 458084 86421 458148
rect 86355 458083 86421 458084
rect 86726 456925 86786 459310
rect 87830 458149 87890 459310
rect 87827 458148 87893 458149
rect 87827 458084 87828 458148
rect 87892 458084 87893 458148
rect 87827 458083 87893 458084
rect 88014 456925 88074 459310
rect 88934 459310 89054 459370
rect 88934 458149 88994 459310
rect 88931 458148 88997 458149
rect 88931 458084 88932 458148
rect 88996 458084 88997 458148
rect 88931 458083 88997 458084
rect 89118 456925 89178 460020
rect 90162 459370 90222 460020
rect 90162 459310 90282 459370
rect 90222 458149 90282 459310
rect 90219 458148 90285 458149
rect 90219 458084 90220 458148
rect 90284 458084 90285 458148
rect 90219 458083 90285 458084
rect 90590 456925 90650 460330
rect 91330 459370 91390 460020
rect 91326 459310 91390 459370
rect 91454 459370 91514 460020
rect 92498 459370 92558 460020
rect 91454 459310 91570 459370
rect 91326 458149 91386 459310
rect 91323 458148 91389 458149
rect 91323 458084 91324 458148
rect 91388 458084 91389 458148
rect 91323 458083 91389 458084
rect 84331 456924 84397 456925
rect 84331 456860 84332 456924
rect 84396 456860 84397 456924
rect 84331 456859 84397 456860
rect 85619 456924 85685 456925
rect 85619 456860 85620 456924
rect 85684 456860 85685 456924
rect 85619 456859 85685 456860
rect 86723 456924 86789 456925
rect 86723 456860 86724 456924
rect 86788 456860 86789 456924
rect 86723 456859 86789 456860
rect 88011 456924 88077 456925
rect 88011 456860 88012 456924
rect 88076 456860 88077 456924
rect 88011 456859 88077 456860
rect 89115 456924 89181 456925
rect 89115 456860 89116 456924
rect 89180 456860 89181 456924
rect 89115 456859 89181 456860
rect 90587 456924 90653 456925
rect 90587 456860 90588 456924
rect 90652 456860 90653 456924
rect 90587 456859 90653 456860
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 443000 84204 444698
rect 90804 452454 91404 457000
rect 91510 456925 91570 459310
rect 92430 459310 92558 459370
rect 92430 458149 92490 459310
rect 92427 458148 92493 458149
rect 92427 458084 92428 458148
rect 92492 458084 92493 458148
rect 92427 458083 92493 458084
rect 93166 457061 93226 460330
rect 93534 460330 93696 460390
rect 93534 458149 93594 460330
rect 93790 459370 93850 460020
rect 94834 459370 94894 460020
rect 93718 459310 93850 459370
rect 94822 459310 94894 459370
rect 94958 459370 95018 460020
rect 94958 459310 95066 459370
rect 93531 458148 93597 458149
rect 93531 458084 93532 458148
rect 93596 458084 93597 458148
rect 93531 458083 93597 458084
rect 93163 457060 93229 457061
rect 93163 456996 93164 457060
rect 93228 456996 93229 457060
rect 93163 456995 93229 456996
rect 93718 456925 93778 459310
rect 94822 458149 94882 459310
rect 94819 458148 94885 458149
rect 94819 458084 94820 458148
rect 94884 458084 94885 458148
rect 94819 458083 94885 458084
rect 95006 457197 95066 459310
rect 95742 458149 95802 460670
rect 97324 460330 97826 460390
rect 99660 460330 100218 460390
rect 96126 459370 96186 460020
rect 96110 459310 96186 459370
rect 97170 459370 97230 460020
rect 97170 459310 97274 459370
rect 95739 458148 95805 458149
rect 95739 458084 95740 458148
rect 95804 458084 95805 458148
rect 95739 458083 95805 458084
rect 95003 457196 95069 457197
rect 95003 457132 95004 457196
rect 95068 457132 95069 457196
rect 95003 457131 95069 457132
rect 91507 456924 91573 456925
rect 91507 456860 91508 456924
rect 91572 456860 91573 456924
rect 91507 456859 91573 456860
rect 93715 456924 93781 456925
rect 93715 456860 93716 456924
rect 93780 456860 93781 456924
rect 93715 456859 93781 456860
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 443000 91404 451898
rect 94404 456054 95004 457000
rect 96110 456925 96170 459310
rect 97214 458149 97274 459310
rect 97211 458148 97277 458149
rect 97211 458084 97212 458148
rect 97276 458084 97277 458148
rect 97211 458083 97277 458084
rect 97766 456925 97826 460330
rect 98338 459370 98398 460020
rect 98318 459310 98398 459370
rect 98462 459370 98522 460020
rect 99506 459370 99566 460020
rect 98462 459310 98562 459370
rect 98318 458149 98378 459310
rect 98315 458148 98381 458149
rect 98315 458084 98316 458148
rect 98380 458084 98381 458148
rect 98315 458083 98381 458084
rect 98502 457197 98562 459310
rect 99422 459310 99566 459370
rect 99422 458149 99482 459310
rect 100158 458149 100218 460330
rect 100526 460330 100704 460390
rect 100828 460330 101506 460390
rect 99419 458148 99485 458149
rect 99419 458084 99420 458148
rect 99484 458084 99485 458148
rect 99419 458083 99485 458084
rect 100155 458148 100221 458149
rect 100155 458084 100156 458148
rect 100220 458084 100221 458148
rect 100155 458083 100221 458084
rect 100526 458013 100586 460330
rect 101446 458013 101506 460330
rect 101842 459370 101902 460020
rect 101814 459310 101902 459370
rect 101966 459370 102026 460020
rect 101966 459310 102058 459370
rect 100523 458012 100589 458013
rect 100523 457948 100524 458012
rect 100588 457948 100589 458012
rect 100523 457947 100589 457948
rect 101443 458012 101509 458013
rect 101443 457948 101444 458012
rect 101508 457948 101509 458012
rect 101443 457947 101509 457948
rect 101814 457877 101874 459310
rect 101998 458149 102058 459310
rect 102734 458149 102794 460670
rect 104332 460330 104818 460390
rect 106668 460330 107210 460390
rect 107836 460330 108498 460390
rect 103134 459370 103194 460020
rect 103102 459310 103194 459370
rect 104178 459370 104238 460020
rect 104178 459310 104266 459370
rect 103102 458149 103162 459310
rect 104206 458149 104266 459310
rect 104758 458149 104818 460330
rect 105346 459370 105406 460020
rect 105310 459310 105406 459370
rect 105470 459370 105530 460020
rect 106514 459370 106574 460020
rect 105470 459310 105554 459370
rect 105310 458149 105370 459310
rect 105494 458149 105554 459310
rect 106414 459310 106574 459370
rect 101995 458148 102061 458149
rect 101995 458084 101996 458148
rect 102060 458084 102061 458148
rect 101995 458083 102061 458084
rect 102731 458148 102797 458149
rect 102731 458084 102732 458148
rect 102796 458084 102797 458148
rect 102731 458083 102797 458084
rect 103099 458148 103165 458149
rect 103099 458084 103100 458148
rect 103164 458084 103165 458148
rect 103099 458083 103165 458084
rect 104203 458148 104269 458149
rect 104203 458084 104204 458148
rect 104268 458084 104269 458148
rect 104203 458083 104269 458084
rect 104755 458148 104821 458149
rect 104755 458084 104756 458148
rect 104820 458084 104821 458148
rect 104755 458083 104821 458084
rect 105307 458148 105373 458149
rect 105307 458084 105308 458148
rect 105372 458084 105373 458148
rect 105307 458083 105373 458084
rect 105491 458148 105557 458149
rect 105491 458084 105492 458148
rect 105556 458084 105557 458148
rect 105491 458083 105557 458084
rect 106414 458013 106474 459310
rect 107150 458149 107210 460330
rect 107682 459370 107742 460020
rect 107682 459310 107762 459370
rect 107147 458148 107213 458149
rect 107147 458084 107148 458148
rect 107212 458084 107213 458148
rect 107147 458083 107213 458084
rect 107702 458013 107762 459310
rect 108438 458013 108498 460330
rect 108850 459370 108910 460020
rect 108806 459310 108910 459370
rect 108806 458149 108866 459310
rect 108990 458149 109050 460390
rect 108803 458148 108869 458149
rect 108803 458084 108804 458148
rect 108868 458084 108869 458148
rect 108803 458083 108869 458084
rect 108987 458148 109053 458149
rect 108987 458084 108988 458148
rect 109052 458084 109053 458148
rect 108987 458083 109053 458084
rect 106411 458012 106477 458013
rect 106411 457948 106412 458012
rect 106476 457948 106477 458012
rect 106411 457947 106477 457948
rect 107699 458012 107765 458013
rect 107699 457948 107700 458012
rect 107764 457948 107765 458012
rect 107699 457947 107765 457948
rect 108435 458012 108501 458013
rect 108435 457948 108436 458012
rect 108500 457948 108501 458012
rect 108435 457947 108501 457948
rect 101811 457876 101877 457877
rect 101811 457812 101812 457876
rect 101876 457812 101877 457876
rect 101811 457811 101877 457812
rect 98499 457196 98565 457197
rect 98499 457132 98500 457196
rect 98564 457132 98565 457196
rect 98499 457131 98565 457132
rect 96107 456924 96173 456925
rect 96107 456860 96108 456924
rect 96172 456860 96173 456924
rect 96107 456859 96173 456860
rect 97763 456924 97829 456925
rect 97763 456860 97764 456924
rect 97828 456860 97829 456924
rect 97763 456859 97829 456860
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 443000 95004 455498
rect 98004 443000 98604 457000
rect 101604 443000 102204 457000
rect 108804 443000 109404 457000
rect 112404 443000 113004 457000
rect 116004 443000 116604 457000
rect 119604 445254 120204 457000
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 443000 120204 444698
rect 126804 452454 127404 457000
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 443000 127404 451898
rect 130404 456054 131004 457000
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 443000 131004 455498
rect 134004 443000 134604 457000
rect 137604 443000 138204 457000
rect 144804 443000 145404 469898
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 443000 149004 473498
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 443000 152604 477098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 443000 156204 444698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 443000 163404 451898
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 443000 167004 455498
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 443000 170604 459098
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 443000 174204 462698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 443000 181404 469898
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 554247 188604 585098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 554247 192204 588698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 554247 199404 559898
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 554247 203004 563498
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 554247 206604 567098
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 554247 210204 570698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 554247 217404 577898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 554247 221004 581498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 554247 224604 585098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 554247 228204 588698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 554247 235404 559898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 554247 239004 563498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 554247 242604 567098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 554247 246204 570698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 554247 253404 577898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 554247 257004 581498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 554247 260604 585098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 554247 264204 588698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 259131 553484 259197 553485
rect 259131 553420 259132 553484
rect 259196 553420 259197 553484
rect 259131 553419 259197 553420
rect 263731 553484 263797 553485
rect 263731 553420 263732 553484
rect 263796 553420 263797 553484
rect 263731 553419 263797 553420
rect 259134 551170 259194 553419
rect 263734 551170 263794 553419
rect 258608 551110 259194 551170
rect 263603 551110 263794 551170
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 266494 546054 266814 546076
rect 266494 545818 266536 546054
rect 266772 545818 266814 546054
rect 266494 545734 266814 545818
rect 266494 545498 266536 545734
rect 266772 545498 266814 545734
rect 266494 545476 266814 545498
rect 266494 542454 266814 542476
rect 266494 542218 266536 542454
rect 266772 542218 266814 542454
rect 266494 542134 266814 542218
rect 266494 541898 266536 542134
rect 266772 541898 266814 542134
rect 266494 541876 266814 541898
rect 266938 535254 267262 535276
rect 266938 535018 266982 535254
rect 267218 535018 267262 535254
rect 266938 534934 267262 535018
rect 266938 534698 266982 534934
rect 267218 534698 267262 534934
rect 266938 534676 267262 534698
rect 266938 531654 267262 531676
rect 266938 531418 266982 531654
rect 267218 531418 267262 531654
rect 266938 531334 267262 531418
rect 266938 531098 266982 531334
rect 267218 531098 267262 531334
rect 266938 531076 267262 531098
rect 266938 528054 267262 528076
rect 266938 527818 266982 528054
rect 267218 527818 267262 528054
rect 266938 527734 267262 527818
rect 266938 527498 266982 527734
rect 267218 527498 267262 527734
rect 266938 527476 267262 527498
rect 266938 524454 267262 524476
rect 266938 524218 266982 524454
rect 267218 524218 267262 524454
rect 266938 524134 267262 524218
rect 266938 523898 266982 524134
rect 267218 523898 267262 524134
rect 266938 523876 267262 523898
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 266494 517254 266814 517276
rect 266494 517018 266536 517254
rect 266772 517018 266814 517254
rect 266494 516934 266814 517018
rect 266494 516698 266536 516934
rect 266772 516698 266814 516934
rect 266494 516676 266814 516698
rect 266494 513654 266814 513676
rect 266494 513418 266536 513654
rect 266772 513418 266814 513654
rect 266494 513334 266814 513418
rect 266494 513098 266536 513334
rect 266772 513098 266814 513334
rect 266494 513076 266814 513098
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 266494 510054 266814 510076
rect 266494 509818 266536 510054
rect 266772 509818 266814 510054
rect 266494 509734 266814 509818
rect 266494 509498 266536 509734
rect 266772 509498 266814 509734
rect 266494 509476 266814 509498
rect 266494 506454 266814 506476
rect 266494 506218 266536 506454
rect 266772 506218 266814 506454
rect 266494 506134 266814 506218
rect 266494 505898 266536 506134
rect 266772 505898 266814 506134
rect 266494 505876 266814 505898
rect 266938 499254 267262 499276
rect 266938 499018 266982 499254
rect 267218 499018 267262 499254
rect 266938 498934 267262 499018
rect 266938 498698 266982 498934
rect 267218 498698 267262 498934
rect 266938 498676 267262 498698
rect 266938 495654 267262 495676
rect 266938 495418 266982 495654
rect 267218 495418 267262 495654
rect 266938 495334 267262 495418
rect 266938 495098 266982 495334
rect 267218 495098 267262 495334
rect 266938 495076 267262 495098
rect 266938 492054 267262 492076
rect 266938 491818 266982 492054
rect 267218 491818 267262 492054
rect 266938 491734 267262 491818
rect 266938 491498 266982 491734
rect 267218 491498 267262 491734
rect 266938 491476 267262 491498
rect 266938 488454 267262 488476
rect 266938 488218 266982 488454
rect 267218 488218 267262 488454
rect 266938 488134 267262 488218
rect 266938 487898 266982 488134
rect 267218 487898 267262 488134
rect 266938 487876 267262 487898
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 266494 481254 266814 481276
rect 266494 481018 266536 481254
rect 266772 481018 266814 481254
rect 266494 480934 266814 481018
rect 266494 480698 266536 480934
rect 266772 480698 266814 480934
rect 266494 480676 266814 480698
rect 266494 477654 266814 477676
rect 266494 477418 266536 477654
rect 266772 477418 266814 477654
rect 266494 477334 266814 477418
rect 266494 477098 266536 477334
rect 266772 477098 266814 477334
rect 266494 477076 266814 477098
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 443000 185004 473498
rect 266494 474054 266814 474076
rect 266494 473818 266536 474054
rect 266772 473818 266814 474054
rect 266494 473734 266814 473818
rect 266494 473498 266536 473734
rect 266772 473498 266814 473734
rect 266494 473476 266814 473498
rect 266494 470454 266814 470476
rect 266494 470218 266536 470454
rect 266772 470218 266814 470454
rect 266494 470134 266814 470218
rect 266494 469898 266536 470134
rect 266772 469898 266814 470134
rect 266494 469876 266814 469898
rect 266938 463254 267262 463276
rect 266938 463018 266982 463254
rect 267218 463018 267262 463254
rect 266938 462934 267262 463018
rect 266938 462698 266982 462934
rect 267218 462698 267262 462934
rect 266938 462676 267262 462698
rect 207062 460670 207344 460730
rect 210558 460670 210848 460730
rect 214054 460670 214352 460730
rect 217550 460670 217856 460730
rect 197494 460330 198000 460390
rect 202462 460330 202672 460390
rect 205132 460330 205466 460390
rect 193803 459370 193863 460020
rect 196802 459370 196862 460020
rect 193803 459310 193874 459370
rect 193814 458149 193874 459310
rect 196758 459310 196862 459370
rect 193811 458148 193877 458149
rect 193811 458084 193812 458148
rect 193876 458084 193877 458148
rect 193811 458083 193877 458084
rect 196758 457605 196818 459310
rect 197494 458013 197554 460330
rect 199138 459370 199198 460020
rect 200306 459370 200366 460020
rect 199138 459310 199210 459370
rect 199150 458013 199210 459310
rect 200254 459310 200366 459370
rect 201474 459370 201534 460020
rect 201474 459310 201602 459370
rect 200254 458149 200314 459310
rect 200251 458148 200317 458149
rect 200251 458084 200252 458148
rect 200316 458084 200317 458148
rect 200251 458083 200317 458084
rect 197491 458012 197557 458013
rect 197491 457948 197492 458012
rect 197556 457948 197557 458012
rect 197491 457947 197557 457948
rect 199147 458012 199213 458013
rect 199147 457948 199148 458012
rect 199212 457948 199213 458012
rect 199147 457947 199213 457948
rect 201542 457741 201602 459310
rect 201539 457740 201605 457741
rect 201539 457676 201540 457740
rect 201604 457676 201605 457740
rect 201539 457675 201605 457676
rect 196755 457604 196821 457605
rect 196755 457540 196756 457604
rect 196820 457540 196821 457604
rect 196755 457539 196821 457540
rect 202462 457197 202522 460330
rect 202766 459370 202826 460020
rect 203810 459370 203870 460020
rect 202646 459310 202826 459370
rect 203750 459310 203870 459370
rect 202646 457197 202706 459310
rect 202459 457196 202525 457197
rect 202459 457132 202460 457196
rect 202524 457132 202525 457196
rect 202459 457131 202525 457132
rect 202643 457196 202709 457197
rect 202643 457132 202644 457196
rect 202708 457132 202709 457196
rect 202643 457131 202709 457132
rect 188004 443000 188604 457000
rect 191604 445254 192204 457000
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 443000 192204 444698
rect 198804 452454 199404 457000
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 443000 199404 451898
rect 202404 456054 203004 457000
rect 203750 456925 203810 459310
rect 203934 456925 203994 460020
rect 204978 459370 205038 460020
rect 204978 459310 205098 459370
rect 205038 457061 205098 459310
rect 205035 457060 205101 457061
rect 205035 456996 205036 457060
rect 205100 456996 205101 457060
rect 205035 456995 205101 456996
rect 205406 456925 205466 460330
rect 206146 459370 206206 460020
rect 206142 459310 206206 459370
rect 206270 459370 206330 460020
rect 206270 459310 206386 459370
rect 206142 457333 206202 459310
rect 206139 457332 206205 457333
rect 206139 457268 206140 457332
rect 206204 457268 206205 457332
rect 206139 457267 206205 457268
rect 206326 457197 206386 459310
rect 207062 458013 207122 460670
rect 208636 460330 209330 460390
rect 207438 459370 207498 460020
rect 207430 459310 207498 459370
rect 208482 459370 208542 460020
rect 208482 459310 208594 459370
rect 207059 458012 207125 458013
rect 207059 457948 207060 458012
rect 207124 457948 207125 458012
rect 207059 457947 207125 457948
rect 206323 457196 206389 457197
rect 206323 457132 206324 457196
rect 206388 457132 206389 457196
rect 206323 457131 206389 457132
rect 203747 456924 203813 456925
rect 203747 456860 203748 456924
rect 203812 456860 203813 456924
rect 203747 456859 203813 456860
rect 203931 456924 203997 456925
rect 203931 456860 203932 456924
rect 203996 456860 203997 456924
rect 203931 456859 203997 456860
rect 205403 456924 205469 456925
rect 205403 456860 205404 456924
rect 205468 456860 205469 456924
rect 205403 456859 205469 456860
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 443000 203004 455498
rect 206004 443000 206604 457000
rect 207430 456925 207490 459310
rect 208534 457469 208594 459310
rect 208531 457468 208597 457469
rect 208531 457404 208532 457468
rect 208596 457404 208597 457468
rect 208531 457403 208597 457404
rect 209270 456925 209330 460330
rect 209650 459370 209710 460020
rect 209638 459310 209710 459370
rect 209774 459370 209834 460020
rect 209774 459310 209882 459370
rect 209638 457741 209698 459310
rect 209635 457740 209701 457741
rect 209635 457676 209636 457740
rect 209700 457676 209701 457740
rect 209635 457675 209701 457676
rect 209822 457197 209882 459310
rect 210558 458149 210618 460670
rect 212140 460330 212458 460390
rect 210942 459370 211002 460020
rect 210926 459310 211002 459370
rect 211986 459370 212046 460020
rect 211986 459310 212090 459370
rect 210555 458148 210621 458149
rect 210555 458084 210556 458148
rect 210620 458084 210621 458148
rect 210555 458083 210621 458084
rect 209819 457196 209885 457197
rect 209819 457132 209820 457196
rect 209884 457132 209885 457196
rect 209819 457131 209885 457132
rect 207427 456924 207493 456925
rect 207427 456860 207428 456924
rect 207492 456860 207493 456924
rect 207427 456859 207493 456860
rect 209267 456924 209333 456925
rect 209267 456860 209268 456924
rect 209332 456860 209333 456924
rect 209267 456859 209333 456860
rect 209604 443000 210204 457000
rect 210926 456925 210986 459310
rect 212030 458149 212090 459310
rect 212027 458148 212093 458149
rect 212027 458084 212028 458148
rect 212092 458084 212093 458148
rect 212027 458083 212093 458084
rect 212398 456925 212458 460330
rect 213154 459370 213214 460020
rect 213134 459310 213214 459370
rect 213278 459370 213338 460020
rect 213278 459310 213378 459370
rect 213134 458149 213194 459310
rect 213131 458148 213197 458149
rect 213131 458084 213132 458148
rect 213196 458084 213197 458148
rect 213131 458083 213197 458084
rect 213318 456925 213378 459310
rect 214054 458149 214114 460670
rect 215342 460330 215520 460390
rect 215644 460330 216322 460390
rect 214446 459370 214506 460020
rect 214422 459310 214506 459370
rect 214051 458148 214117 458149
rect 214051 458084 214052 458148
rect 214116 458084 214117 458148
rect 214051 458083 214117 458084
rect 214422 457197 214482 459310
rect 215342 458149 215402 460330
rect 215339 458148 215405 458149
rect 215339 458084 215340 458148
rect 215404 458084 215405 458148
rect 215339 458083 215405 458084
rect 216262 457469 216322 460330
rect 216658 459370 216718 460020
rect 216630 459310 216718 459370
rect 216782 459370 216842 460020
rect 216782 459310 216874 459370
rect 216630 458149 216690 459310
rect 216627 458148 216693 458149
rect 216627 458084 216628 458148
rect 216692 458084 216693 458148
rect 216627 458083 216693 458084
rect 216259 457468 216325 457469
rect 216259 457404 216260 457468
rect 216324 457404 216325 457468
rect 216259 457403 216325 457404
rect 216814 457197 216874 459310
rect 217550 458149 217610 460670
rect 218838 460330 219024 460390
rect 221484 460330 222026 460390
rect 222652 460330 223314 460390
rect 217950 459370 218010 460020
rect 217918 459310 218010 459370
rect 217547 458148 217613 458149
rect 217547 458084 217548 458148
rect 217612 458084 217613 458148
rect 217547 458083 217613 458084
rect 214419 457196 214485 457197
rect 214419 457132 214420 457196
rect 214484 457132 214485 457196
rect 214419 457131 214485 457132
rect 216811 457196 216877 457197
rect 216811 457132 216812 457196
rect 216876 457132 216877 457196
rect 216811 457131 216877 457132
rect 210923 456924 210989 456925
rect 210923 456860 210924 456924
rect 210988 456860 210989 456924
rect 210923 456859 210989 456860
rect 212395 456924 212461 456925
rect 212395 456860 212396 456924
rect 212460 456860 212461 456924
rect 212395 456859 212461 456860
rect 213315 456924 213381 456925
rect 213315 456860 213316 456924
rect 213380 456860 213381 456924
rect 213315 456859 213381 456860
rect 216804 443000 217404 457000
rect 217918 456925 217978 459310
rect 218838 458149 218898 460330
rect 219118 459370 219178 460020
rect 220162 459370 220222 460020
rect 219118 459310 219266 459370
rect 218835 458148 218901 458149
rect 218835 458084 218836 458148
rect 218900 458084 218901 458148
rect 218835 458083 218901 458084
rect 219206 456925 219266 459310
rect 220126 459310 220222 459370
rect 220286 459370 220346 460020
rect 221330 459370 221390 460020
rect 220286 459310 220370 459370
rect 221330 459310 221474 459370
rect 220126 458149 220186 459310
rect 220123 458148 220189 458149
rect 220123 458084 220124 458148
rect 220188 458084 220189 458148
rect 220123 458083 220189 458084
rect 220310 457197 220370 459310
rect 221414 458149 221474 459310
rect 221411 458148 221477 458149
rect 221411 458084 221412 458148
rect 221476 458084 221477 458148
rect 221411 458083 221477 458084
rect 220307 457196 220373 457197
rect 220307 457132 220308 457196
rect 220372 457132 220373 457196
rect 220307 457131 220373 457132
rect 217915 456924 217981 456925
rect 217915 456860 217916 456924
rect 217980 456860 217981 456924
rect 217915 456859 217981 456860
rect 219203 456924 219269 456925
rect 219203 456860 219204 456924
rect 219268 456860 219269 456924
rect 219203 456859 219269 456860
rect 220404 443000 221004 457000
rect 221966 456925 222026 460330
rect 222498 459370 222558 460020
rect 222498 459310 222578 459370
rect 222518 458149 222578 459310
rect 222515 458148 222581 458149
rect 222515 458084 222516 458148
rect 222580 458084 222581 458148
rect 222515 458083 222581 458084
rect 223254 456925 223314 460330
rect 224358 460330 224864 460390
rect 224988 460330 225706 460390
rect 223666 459370 223726 460020
rect 223622 459310 223726 459370
rect 223790 459370 223850 460020
rect 223790 459310 223866 459370
rect 223622 458149 223682 459310
rect 223619 458148 223685 458149
rect 223619 458084 223620 458148
rect 223684 458084 223685 458148
rect 223619 458083 223685 458084
rect 223806 456925 223866 459310
rect 224358 458149 224418 460330
rect 224355 458148 224421 458149
rect 224355 458084 224356 458148
rect 224420 458084 224421 458148
rect 224355 458083 224421 458084
rect 225646 457061 225706 460330
rect 225830 460330 226032 460390
rect 228492 460330 229018 460390
rect 231996 460330 232698 460390
rect 225830 458149 225890 460330
rect 226126 459370 226186 460020
rect 227170 459370 227230 460020
rect 226126 459310 226258 459370
rect 225827 458148 225893 458149
rect 225827 458084 225828 458148
rect 225892 458084 225893 458148
rect 225827 458083 225893 458084
rect 225643 457060 225709 457061
rect 221963 456924 222029 456925
rect 221963 456860 221964 456924
rect 222028 456860 222029 456924
rect 221963 456859 222029 456860
rect 223251 456924 223317 456925
rect 223251 456860 223252 456924
rect 223316 456860 223317 456924
rect 223251 456859 223317 456860
rect 223803 456924 223869 456925
rect 223803 456860 223804 456924
rect 223868 456860 223869 456924
rect 223803 456859 223869 456860
rect 224004 443000 224604 457000
rect 225643 456996 225644 457060
rect 225708 456996 225709 457060
rect 225643 456995 225709 456996
rect 226198 456925 226258 459310
rect 227118 459310 227230 459370
rect 227294 459370 227354 460020
rect 228338 459370 228398 460020
rect 227294 459310 227362 459370
rect 228338 459310 228466 459370
rect 227118 458149 227178 459310
rect 227115 458148 227181 458149
rect 227115 458084 227116 458148
rect 227180 458084 227181 458148
rect 227115 458083 227181 458084
rect 227302 456925 227362 459310
rect 228406 458149 228466 459310
rect 228403 458148 228469 458149
rect 228403 458084 228404 458148
rect 228468 458084 228469 458148
rect 228403 458083 228469 458084
rect 226195 456924 226261 456925
rect 226195 456860 226196 456924
rect 226260 456860 226261 456924
rect 226195 456859 226261 456860
rect 227299 456924 227365 456925
rect 227299 456860 227300 456924
rect 227364 456860 227365 456924
rect 227299 456859 227365 456860
rect 227604 445254 228204 457000
rect 228958 456925 229018 460330
rect 229506 459370 229566 460020
rect 229630 459370 229690 460020
rect 230674 459370 230734 460020
rect 229506 459310 229570 459370
rect 229630 459310 229754 459370
rect 229510 458149 229570 459310
rect 229507 458148 229573 458149
rect 229507 458084 229508 458148
rect 229572 458084 229573 458148
rect 229507 458083 229573 458084
rect 229694 456925 229754 459310
rect 230614 459310 230734 459370
rect 230614 457605 230674 459310
rect 230611 457604 230677 457605
rect 230611 457540 230612 457604
rect 230676 457540 230677 457604
rect 230611 457539 230677 457540
rect 230798 456925 230858 460020
rect 231842 459370 231902 460020
rect 231842 459310 231962 459370
rect 231902 457877 231962 459310
rect 231899 457876 231965 457877
rect 231899 457812 231900 457876
rect 231964 457812 231965 457876
rect 231899 457811 231965 457812
rect 232638 457061 232698 460330
rect 232822 460330 233040 460390
rect 233558 460330 234208 460390
rect 234662 460330 235376 460390
rect 235500 460330 235826 460390
rect 232822 458149 232882 460330
rect 233134 459370 233194 460020
rect 233006 459310 233194 459370
rect 232819 458148 232885 458149
rect 232819 458084 232820 458148
rect 232884 458084 232885 458148
rect 232819 458083 232885 458084
rect 232635 457060 232701 457061
rect 232635 456996 232636 457060
rect 232700 456996 232701 457060
rect 232635 456995 232701 456996
rect 233006 456925 233066 459310
rect 233558 458149 233618 460330
rect 234302 459370 234362 460020
rect 234294 459310 234362 459370
rect 233555 458148 233621 458149
rect 233555 458084 233556 458148
rect 233620 458084 233621 458148
rect 233555 458083 233621 458084
rect 234294 456925 234354 459310
rect 234662 458013 234722 460330
rect 234659 458012 234725 458013
rect 234659 457948 234660 458012
rect 234724 457948 234725 458012
rect 234659 457947 234725 457948
rect 228955 456924 229021 456925
rect 228955 456860 228956 456924
rect 229020 456860 229021 456924
rect 228955 456859 229021 456860
rect 229691 456924 229757 456925
rect 229691 456860 229692 456924
rect 229756 456860 229757 456924
rect 229691 456859 229757 456860
rect 230795 456924 230861 456925
rect 230795 456860 230796 456924
rect 230860 456860 230861 456924
rect 230795 456859 230861 456860
rect 233003 456924 233069 456925
rect 233003 456860 233004 456924
rect 233068 456860 233069 456924
rect 233003 456859 233069 456860
rect 234291 456924 234357 456925
rect 234291 456860 234292 456924
rect 234356 456860 234357 456924
rect 234291 456859 234357 456860
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 443000 228204 444698
rect 234804 452454 235404 457000
rect 235766 456925 235826 460330
rect 237422 460330 237712 460390
rect 239004 460330 239690 460390
rect 236514 459370 236574 460020
rect 236502 459310 236574 459370
rect 236638 459370 236698 460020
rect 236638 459310 236746 459370
rect 236502 457877 236562 459310
rect 236499 457876 236565 457877
rect 236499 457812 236500 457876
rect 236564 457812 236565 457876
rect 236499 457811 236565 457812
rect 236686 456925 236746 459310
rect 237422 457741 237482 460330
rect 237806 459370 237866 460020
rect 237790 459310 237866 459370
rect 238850 459370 238910 460020
rect 238850 459310 238954 459370
rect 237419 457740 237485 457741
rect 237419 457676 237420 457740
rect 237484 457676 237485 457740
rect 237419 457675 237485 457676
rect 237790 456925 237850 459310
rect 238894 457741 238954 459310
rect 238891 457740 238957 457741
rect 238891 457676 238892 457740
rect 238956 457676 238957 457740
rect 238891 457675 238957 457676
rect 235763 456924 235829 456925
rect 235763 456860 235764 456924
rect 235828 456860 235829 456924
rect 235763 456859 235829 456860
rect 236683 456924 236749 456925
rect 236683 456860 236684 456924
rect 236748 456860 236749 456924
rect 236683 456859 236749 456860
rect 237787 456924 237853 456925
rect 237787 456860 237788 456924
rect 237852 456860 237853 456924
rect 237787 456859 237853 456860
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 443000 235404 451898
rect 238404 456054 239004 457000
rect 239630 456925 239690 460330
rect 239627 456924 239693 456925
rect 239627 456860 239628 456924
rect 239692 456860 239693 456924
rect 239627 456859 239693 456860
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 443000 239004 455498
rect 242004 443000 242604 457000
rect 245604 443000 246204 457000
rect 252804 443000 253404 457000
rect 256404 443000 257004 457000
rect 260004 443000 260604 457000
rect 263604 445254 264204 457000
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 443000 264204 444698
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 443000 271404 451898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 443000 275004 455498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 443000 278604 459098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 443000 282204 462698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 443000 289404 469898
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 443000 293004 473498
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299427 673844 299493 673845
rect 299427 673780 299428 673844
rect 299492 673780 299493 673844
rect 299427 673779 299493 673780
rect 299430 673573 299490 673779
rect 299427 673572 299493 673573
rect 299427 673508 299428 673572
rect 299492 673508 299493 673572
rect 299427 673507 299493 673508
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299427 650316 299493 650317
rect 299427 650252 299428 650316
rect 299492 650252 299493 650316
rect 299427 650251 299493 650252
rect 299430 650045 299490 650251
rect 299427 650044 299493 650045
rect 299427 649980 299428 650044
rect 299492 649980 299493 650044
rect 299427 649979 299493 649980
rect 299427 626924 299493 626925
rect 299427 626860 299428 626924
rect 299492 626860 299493 626924
rect 299427 626859 299493 626860
rect 299430 626653 299490 626859
rect 299427 626652 299493 626653
rect 299427 626588 299428 626652
rect 299492 626588 299493 626652
rect 299427 626587 299493 626588
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299427 603396 299493 603397
rect 299427 603332 299428 603396
rect 299492 603332 299493 603396
rect 299427 603331 299493 603332
rect 299430 603125 299490 603331
rect 299427 603124 299493 603125
rect 299427 603060 299428 603124
rect 299492 603060 299493 603124
rect 299427 603059 299493 603060
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 443000 296604 477098
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 554247 307404 559898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 554247 311004 563498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 554247 314604 567098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 554247 318204 570698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 554247 325404 577898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 554247 329004 581498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 554247 332604 585098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 554247 336204 588698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 554247 343404 559898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 554247 347004 563498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 554247 350604 567098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 554247 354204 570698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 554247 361404 577898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 554247 365004 581498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 554247 368604 585098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 554247 372204 588698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 554247 379404 559898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 554247 383004 563498
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 554247 386604 567098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 554247 390204 570698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 378547 553484 378613 553485
rect 378547 553420 378548 553484
rect 378612 553420 378613 553484
rect 378547 553419 378613 553420
rect 382963 553484 383029 553485
rect 382963 553420 382964 553484
rect 383028 553420 383029 553484
rect 382963 553419 383029 553420
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 378550 551110 378610 553419
rect 382966 551170 383026 553419
rect 382966 551110 383603 551170
rect 386494 546054 386814 546076
rect 386494 545818 386536 546054
rect 386772 545818 386814 546054
rect 386494 545734 386814 545818
rect 386494 545498 386536 545734
rect 386772 545498 386814 545734
rect 386494 545476 386814 545498
rect 386494 542454 386814 542476
rect 386494 542218 386536 542454
rect 386772 542218 386814 542454
rect 386494 542134 386814 542218
rect 386494 541898 386536 542134
rect 386772 541898 386814 542134
rect 386494 541876 386814 541898
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 386938 535254 387262 535276
rect 386938 535018 386982 535254
rect 387218 535018 387262 535254
rect 386938 534934 387262 535018
rect 386938 534698 386982 534934
rect 387218 534698 387262 534934
rect 386938 534676 387262 534698
rect 386938 531654 387262 531676
rect 386938 531418 386982 531654
rect 387218 531418 387262 531654
rect 386938 531334 387262 531418
rect 386938 531098 386982 531334
rect 387218 531098 387262 531334
rect 386938 531076 387262 531098
rect 386938 528054 387262 528076
rect 386938 527818 386982 528054
rect 387218 527818 387262 528054
rect 386938 527734 387262 527818
rect 386938 527498 386982 527734
rect 387218 527498 387262 527734
rect 386938 527476 387262 527498
rect 386938 524454 387262 524476
rect 386938 524218 386982 524454
rect 387218 524218 387262 524454
rect 386938 524134 387262 524218
rect 386938 523898 386982 524134
rect 387218 523898 387262 524134
rect 386938 523876 387262 523898
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 386494 517254 386814 517276
rect 386494 517018 386536 517254
rect 386772 517018 386814 517254
rect 386494 516934 386814 517018
rect 386494 516698 386536 516934
rect 386772 516698 386814 516934
rect 386494 516676 386814 516698
rect 386494 513654 386814 513676
rect 386494 513418 386536 513654
rect 386772 513418 386814 513654
rect 386494 513334 386814 513418
rect 386494 513098 386536 513334
rect 386772 513098 386814 513334
rect 386494 513076 386814 513098
rect 386494 510054 386814 510076
rect 386494 509818 386536 510054
rect 386772 509818 386814 510054
rect 386494 509734 386814 509818
rect 386494 509498 386536 509734
rect 386772 509498 386814 509734
rect 386494 509476 386814 509498
rect 386494 506454 386814 506476
rect 386494 506218 386536 506454
rect 386772 506218 386814 506454
rect 386494 506134 386814 506218
rect 386494 505898 386536 506134
rect 386772 505898 386814 506134
rect 386494 505876 386814 505898
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 386938 499254 387262 499276
rect 386938 499018 386982 499254
rect 387218 499018 387262 499254
rect 386938 498934 387262 499018
rect 386938 498698 386982 498934
rect 387218 498698 387262 498934
rect 386938 498676 387262 498698
rect 386938 495654 387262 495676
rect 386938 495418 386982 495654
rect 387218 495418 387262 495654
rect 386938 495334 387262 495418
rect 386938 495098 386982 495334
rect 387218 495098 387262 495334
rect 386938 495076 387262 495098
rect 386938 492054 387262 492076
rect 386938 491818 386982 492054
rect 387218 491818 387262 492054
rect 386938 491734 387262 491818
rect 386938 491498 386982 491734
rect 387218 491498 387262 491734
rect 386938 491476 387262 491498
rect 386938 488454 387262 488476
rect 386938 488218 386982 488454
rect 387218 488218 387262 488454
rect 386938 488134 387262 488218
rect 386938 487898 386982 488134
rect 387218 487898 387262 488134
rect 386938 487876 387262 487898
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 386494 481254 386814 481276
rect 386494 481018 386536 481254
rect 386772 481018 386814 481254
rect 386494 480934 386814 481018
rect 386494 480698 386536 480934
rect 386772 480698 386814 480934
rect 386494 480676 386814 480698
rect 386494 477654 386814 477676
rect 386494 477418 386536 477654
rect 386772 477418 386814 477654
rect 386494 477334 386814 477418
rect 386494 477098 386536 477334
rect 386772 477098 386814 477334
rect 386494 477076 386814 477098
rect 386494 474054 386814 474076
rect 386494 473818 386536 474054
rect 386772 473818 386814 474054
rect 386494 473734 386814 473818
rect 386494 473498 386536 473734
rect 386772 473498 386814 473734
rect 386494 473476 386814 473498
rect 386494 470454 386814 470476
rect 386494 470218 386536 470454
rect 386772 470218 386814 470454
rect 386494 470134 386814 470218
rect 386494 469898 386536 470134
rect 386772 469898 386814 470134
rect 386494 469876 386814 469898
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 386938 463254 387262 463276
rect 386938 463018 386982 463254
rect 387218 463018 387262 463254
rect 386938 462934 387262 463018
rect 386938 462698 386982 462934
rect 387218 462698 387262 462934
rect 386938 462676 387262 462698
rect 323534 460670 323840 460730
rect 334022 460670 334352 460730
rect 339910 460670 340192 460730
rect 346902 460670 347200 460730
rect 357390 460670 357712 460730
rect 316174 460330 316832 460390
rect 317462 460330 318000 460390
rect 320958 460330 321504 460390
rect 313803 459370 313863 460020
rect 313782 459310 313863 459370
rect 313782 458149 313842 459310
rect 313779 458148 313845 458149
rect 313779 458084 313780 458148
rect 313844 458084 313845 458148
rect 313779 458083 313845 458084
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 443000 300204 444698
rect 306804 452454 307404 457000
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 59126 438910 59370 438970
rect 59126 297941 59186 438910
rect 64208 434454 64528 434476
rect 64208 434218 64250 434454
rect 64486 434218 64528 434454
rect 64208 434134 64528 434218
rect 64208 433898 64250 434134
rect 64486 433898 64528 434134
rect 64208 433876 64528 433898
rect 79568 427254 79888 427276
rect 79568 427018 79610 427254
rect 79846 427018 79888 427254
rect 79568 426934 79888 427018
rect 79568 426698 79610 426934
rect 79846 426698 79888 426934
rect 79568 426676 79888 426698
rect 79568 423654 79888 423676
rect 79568 423418 79610 423654
rect 79846 423418 79888 423654
rect 79568 423334 79888 423418
rect 79568 423098 79610 423334
rect 79846 423098 79888 423334
rect 79568 423076 79888 423098
rect 79568 420054 79888 420076
rect 79568 419818 79610 420054
rect 79846 419818 79888 420054
rect 79568 419734 79888 419818
rect 79568 419498 79610 419734
rect 79846 419498 79888 419734
rect 79568 419476 79888 419498
rect 79568 416454 79888 416476
rect 79568 416218 79610 416454
rect 79846 416218 79888 416454
rect 79568 416134 79888 416218
rect 79568 415898 79610 416134
rect 79846 415898 79888 416134
rect 79568 415876 79888 415898
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 64208 409254 64528 409276
rect 64208 409018 64250 409254
rect 64486 409018 64528 409254
rect 64208 408934 64528 409018
rect 64208 408698 64250 408934
rect 64486 408698 64528 408934
rect 64208 408676 64528 408698
rect 64208 405654 64528 405676
rect 64208 405418 64250 405654
rect 64486 405418 64528 405654
rect 64208 405334 64528 405418
rect 64208 405098 64250 405334
rect 64486 405098 64528 405334
rect 64208 405076 64528 405098
rect 64208 402054 64528 402076
rect 64208 401818 64250 402054
rect 64486 401818 64528 402054
rect 64208 401734 64528 401818
rect 64208 401498 64250 401734
rect 64486 401498 64528 401734
rect 64208 401476 64528 401498
rect 64208 398454 64528 398476
rect 64208 398218 64250 398454
rect 64486 398218 64528 398454
rect 64208 398134 64528 398218
rect 64208 397898 64250 398134
rect 64486 397898 64528 398134
rect 64208 397876 64528 397898
rect 79568 391254 79888 391276
rect 79568 391018 79610 391254
rect 79846 391018 79888 391254
rect 79568 390934 79888 391018
rect 79568 390698 79610 390934
rect 79846 390698 79888 390934
rect 79568 390676 79888 390698
rect 79568 387654 79888 387676
rect 79568 387418 79610 387654
rect 79846 387418 79888 387654
rect 79568 387334 79888 387418
rect 79568 387098 79610 387334
rect 79846 387098 79888 387334
rect 79568 387076 79888 387098
rect 79568 384054 79888 384076
rect 79568 383818 79610 384054
rect 79846 383818 79888 384054
rect 79568 383734 79888 383818
rect 79568 383498 79610 383734
rect 79846 383498 79888 383734
rect 79568 383476 79888 383498
rect 79568 380454 79888 380476
rect 79568 380218 79610 380454
rect 79846 380218 79888 380454
rect 79568 380134 79888 380218
rect 79568 379898 79610 380134
rect 79846 379898 79888 380134
rect 79568 379876 79888 379898
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 64208 373254 64528 373276
rect 64208 373018 64250 373254
rect 64486 373018 64528 373254
rect 64208 372934 64528 373018
rect 64208 372698 64250 372934
rect 64486 372698 64528 372934
rect 64208 372676 64528 372698
rect 64208 369654 64528 369676
rect 64208 369418 64250 369654
rect 64486 369418 64528 369654
rect 64208 369334 64528 369418
rect 64208 369098 64250 369334
rect 64486 369098 64528 369334
rect 64208 369076 64528 369098
rect 64208 366054 64528 366076
rect 64208 365818 64250 366054
rect 64486 365818 64528 366054
rect 64208 365734 64528 365818
rect 64208 365498 64250 365734
rect 64486 365498 64528 365734
rect 64208 365476 64528 365498
rect 64208 362454 64528 362476
rect 64208 362218 64250 362454
rect 64486 362218 64528 362454
rect 64208 362134 64528 362218
rect 64208 361898 64250 362134
rect 64486 361898 64528 362134
rect 64208 361876 64528 361898
rect 79568 355254 79888 355276
rect 79568 355018 79610 355254
rect 79846 355018 79888 355254
rect 79568 354934 79888 355018
rect 79568 354698 79610 354934
rect 79846 354698 79888 354934
rect 79568 354676 79888 354698
rect 79568 351654 79888 351676
rect 79568 351418 79610 351654
rect 79846 351418 79888 351654
rect 79568 351334 79888 351418
rect 79568 351098 79610 351334
rect 79846 351098 79888 351334
rect 79568 351076 79888 351098
rect 79568 348054 79888 348076
rect 79568 347818 79610 348054
rect 79846 347818 79888 348054
rect 79568 347734 79888 347818
rect 79568 347498 79610 347734
rect 79846 347498 79888 347734
rect 79568 347476 79888 347498
rect 79568 344454 79888 344476
rect 79568 344218 79610 344454
rect 79846 344218 79888 344454
rect 79568 344134 79888 344218
rect 79568 343898 79610 344134
rect 79846 343898 79888 344134
rect 79568 343876 79888 343898
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 64208 337254 64528 337276
rect 64208 337018 64250 337254
rect 64486 337018 64528 337254
rect 64208 336934 64528 337018
rect 64208 336698 64250 336934
rect 64486 336698 64528 336934
rect 64208 336676 64528 336698
rect 64208 333654 64528 333676
rect 64208 333418 64250 333654
rect 64486 333418 64528 333654
rect 64208 333334 64528 333418
rect 64208 333098 64250 333334
rect 64486 333098 64528 333334
rect 64208 333076 64528 333098
rect 64208 330054 64528 330076
rect 64208 329818 64250 330054
rect 64486 329818 64528 330054
rect 64208 329734 64528 329818
rect 64208 329498 64250 329734
rect 64486 329498 64528 329734
rect 64208 329476 64528 329498
rect 64208 326454 64528 326476
rect 64208 326218 64250 326454
rect 64486 326218 64528 326454
rect 64208 326134 64528 326218
rect 64208 325898 64250 326134
rect 64486 325898 64528 326134
rect 64208 325876 64528 325898
rect 79568 319254 79888 319276
rect 79568 319018 79610 319254
rect 79846 319018 79888 319254
rect 79568 318934 79888 319018
rect 79568 318698 79610 318934
rect 79846 318698 79888 318934
rect 79568 318676 79888 318698
rect 79568 315654 79888 315676
rect 79568 315418 79610 315654
rect 79846 315418 79888 315654
rect 79568 315334 79888 315418
rect 79568 315098 79610 315334
rect 79846 315098 79888 315334
rect 79568 315076 79888 315098
rect 79568 312054 79888 312076
rect 79568 311818 79610 312054
rect 79846 311818 79888 312054
rect 79568 311734 79888 311818
rect 79568 311498 79610 311734
rect 79846 311498 79888 311734
rect 79568 311476 79888 311498
rect 79568 308454 79888 308476
rect 79568 308218 79610 308454
rect 79846 308218 79888 308454
rect 79568 308134 79888 308218
rect 79568 307898 79610 308134
rect 79846 307898 79888 308134
rect 79568 307876 79888 307898
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 64208 301254 64528 301276
rect 64208 301018 64250 301254
rect 64486 301018 64528 301254
rect 64208 300934 64528 301018
rect 64208 300698 64250 300934
rect 64486 300698 64528 300934
rect 64208 300676 64528 300698
rect 59123 297940 59189 297941
rect 59123 297876 59124 297940
rect 59188 297876 59189 297940
rect 59123 297875 59189 297876
rect 64208 297654 64528 297676
rect 64208 297418 64250 297654
rect 64486 297418 64528 297654
rect 64208 297334 64528 297418
rect 64208 297098 64250 297334
rect 64486 297098 64528 297334
rect 64208 297076 64528 297098
rect 64208 294054 64528 294076
rect 64208 293818 64250 294054
rect 64486 293818 64528 294054
rect 64208 293734 64528 293818
rect 64208 293498 64250 293734
rect 64486 293498 64528 293734
rect 64208 293476 64528 293498
rect 64208 290454 64528 290476
rect 64208 290218 64250 290454
rect 64486 290218 64528 290454
rect 64208 290134 64528 290218
rect 64208 289898 64250 290134
rect 64486 289898 64528 290134
rect 64208 289876 64528 289898
rect 79568 283254 79888 283276
rect 79568 283018 79610 283254
rect 79846 283018 79888 283254
rect 79568 282934 79888 283018
rect 79568 282698 79610 282934
rect 79846 282698 79888 282934
rect 79568 282676 79888 282698
rect 79568 279654 79888 279676
rect 79568 279418 79610 279654
rect 79846 279418 79888 279654
rect 79568 279334 79888 279418
rect 79568 279098 79610 279334
rect 79846 279098 79888 279334
rect 79568 279076 79888 279098
rect 58939 278900 59005 278901
rect 58939 278836 58940 278900
rect 59004 278836 59005 278900
rect 58939 278835 59005 278836
rect 79568 276054 79888 276076
rect 79568 275818 79610 276054
rect 79846 275818 79888 276054
rect 79568 275734 79888 275818
rect 79568 275498 79610 275734
rect 79846 275498 79888 275734
rect 79568 275476 79888 275498
rect 79568 272454 79888 272476
rect 79568 272218 79610 272454
rect 79846 272218 79888 272454
rect 79568 272134 79888 272218
rect 79568 271898 79610 272134
rect 79846 271898 79888 272134
rect 79568 271876 79888 271898
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 57099 266252 57165 266253
rect 57099 266188 57100 266252
rect 57164 266188 57165 266252
rect 57099 266187 57165 266188
rect 64208 265254 64528 265276
rect 64208 265018 64250 265254
rect 64486 265018 64528 265254
rect 64208 264934 64528 265018
rect 64208 264698 64250 264934
rect 64486 264698 64528 264934
rect 64208 264676 64528 264698
rect 64208 261654 64528 261676
rect 64208 261418 64250 261654
rect 64486 261418 64528 261654
rect 64208 261334 64528 261418
rect 64208 261098 64250 261334
rect 64486 261098 64528 261334
rect 64208 261076 64528 261098
rect 64208 258054 64528 258076
rect 64208 257818 64250 258054
rect 64486 257818 64528 258054
rect 64208 257734 64528 257818
rect 64208 257498 64250 257734
rect 64486 257498 64528 257734
rect 64208 257476 64528 257498
rect 64208 254454 64528 254476
rect 64208 254218 64250 254454
rect 64486 254218 64528 254454
rect 64208 254134 64528 254218
rect 64208 253898 64250 254134
rect 64486 253898 64528 254134
rect 64208 253876 64528 253898
rect 57651 249524 57717 249525
rect 57651 249460 57652 249524
rect 57716 249460 57717 249524
rect 57651 249459 57717 249460
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 56915 213620 56981 213621
rect 56915 213556 56916 213620
rect 56980 213556 56981 213620
rect 56915 213555 56981 213556
rect 56731 205188 56797 205189
rect 56731 205124 56732 205188
rect 56796 205124 56797 205188
rect 56731 205123 56797 205124
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 56734 29341 56794 205123
rect 56918 110805 56978 213555
rect 57283 211580 57349 211581
rect 57283 211516 57284 211580
rect 57348 211516 57349 211580
rect 57283 211515 57349 211516
rect 57099 209404 57165 209405
rect 57099 209340 57100 209404
rect 57164 209340 57165 209404
rect 57099 209339 57165 209340
rect 56915 110804 56981 110805
rect 56915 110740 56916 110804
rect 56980 110740 56981 110804
rect 56915 110739 56981 110740
rect 57102 87277 57162 209339
rect 57099 87276 57165 87277
rect 57099 87212 57100 87276
rect 57164 87212 57165 87276
rect 57099 87211 57165 87212
rect 57286 76261 57346 211515
rect 57467 207364 57533 207365
rect 57467 207300 57468 207364
rect 57532 207300 57533 207364
rect 57467 207299 57533 207300
rect 57283 76260 57349 76261
rect 57283 76196 57284 76260
rect 57348 76196 57349 76260
rect 57283 76195 57349 76196
rect 57470 63885 57530 207299
rect 57654 205053 57714 249459
rect 57835 247348 57901 247349
rect 57835 247284 57836 247348
rect 57900 247284 57901 247348
rect 57835 247283 57901 247284
rect 57651 205052 57717 205053
rect 57651 204988 57652 205052
rect 57716 204988 57717 205052
rect 57651 204987 57717 204988
rect 57651 203148 57717 203149
rect 57651 203084 57652 203148
rect 57716 203084 57717 203148
rect 57651 203083 57717 203084
rect 57467 63884 57533 63885
rect 57467 63820 57468 63884
rect 57532 63820 57533 63884
rect 57467 63819 57533 63820
rect 57654 40357 57714 203083
rect 57838 200701 57898 247283
rect 79568 247254 79888 247276
rect 79568 247018 79610 247254
rect 79846 247018 79888 247254
rect 79568 246934 79888 247018
rect 79568 246698 79610 246934
rect 79846 246698 79888 246934
rect 79568 246676 79888 246698
rect 79568 243654 79888 243676
rect 79568 243418 79610 243654
rect 79846 243418 79888 243654
rect 79568 243334 79888 243418
rect 79568 243098 79610 243334
rect 79846 243098 79888 243334
rect 79568 243076 79888 243098
rect 79568 240054 79888 240076
rect 79568 239818 79610 240054
rect 79846 239818 79888 240054
rect 79568 239734 79888 239818
rect 79568 239498 79610 239734
rect 79846 239498 79888 239734
rect 79568 239476 79888 239498
rect 79568 236454 79888 236476
rect 79568 236218 79610 236454
rect 79846 236218 79888 236454
rect 79568 236134 79888 236218
rect 79568 235898 79610 236134
rect 79846 235898 79888 236134
rect 79568 235876 79888 235898
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 64208 229254 64528 229276
rect 64208 229018 64250 229254
rect 64486 229018 64528 229254
rect 64208 228934 64528 229018
rect 64208 228698 64250 228934
rect 64486 228698 64528 228934
rect 64208 228676 64528 228698
rect 64208 225654 64528 225676
rect 64208 225418 64250 225654
rect 64486 225418 64528 225654
rect 64208 225334 64528 225418
rect 64208 225098 64250 225334
rect 64486 225098 64528 225334
rect 64208 225076 64528 225098
rect 64208 222054 64528 222076
rect 64208 221818 64250 222054
rect 64486 221818 64528 222054
rect 64208 221734 64528 221818
rect 64208 221498 64250 221734
rect 64486 221498 64528 221734
rect 64208 221476 64528 221498
rect 64208 218454 64528 218476
rect 64208 218218 64250 218454
rect 64486 218218 64528 218454
rect 64208 218134 64528 218218
rect 64208 217898 64250 218134
rect 64486 217898 64528 218134
rect 64208 217876 64528 217898
rect 79568 211254 79888 211276
rect 79568 211018 79610 211254
rect 79846 211018 79888 211254
rect 79568 210934 79888 211018
rect 79568 210698 79610 210934
rect 79846 210698 79888 210934
rect 79568 210676 79888 210698
rect 79568 207654 79888 207676
rect 79568 207418 79610 207654
rect 79846 207418 79888 207654
rect 79568 207334 79888 207418
rect 79568 207098 79610 207334
rect 79846 207098 79888 207334
rect 79568 207076 79888 207098
rect 79568 204054 79888 204076
rect 79568 203818 79610 204054
rect 79846 203818 79888 204054
rect 79568 203734 79888 203818
rect 79568 203498 79610 203734
rect 79846 203498 79888 203734
rect 79568 203476 79888 203498
rect 57835 200700 57901 200701
rect 57835 200636 57836 200700
rect 57900 200636 57901 200700
rect 57835 200635 57901 200636
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 58404 168054 59004 197000
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 57651 40356 57717 40357
rect 57651 40292 57652 40356
rect 57716 40292 57717 40356
rect 57651 40291 57717 40292
rect 56731 29340 56797 29341
rect 56731 29276 56732 29340
rect 56796 29276 56797 29340
rect 56731 29275 56797 29276
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 171654 62604 197000
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 175254 66204 197000
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 182454 73404 197000
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 186054 77004 197000
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 189654 80604 197000
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 193254 84204 197000
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 164454 91404 197000
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 168054 95004 197000
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 171654 98604 197000
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 175254 102204 197000
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 182454 109404 197000
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 186054 113004 197000
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 116004 189654 116604 197000
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 115795 110940 115861 110941
rect 115795 110876 115796 110940
rect 115860 110876 115861 110940
rect 115795 110875 115861 110876
rect 115798 110533 115858 110875
rect 115795 110532 115861 110533
rect 115795 110468 115796 110532
rect 115860 110468 115861 110532
rect 115795 110467 115861 110468
rect 115795 87412 115861 87413
rect 115795 87348 115796 87412
rect 115860 87348 115861 87412
rect 115795 87347 115861 87348
rect 115798 87005 115858 87347
rect 115795 87004 115861 87005
rect 115795 86940 115796 87004
rect 115860 86940 115861 87004
rect 115795 86939 115861 86940
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 115795 76396 115861 76397
rect 115795 76332 115796 76396
rect 115860 76332 115861 76396
rect 115795 76331 115861 76332
rect 115798 75989 115858 76331
rect 115795 75988 115861 75989
rect 115795 75924 115796 75988
rect 115860 75924 115861 75988
rect 115795 75923 115861 75924
rect 115795 64020 115861 64021
rect 115795 63956 115796 64020
rect 115860 63956 115861 64020
rect 115795 63955 115861 63956
rect 115798 63613 115858 63955
rect 115795 63612 115861 63613
rect 115795 63548 115796 63612
rect 115860 63548 115861 63612
rect 115795 63547 115861 63548
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 115795 40492 115861 40493
rect 115795 40428 115796 40492
rect 115860 40428 115861 40492
rect 115795 40427 115861 40428
rect 115798 40085 115858 40427
rect 115795 40084 115861 40085
rect 115795 40020 115796 40084
rect 115860 40020 115861 40084
rect 115795 40019 115861 40020
rect 115795 29476 115861 29477
rect 115795 29412 115796 29476
rect 115860 29412 115861 29476
rect 115795 29411 115861 29412
rect 115798 29069 115858 29411
rect 115795 29068 115861 29069
rect 115795 29004 115796 29068
rect 115860 29004 115861 29068
rect 115795 29003 115861 29004
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 193254 120204 197000
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 126804 164454 127404 197000
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 125547 111076 125613 111077
rect 125547 111012 125548 111076
rect 125612 111012 125613 111076
rect 125547 111011 125613 111012
rect 125550 110805 125610 111011
rect 125547 110804 125613 110805
rect 125547 110740 125548 110804
rect 125612 110740 125613 110804
rect 125547 110739 125613 110740
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 125547 76532 125613 76533
rect 125547 76468 125548 76532
rect 125612 76468 125613 76532
rect 125547 76467 125613 76468
rect 125550 76261 125610 76467
rect 125547 76260 125613 76261
rect 125547 76196 125548 76260
rect 125612 76196 125613 76260
rect 125547 76195 125613 76196
rect 125547 64156 125613 64157
rect 125547 64092 125548 64156
rect 125612 64092 125613 64156
rect 125547 64091 125613 64092
rect 125550 63885 125610 64091
rect 125547 63884 125613 63885
rect 125547 63820 125548 63884
rect 125612 63820 125613 63884
rect 125547 63819 125613 63820
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 125547 40628 125613 40629
rect 125547 40564 125548 40628
rect 125612 40564 125613 40628
rect 125547 40563 125613 40564
rect 125550 40357 125610 40563
rect 125547 40356 125613 40357
rect 125547 40292 125548 40356
rect 125612 40292 125613 40356
rect 125547 40291 125613 40292
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 168054 131004 197000
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 134004 171654 134604 197000
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 133827 87412 133893 87413
rect 133827 87348 133828 87412
rect 133892 87348 133893 87412
rect 133827 87347 133893 87348
rect 133830 87141 133890 87347
rect 133827 87140 133893 87141
rect 133827 87076 133828 87140
rect 133892 87076 133893 87140
rect 133827 87075 133893 87076
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 133827 29476 133893 29477
rect 133827 29412 133828 29476
rect 133892 29412 133893 29476
rect 133827 29411 133893 29412
rect 133830 29205 133890 29411
rect 133827 29204 133893 29205
rect 133827 29140 133828 29204
rect 133892 29140 133893 29204
rect 133827 29139 133893 29140
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 175254 138204 197000
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 182454 145404 197000
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 186054 149004 197000
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 189654 152604 197000
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 193254 156204 197000
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 164454 163404 197000
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 168054 167004 197000
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 171654 170604 197000
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 175254 174204 197000
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 182454 181404 197000
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 186054 185004 197000
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 189654 188604 197000
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 193254 192204 197000
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 164454 199404 197000
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 168054 203004 197000
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 171654 206604 197000
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 175254 210204 197000
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 182454 217404 197000
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 186054 221004 197000
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 189654 224604 197000
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 193254 228204 197000
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 164454 235404 197000
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 168054 239004 197000
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 171654 242604 197000
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 175254 246204 197000
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 182454 253404 197000
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 186054 257004 197000
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 189654 260604 197000
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 193254 264204 197000
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 164454 271404 197000
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 168054 275004 197000
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 171654 278604 197000
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 175254 282204 197000
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 182454 289404 197000
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 186054 293004 197000
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 189654 296604 197000
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 193254 300204 197000
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 456054 311004 457000
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 423654 314604 457000
rect 316174 456925 316234 460330
rect 317462 457877 317522 460330
rect 319138 459370 319198 460020
rect 320306 459370 320366 460020
rect 319118 459310 319198 459370
rect 320222 459310 320366 459370
rect 317459 457876 317525 457877
rect 317459 457812 317460 457876
rect 317524 457812 317525 457876
rect 317459 457811 317525 457812
rect 316171 456924 316237 456925
rect 316171 456860 316172 456924
rect 316236 456860 316237 456924
rect 316171 456859 316237 456860
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 427254 318204 457000
rect 319118 456925 319178 459310
rect 320222 456925 320282 459310
rect 320958 457061 321018 460330
rect 322642 459370 322702 460020
rect 322614 459310 322702 459370
rect 322766 459370 322826 460020
rect 322766 459310 322858 459370
rect 322614 458013 322674 459310
rect 322798 458149 322858 459310
rect 322795 458148 322861 458149
rect 322795 458084 322796 458148
rect 322860 458084 322861 458148
rect 322795 458083 322861 458084
rect 323534 458013 323594 460670
rect 324822 460330 325008 460390
rect 323934 459370 323994 460020
rect 323902 459310 323994 459370
rect 323902 458149 323962 459310
rect 323899 458148 323965 458149
rect 323899 458084 323900 458148
rect 323964 458084 323965 458148
rect 323899 458083 323965 458084
rect 322611 458012 322677 458013
rect 322611 457948 322612 458012
rect 322676 457948 322677 458012
rect 322611 457947 322677 457948
rect 323531 458012 323597 458013
rect 323531 457948 323532 458012
rect 323596 457948 323597 458012
rect 323531 457947 323597 457948
rect 324822 457877 324882 460330
rect 325102 459370 325162 460020
rect 326146 459370 326206 460020
rect 325006 459310 325162 459370
rect 326110 459310 326206 459370
rect 326270 459370 326330 460020
rect 327314 459509 327374 460020
rect 327311 459508 327377 459509
rect 327311 459444 327312 459508
rect 327376 459444 327377 459508
rect 327311 459443 327377 459444
rect 327438 459370 327498 460020
rect 328482 459509 328542 460020
rect 328479 459508 328545 459509
rect 328479 459444 328480 459508
rect 328544 459444 328545 459508
rect 328479 459443 328545 459444
rect 328606 459370 328666 460020
rect 328867 459508 328933 459509
rect 328867 459444 328868 459508
rect 328932 459444 328933 459508
rect 328867 459443 328933 459444
rect 326270 459310 326354 459370
rect 324819 457876 324885 457877
rect 324819 457812 324820 457876
rect 324884 457812 324885 457876
rect 324819 457811 324885 457812
rect 325006 457197 325066 459310
rect 326110 457877 326170 459310
rect 326294 458149 326354 459310
rect 327398 459310 327498 459370
rect 328502 459310 328666 459370
rect 327398 458149 327458 459310
rect 326291 458148 326357 458149
rect 326291 458084 326292 458148
rect 326356 458084 326357 458148
rect 326291 458083 326357 458084
rect 327395 458148 327461 458149
rect 327395 458084 327396 458148
rect 327460 458084 327461 458148
rect 327395 458083 327461 458084
rect 326107 457876 326173 457877
rect 326107 457812 326108 457876
rect 326172 457812 326173 457876
rect 326107 457811 326173 457812
rect 328502 457197 328562 459310
rect 328870 458149 328930 459443
rect 329650 459370 329710 460020
rect 329606 459310 329710 459370
rect 328867 458148 328933 458149
rect 328867 458084 328868 458148
rect 328932 458084 328933 458148
rect 328867 458083 328933 458084
rect 329606 458013 329666 459310
rect 329603 458012 329669 458013
rect 329603 457948 329604 458012
rect 329668 457948 329669 458012
rect 329603 457947 329669 457948
rect 329790 457333 329850 460390
rect 330526 460330 330848 460390
rect 331814 460330 332016 460390
rect 330526 457877 330586 460330
rect 330942 459370 331002 460020
rect 330894 459310 331002 459370
rect 330894 458149 330954 459310
rect 331814 458149 331874 460330
rect 332110 459370 332170 460020
rect 333154 459370 333214 460020
rect 331998 459310 332170 459370
rect 333102 459310 333214 459370
rect 333278 459370 333338 460020
rect 333278 459310 333346 459370
rect 330891 458148 330957 458149
rect 330891 458084 330892 458148
rect 330956 458084 330957 458148
rect 330891 458083 330957 458084
rect 331811 458148 331877 458149
rect 331811 458084 331812 458148
rect 331876 458084 331877 458148
rect 331811 458083 331877 458084
rect 330523 457876 330589 457877
rect 330523 457812 330524 457876
rect 330588 457812 330589 457876
rect 330523 457811 330589 457812
rect 331998 457741 332058 459310
rect 333102 458149 333162 459310
rect 333099 458148 333165 458149
rect 333099 458084 333100 458148
rect 333164 458084 333165 458148
rect 333099 458083 333165 458084
rect 331995 457740 332061 457741
rect 331995 457676 331996 457740
rect 332060 457676 332061 457740
rect 331995 457675 332061 457676
rect 329787 457332 329853 457333
rect 329787 457268 329788 457332
rect 329852 457268 329853 457332
rect 329787 457267 329853 457268
rect 325003 457196 325069 457197
rect 325003 457132 325004 457196
rect 325068 457132 325069 457196
rect 325003 457131 325069 457132
rect 328499 457196 328565 457197
rect 328499 457132 328500 457196
rect 328564 457132 328565 457196
rect 328499 457131 328565 457132
rect 320955 457060 321021 457061
rect 320955 456996 320956 457060
rect 321020 456996 321021 457060
rect 320955 456995 321021 456996
rect 319115 456924 319181 456925
rect 319115 456860 319116 456924
rect 319180 456860 319181 456924
rect 319115 456859 319181 456860
rect 320219 456924 320285 456925
rect 320219 456860 320220 456924
rect 320284 456860 320285 456924
rect 320219 456859 320285 456860
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 434454 325404 457000
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 438054 329004 457000
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 441654 332604 457000
rect 333286 456925 333346 459310
rect 334022 458149 334082 460670
rect 335310 460330 335520 460390
rect 337702 460330 337856 460390
rect 334446 459370 334506 460020
rect 334390 459310 334506 459370
rect 334019 458148 334085 458149
rect 334019 458084 334020 458148
rect 334084 458084 334085 458148
rect 334019 458083 334085 458084
rect 334390 456925 334450 459310
rect 335310 458149 335370 460330
rect 335614 459370 335674 460020
rect 336658 459370 336718 460020
rect 335494 459310 335674 459370
rect 336598 459310 336718 459370
rect 335307 458148 335373 458149
rect 335307 458084 335308 458148
rect 335372 458084 335373 458148
rect 335307 458083 335373 458084
rect 335494 457197 335554 459310
rect 336598 458149 336658 459310
rect 336595 458148 336661 458149
rect 336595 458084 336596 458148
rect 336660 458084 336661 458148
rect 336595 458083 336661 458084
rect 335491 457196 335557 457197
rect 335491 457132 335492 457196
rect 335556 457132 335557 457196
rect 335491 457131 335557 457132
rect 333283 456924 333349 456925
rect 333283 456860 333284 456924
rect 333348 456860 333349 456924
rect 333283 456859 333349 456860
rect 334387 456924 334453 456925
rect 334387 456860 334388 456924
rect 334452 456860 334453 456924
rect 334387 456859 334453 456860
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 445254 336204 457000
rect 336782 456925 336842 460020
rect 337702 458149 337762 460330
rect 337950 459370 338010 460020
rect 338994 459370 339054 460020
rect 337886 459310 338010 459370
rect 338990 459310 339054 459370
rect 339118 459370 339178 460020
rect 339118 459310 339234 459370
rect 337699 458148 337765 458149
rect 337699 458084 337700 458148
rect 337764 458084 337765 458148
rect 337699 458083 337765 458084
rect 337886 457061 337946 459310
rect 338990 458149 339050 459310
rect 338987 458148 339053 458149
rect 338987 458084 338988 458148
rect 339052 458084 339053 458148
rect 338987 458083 339053 458084
rect 337883 457060 337949 457061
rect 337883 456996 337884 457060
rect 337948 456996 337949 457060
rect 337883 456995 337949 456996
rect 339174 456925 339234 459310
rect 339910 458149 339970 460670
rect 341198 460330 341360 460390
rect 343820 460330 344018 460390
rect 340286 459370 340346 460020
rect 340278 459310 340346 459370
rect 339907 458148 339973 458149
rect 339907 458084 339908 458148
rect 339972 458084 339973 458148
rect 339907 458083 339973 458084
rect 340278 456925 340338 459310
rect 341198 458149 341258 460330
rect 341454 459370 341514 460020
rect 342498 459370 342558 460020
rect 341382 459310 341514 459370
rect 342486 459310 342558 459370
rect 342622 459370 342682 460020
rect 343666 459370 343726 460020
rect 342622 459310 342730 459370
rect 341195 458148 341261 458149
rect 341195 458084 341196 458148
rect 341260 458084 341261 458148
rect 341195 458083 341261 458084
rect 341382 457197 341442 459310
rect 342486 458013 342546 459310
rect 342670 458149 342730 459310
rect 343590 459310 343726 459370
rect 342667 458148 342733 458149
rect 342667 458084 342668 458148
rect 342732 458084 342733 458148
rect 342667 458083 342733 458084
rect 343590 458013 343650 459310
rect 343958 458149 344018 460330
rect 344694 460330 344864 460390
rect 344694 458149 344754 460330
rect 344958 459370 345018 460020
rect 346002 459370 346062 460020
rect 344878 459310 345018 459370
rect 345982 459310 346062 459370
rect 346126 459370 346186 460020
rect 346126 459310 346226 459370
rect 343955 458148 344021 458149
rect 343955 458084 343956 458148
rect 344020 458084 344021 458148
rect 343955 458083 344021 458084
rect 344691 458148 344757 458149
rect 344691 458084 344692 458148
rect 344756 458084 344757 458148
rect 344691 458083 344757 458084
rect 342483 458012 342549 458013
rect 342483 457948 342484 458012
rect 342548 457948 342549 458012
rect 342483 457947 342549 457948
rect 343587 458012 343653 458013
rect 343587 457948 343588 458012
rect 343652 457948 343653 458012
rect 343587 457947 343653 457948
rect 344878 457741 344938 459310
rect 345982 458013 346042 459310
rect 346166 458149 346226 459310
rect 346163 458148 346229 458149
rect 346163 458084 346164 458148
rect 346228 458084 346229 458148
rect 346163 458083 346229 458084
rect 346902 458013 346962 460670
rect 348190 460330 348368 460390
rect 350828 460330 351010 460390
rect 347294 459370 347354 460020
rect 347270 459310 347354 459370
rect 347270 458149 347330 459310
rect 347267 458148 347333 458149
rect 347267 458084 347268 458148
rect 347332 458084 347333 458148
rect 347267 458083 347333 458084
rect 348190 458013 348250 460330
rect 348462 459370 348522 460020
rect 349506 459370 349566 460020
rect 348374 459310 348522 459370
rect 349478 459310 349566 459370
rect 349630 459370 349690 460020
rect 350674 459370 350734 460020
rect 349630 459310 349722 459370
rect 348374 458149 348434 459310
rect 348371 458148 348437 458149
rect 348371 458084 348372 458148
rect 348436 458084 348437 458148
rect 348371 458083 348437 458084
rect 349478 458013 349538 459310
rect 349662 458149 349722 459310
rect 350582 459310 350734 459370
rect 349659 458148 349725 458149
rect 349659 458084 349660 458148
rect 349724 458084 349725 458148
rect 349659 458083 349725 458084
rect 350582 458013 350642 459310
rect 345979 458012 346045 458013
rect 345979 457948 345980 458012
rect 346044 457948 346045 458012
rect 345979 457947 346045 457948
rect 346899 458012 346965 458013
rect 346899 457948 346900 458012
rect 346964 457948 346965 458012
rect 346899 457947 346965 457948
rect 348187 458012 348253 458013
rect 348187 457948 348188 458012
rect 348252 457948 348253 458012
rect 348187 457947 348253 457948
rect 349475 458012 349541 458013
rect 349475 457948 349476 458012
rect 349540 457948 349541 458012
rect 349475 457947 349541 457948
rect 350579 458012 350645 458013
rect 350579 457948 350580 458012
rect 350644 457948 350645 458012
rect 350579 457947 350645 457948
rect 344875 457740 344941 457741
rect 344875 457676 344876 457740
rect 344940 457676 344941 457740
rect 344875 457675 344941 457676
rect 341379 457196 341445 457197
rect 341379 457132 341380 457196
rect 341444 457132 341445 457196
rect 341379 457131 341445 457132
rect 336779 456924 336845 456925
rect 336779 456860 336780 456924
rect 336844 456860 336845 456924
rect 336779 456859 336845 456860
rect 339171 456924 339237 456925
rect 339171 456860 339172 456924
rect 339236 456860 339237 456924
rect 339171 456859 339237 456860
rect 340275 456924 340341 456925
rect 340275 456860 340276 456924
rect 340340 456860 340341 456924
rect 340275 456859 340341 456860
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 452454 343404 457000
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 456054 347004 457000
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 423654 350604 457000
rect 350950 456925 351010 460330
rect 353526 460330 354208 460390
rect 355182 460330 355376 460390
rect 351842 459645 351902 460020
rect 351839 459644 351905 459645
rect 351839 459580 351840 459644
rect 351904 459580 351905 459644
rect 351839 459579 351905 459580
rect 351966 459370 352026 460020
rect 353010 459370 353070 460020
rect 351870 459310 352026 459370
rect 352974 459310 353070 459370
rect 353134 459370 353194 460020
rect 353134 459310 353218 459370
rect 351870 456925 351930 459310
rect 352974 458149 353034 459310
rect 352971 458148 353037 458149
rect 352971 458084 352972 458148
rect 353036 458084 353037 458148
rect 352971 458083 353037 458084
rect 353158 457061 353218 459310
rect 353526 458149 353586 460330
rect 354302 459370 354362 460020
rect 354262 459310 354362 459370
rect 353523 458148 353589 458149
rect 353523 458084 353524 458148
rect 353588 458084 353589 458148
rect 353523 458083 353589 458084
rect 354262 457197 354322 459310
rect 355182 457877 355242 460330
rect 355470 459370 355530 460020
rect 356514 459370 356574 460020
rect 355366 459310 355530 459370
rect 356470 459310 356574 459370
rect 356638 459370 356698 460020
rect 356638 459310 356714 459370
rect 355179 457876 355245 457877
rect 355179 457812 355180 457876
rect 355244 457812 355245 457876
rect 355179 457811 355245 457812
rect 354259 457196 354325 457197
rect 354259 457132 354260 457196
rect 354324 457132 354325 457196
rect 354259 457131 354325 457132
rect 353155 457060 353221 457061
rect 353155 456996 353156 457060
rect 353220 456996 353221 457060
rect 353155 456995 353221 456996
rect 350947 456924 351013 456925
rect 350947 456860 350948 456924
rect 351012 456860 351013 456924
rect 350947 456859 351013 456860
rect 351867 456924 351933 456925
rect 351867 456860 351868 456924
rect 351932 456860 351933 456924
rect 351867 456859 351933 456860
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 427254 354204 457000
rect 355366 456925 355426 459310
rect 356470 458013 356530 459310
rect 356467 458012 356533 458013
rect 356467 457948 356468 458012
rect 356532 457948 356533 458012
rect 356467 457947 356533 457948
rect 356654 456925 356714 459310
rect 357390 457741 357450 460670
rect 357806 459370 357866 460020
rect 358850 459509 358910 460020
rect 358847 459508 358913 459509
rect 358847 459444 358848 459508
rect 358912 459444 358913 459508
rect 358847 459443 358913 459444
rect 358974 459370 359034 460020
rect 357758 459310 357866 459370
rect 358862 459310 359034 459370
rect 357387 457740 357453 457741
rect 357387 457676 357388 457740
rect 357452 457676 357453 457740
rect 357387 457675 357453 457676
rect 357758 456925 357818 459310
rect 358862 456925 358922 459310
rect 355363 456924 355429 456925
rect 355363 456860 355364 456924
rect 355428 456860 355429 456924
rect 355363 456859 355429 456860
rect 356651 456924 356717 456925
rect 356651 456860 356652 456924
rect 356716 456860 356717 456924
rect 356651 456859 356717 456860
rect 357755 456924 357821 456925
rect 357755 456860 357756 456924
rect 357820 456860 357821 456924
rect 357755 456859 357821 456860
rect 358859 456924 358925 456925
rect 358859 456860 358860 456924
rect 358924 456860 358925 456924
rect 358859 456859 358925 456860
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 434454 361404 457000
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 438054 365004 457000
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 441654 368604 457000
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 445254 372204 457000
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 452454 379404 457000
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 456054 383004 457000
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 423654 386604 457000
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 427254 390204 457000
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 434667 626924 434733 626925
rect 434667 626860 434668 626924
rect 434732 626860 434733 626924
rect 434667 626859 434733 626860
rect 434670 626653 434730 626859
rect 434667 626652 434733 626653
rect 434667 626588 434668 626652
rect 434732 626588 434733 626652
rect 434667 626587 434733 626588
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 434667 603260 434733 603261
rect 434667 603196 434668 603260
rect 434732 603196 434733 603260
rect 434667 603195 434733 603196
rect 434670 602989 434730 603195
rect 434667 602988 434733 602989
rect 434667 602924 434668 602988
rect 434732 602924 434733 602988
rect 434667 602923 434733 602924
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 554247 437004 581498
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 554247 440604 585098
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 554247 444204 588698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 554247 451404 559898
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 554247 455004 563498
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 554247 458604 567098
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 554247 462204 570698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 554247 469404 577898
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 554247 473004 581498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 554247 476604 585098
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 554247 480204 588698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 554247 487404 559898
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 554247 491004 563498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 554247 494604 567098
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 554247 498204 570698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 554247 505404 577898
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 554247 509004 581498
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 554247 512604 585098
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 554247 516204 588698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 507899 553484 507965 553485
rect 507899 553420 507900 553484
rect 507964 553420 507965 553484
rect 507899 553419 507965 553420
rect 513419 553484 513485 553485
rect 513419 553420 513420 553484
rect 513484 553420 513485 553484
rect 513419 553419 513485 553420
rect 507902 551170 507962 553419
rect 513422 551170 513482 553419
rect 507902 551110 508608 551170
rect 513422 551110 514218 551170
rect 514158 550765 514218 551110
rect 514155 550764 514221 550765
rect 514155 550700 514156 550764
rect 514220 550700 514221 550764
rect 514155 550699 514221 550700
rect 516494 546054 516814 546076
rect 516494 545818 516536 546054
rect 516772 545818 516814 546054
rect 516494 545734 516814 545818
rect 516494 545498 516536 545734
rect 516772 545498 516814 545734
rect 516494 545476 516814 545498
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 516494 542454 516814 542476
rect 516494 542218 516536 542454
rect 516772 542218 516814 542454
rect 516494 542134 516814 542218
rect 516494 541898 516536 542134
rect 516772 541898 516814 542134
rect 516494 541876 516814 541898
rect 516938 535254 517262 535276
rect 516938 535018 516982 535254
rect 517218 535018 517262 535254
rect 516938 534934 517262 535018
rect 516938 534698 516982 534934
rect 517218 534698 517262 534934
rect 516938 534676 517262 534698
rect 516938 531654 517262 531676
rect 516938 531418 516982 531654
rect 517218 531418 517262 531654
rect 516938 531334 517262 531418
rect 516938 531098 516982 531334
rect 517218 531098 517262 531334
rect 516938 531076 517262 531098
rect 516938 528054 517262 528076
rect 516938 527818 516982 528054
rect 517218 527818 517262 528054
rect 516938 527734 517262 527818
rect 516938 527498 516982 527734
rect 517218 527498 517262 527734
rect 516938 527476 517262 527498
rect 516938 524454 517262 524476
rect 516938 524218 516982 524454
rect 517218 524218 517262 524454
rect 516938 524134 517262 524218
rect 516938 523898 516982 524134
rect 517218 523898 517262 524134
rect 516938 523876 517262 523898
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 516494 517254 516814 517276
rect 516494 517018 516536 517254
rect 516772 517018 516814 517254
rect 516494 516934 516814 517018
rect 516494 516698 516536 516934
rect 516772 516698 516814 516934
rect 516494 516676 516814 516698
rect 516494 513654 516814 513676
rect 516494 513418 516536 513654
rect 516772 513418 516814 513654
rect 516494 513334 516814 513418
rect 516494 513098 516536 513334
rect 516772 513098 516814 513334
rect 516494 513076 516814 513098
rect 516494 510054 516814 510076
rect 516494 509818 516536 510054
rect 516772 509818 516814 510054
rect 516494 509734 516814 509818
rect 516494 509498 516536 509734
rect 516772 509498 516814 509734
rect 516494 509476 516814 509498
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 516494 506454 516814 506476
rect 516494 506218 516536 506454
rect 516772 506218 516814 506454
rect 516494 506134 516814 506218
rect 516494 505898 516536 506134
rect 516772 505898 516814 506134
rect 516494 505876 516814 505898
rect 516938 499254 517262 499276
rect 516938 499018 516982 499254
rect 517218 499018 517262 499254
rect 516938 498934 517262 499018
rect 516938 498698 516982 498934
rect 517218 498698 517262 498934
rect 516938 498676 517262 498698
rect 516938 495654 517262 495676
rect 516938 495418 516982 495654
rect 517218 495418 517262 495654
rect 516938 495334 517262 495418
rect 516938 495098 516982 495334
rect 517218 495098 517262 495334
rect 516938 495076 517262 495098
rect 516938 492054 517262 492076
rect 516938 491818 516982 492054
rect 517218 491818 517262 492054
rect 516938 491734 517262 491818
rect 516938 491498 516982 491734
rect 517218 491498 517262 491734
rect 516938 491476 517262 491498
rect 516938 488454 517262 488476
rect 516938 488218 516982 488454
rect 517218 488218 517262 488454
rect 516938 488134 517262 488218
rect 516938 487898 516982 488134
rect 517218 487898 517262 488134
rect 516938 487876 517262 487898
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 516494 481254 516814 481276
rect 516494 481018 516536 481254
rect 516772 481018 516814 481254
rect 516494 480934 516814 481018
rect 516494 480698 516536 480934
rect 516772 480698 516814 480934
rect 516494 480676 516814 480698
rect 516494 477654 516814 477676
rect 516494 477418 516536 477654
rect 516772 477418 516814 477654
rect 516494 477334 516814 477418
rect 516494 477098 516536 477334
rect 516772 477098 516814 477334
rect 516494 477076 516814 477098
rect 516494 474054 516814 474076
rect 516494 473818 516536 474054
rect 516772 473818 516814 474054
rect 516494 473734 516814 473818
rect 516494 473498 516536 473734
rect 516772 473498 516814 473734
rect 516494 473476 516814 473498
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 516494 470454 516814 470476
rect 516494 470218 516536 470454
rect 516772 470218 516814 470454
rect 516494 470134 516814 470218
rect 516494 469898 516536 470134
rect 516772 469898 516814 470134
rect 516494 469876 516814 469898
rect 516938 463254 517262 463276
rect 516938 463018 516982 463254
rect 517218 463018 517262 463254
rect 516938 462934 517262 463018
rect 516938 462698 516982 462934
rect 517218 462698 517262 462934
rect 516938 462676 517262 462698
rect 454726 460670 455008 460730
rect 458222 460670 458512 460730
rect 461718 460670 462016 460730
rect 465214 460670 465520 460730
rect 468710 460670 469024 460730
rect 472206 460670 472528 460730
rect 481590 460670 481872 460730
rect 443134 460330 443833 460390
rect 448470 460330 449168 460390
rect 453622 460330 453840 460390
rect 443134 458013 443194 460330
rect 446802 459370 446862 460020
rect 447970 459370 448030 460020
rect 446802 459310 446874 459370
rect 443131 458012 443197 458013
rect 443131 457948 443132 458012
rect 443196 457948 443197 458012
rect 443131 457947 443197 457948
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 438054 437004 457000
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 441654 440604 457000
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 445254 444204 457000
rect 446814 456925 446874 459310
rect 447918 459310 448030 459370
rect 447918 457061 447978 459310
rect 447915 457060 447981 457061
rect 447915 456996 447916 457060
rect 447980 456996 447981 457060
rect 447915 456995 447981 456996
rect 448470 456925 448530 460330
rect 450306 459370 450366 460020
rect 451474 459370 451534 460020
rect 452642 459509 452702 460020
rect 452639 459508 452705 459509
rect 452639 459444 452640 459508
rect 452704 459444 452705 459508
rect 452639 459443 452705 459444
rect 452766 459370 452826 460020
rect 453067 459508 453133 459509
rect 453067 459444 453068 459508
rect 453132 459444 453133 459508
rect 453067 459443 453133 459444
rect 450306 459310 450370 459370
rect 450310 456925 450370 459310
rect 451414 459310 451534 459370
rect 452702 459310 452826 459370
rect 451414 457197 451474 459310
rect 451411 457196 451477 457197
rect 451411 457132 451412 457196
rect 451476 457132 451477 457196
rect 451411 457131 451477 457132
rect 446811 456924 446877 456925
rect 446811 456860 446812 456924
rect 446876 456860 446877 456924
rect 446811 456859 446877 456860
rect 448467 456924 448533 456925
rect 448467 456860 448468 456924
rect 448532 456860 448533 456924
rect 448467 456859 448533 456860
rect 450307 456924 450373 456925
rect 450307 456860 450308 456924
rect 450372 456860 450373 456924
rect 450307 456859 450373 456860
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 452454 451404 457000
rect 452702 456925 452762 459310
rect 453070 456925 453130 459443
rect 453622 456925 453682 460330
rect 453934 459370 453994 460020
rect 453806 459310 453994 459370
rect 453806 457469 453866 459310
rect 453803 457468 453869 457469
rect 453803 457404 453804 457468
rect 453868 457404 453869 457468
rect 453803 457403 453869 457404
rect 454726 457197 454786 460670
rect 456014 460330 456176 460390
rect 455102 459370 455162 460020
rect 455094 459310 455162 459370
rect 455094 457469 455154 459310
rect 455091 457468 455157 457469
rect 455091 457404 455092 457468
rect 455156 457404 455157 457468
rect 455091 457403 455157 457404
rect 454723 457196 454789 457197
rect 454723 457132 454724 457196
rect 454788 457132 454789 457196
rect 454723 457131 454789 457132
rect 456014 457061 456074 460330
rect 456270 459370 456330 460020
rect 457314 459370 457374 460020
rect 456198 459310 456330 459370
rect 457302 459310 457374 459370
rect 457438 459370 457498 460020
rect 457438 459310 457546 459370
rect 456011 457060 456077 457061
rect 452699 456924 452765 456925
rect 452699 456860 452700 456924
rect 452764 456860 452765 456924
rect 452699 456859 452765 456860
rect 453067 456924 453133 456925
rect 453067 456860 453068 456924
rect 453132 456860 453133 456924
rect 453067 456859 453133 456860
rect 453619 456924 453685 456925
rect 453619 456860 453620 456924
rect 453684 456860 453685 456924
rect 453619 456859 453685 456860
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 456054 455004 457000
rect 456011 456996 456012 457060
rect 456076 456996 456077 457060
rect 456011 456995 456077 456996
rect 456198 456925 456258 459310
rect 457302 456925 457362 459310
rect 457486 457605 457546 459310
rect 457483 457604 457549 457605
rect 457483 457540 457484 457604
rect 457548 457540 457549 457604
rect 457483 457539 457549 457540
rect 458222 457197 458282 460670
rect 459510 460330 459680 460390
rect 458606 459370 458666 460020
rect 458590 459310 458666 459370
rect 458590 457877 458650 459310
rect 459510 458013 459570 460330
rect 459774 459370 459834 460020
rect 460818 459370 460878 460020
rect 459694 459310 459834 459370
rect 460798 459310 460878 459370
rect 460942 459370 461002 460020
rect 460942 459310 461042 459370
rect 459507 458012 459573 458013
rect 459507 457948 459508 458012
rect 459572 457948 459573 458012
rect 459507 457947 459573 457948
rect 458587 457876 458653 457877
rect 458587 457812 458588 457876
rect 458652 457812 458653 457876
rect 458587 457811 458653 457812
rect 459694 457605 459754 459310
rect 460798 457741 460858 459310
rect 460795 457740 460861 457741
rect 460795 457676 460796 457740
rect 460860 457676 460861 457740
rect 460795 457675 460861 457676
rect 459691 457604 459757 457605
rect 459691 457540 459692 457604
rect 459756 457540 459757 457604
rect 459691 457539 459757 457540
rect 458219 457196 458285 457197
rect 458219 457132 458220 457196
rect 458284 457132 458285 457196
rect 458219 457131 458285 457132
rect 456195 456924 456261 456925
rect 456195 456860 456196 456924
rect 456260 456860 456261 456924
rect 456195 456859 456261 456860
rect 457299 456924 457365 456925
rect 457299 456860 457300 456924
rect 457364 456860 457365 456924
rect 457299 456859 457365 456860
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 423654 458604 457000
rect 460982 456925 461042 459310
rect 461718 458149 461778 460670
rect 463006 460330 463184 460390
rect 462110 459370 462170 460020
rect 462086 459310 462170 459370
rect 461715 458148 461781 458149
rect 461715 458084 461716 458148
rect 461780 458084 461781 458148
rect 461715 458083 461781 458084
rect 462086 457197 462146 459310
rect 463006 458149 463066 460330
rect 463278 459370 463338 460020
rect 464322 459370 464382 460020
rect 463190 459310 463338 459370
rect 464294 459310 464382 459370
rect 464446 459370 464506 460020
rect 464446 459310 464538 459370
rect 463003 458148 463069 458149
rect 463003 458084 463004 458148
rect 463068 458084 463069 458148
rect 463003 458083 463069 458084
rect 462083 457196 462149 457197
rect 462083 457132 462084 457196
rect 462148 457132 462149 457196
rect 462083 457131 462149 457132
rect 460979 456924 461045 456925
rect 460979 456860 460980 456924
rect 461044 456860 461045 456924
rect 460979 456859 461045 456860
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 427254 462204 457000
rect 463190 456925 463250 459310
rect 464294 458149 464354 459310
rect 464291 458148 464357 458149
rect 464291 458084 464292 458148
rect 464356 458084 464357 458148
rect 464291 458083 464357 458084
rect 464478 456925 464538 459310
rect 465214 458149 465274 460670
rect 466502 460330 466688 460390
rect 465614 459370 465674 460020
rect 465582 459310 465674 459370
rect 465211 458148 465277 458149
rect 465211 458084 465212 458148
rect 465276 458084 465277 458148
rect 465211 458083 465277 458084
rect 465582 456925 465642 459310
rect 466502 457877 466562 460330
rect 466782 459370 466842 460020
rect 467826 459370 467886 460020
rect 466686 459310 466842 459370
rect 467790 459310 467886 459370
rect 467950 459370 468010 460020
rect 467950 459310 468034 459370
rect 466499 457876 466565 457877
rect 466499 457812 466500 457876
rect 466564 457812 466565 457876
rect 466499 457811 466565 457812
rect 466686 456925 466746 459310
rect 467790 458013 467850 459310
rect 467787 458012 467853 458013
rect 467787 457948 467788 458012
rect 467852 457948 467853 458012
rect 467787 457947 467853 457948
rect 467974 456925 468034 459310
rect 468710 458149 468770 460670
rect 469998 460330 470192 460390
rect 469118 459370 469178 460020
rect 469078 459310 469178 459370
rect 468707 458148 468773 458149
rect 468707 458084 468708 458148
rect 468772 458084 468773 458148
rect 468707 458083 468773 458084
rect 469078 457197 469138 459310
rect 469998 458149 470058 460330
rect 470286 459370 470346 460020
rect 471330 459370 471390 460020
rect 470182 459310 470346 459370
rect 471286 459310 471390 459370
rect 471454 459370 471514 460020
rect 471454 459310 471530 459370
rect 469995 458148 470061 458149
rect 469995 458084 469996 458148
rect 470060 458084 470061 458148
rect 469995 458083 470061 458084
rect 469075 457196 469141 457197
rect 469075 457132 469076 457196
rect 469140 457132 469141 457196
rect 469075 457131 469141 457132
rect 463187 456924 463253 456925
rect 463187 456860 463188 456924
rect 463252 456860 463253 456924
rect 463187 456859 463253 456860
rect 464475 456924 464541 456925
rect 464475 456860 464476 456924
rect 464540 456860 464541 456924
rect 464475 456859 464541 456860
rect 465579 456924 465645 456925
rect 465579 456860 465580 456924
rect 465644 456860 465645 456924
rect 465579 456859 465645 456860
rect 466683 456924 466749 456925
rect 466683 456860 466684 456924
rect 466748 456860 466749 456924
rect 466683 456859 466749 456860
rect 467971 456924 468037 456925
rect 467971 456860 467972 456924
rect 468036 456860 468037 456924
rect 467971 456859 468037 456860
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 434454 469404 457000
rect 470182 456925 470242 459310
rect 471286 458149 471346 459310
rect 471283 458148 471349 458149
rect 471283 458084 471284 458148
rect 471348 458084 471349 458148
rect 471283 458083 471349 458084
rect 471470 456925 471530 459310
rect 472206 458149 472266 460670
rect 473494 460330 473696 460390
rect 475518 460330 476032 460390
rect 476990 460330 477200 460390
rect 479382 460330 479536 460390
rect 472622 459370 472682 460020
rect 472574 459310 472682 459370
rect 472203 458148 472269 458149
rect 472203 458084 472204 458148
rect 472268 458084 472269 458148
rect 472203 458083 472269 458084
rect 472574 457197 472634 459310
rect 473494 458149 473554 460330
rect 473790 459370 473850 460020
rect 474834 459370 474894 460020
rect 473678 459310 473850 459370
rect 474782 459310 474894 459370
rect 474958 459370 475018 460020
rect 474958 459310 475026 459370
rect 473491 458148 473557 458149
rect 473491 458084 473492 458148
rect 473556 458084 473557 458148
rect 473491 458083 473557 458084
rect 472571 457196 472637 457197
rect 472571 457132 472572 457196
rect 472636 457132 472637 457196
rect 472571 457131 472637 457132
rect 470179 456924 470245 456925
rect 470179 456860 470180 456924
rect 470244 456860 470245 456924
rect 470179 456859 470245 456860
rect 471467 456924 471533 456925
rect 471467 456860 471468 456924
rect 471532 456860 471533 456924
rect 471467 456859 471533 456860
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 438054 473004 457000
rect 473678 456925 473738 459310
rect 474782 458149 474842 459310
rect 474779 458148 474845 458149
rect 474779 458084 474780 458148
rect 474844 458084 474845 458148
rect 474779 458083 474845 458084
rect 474966 456925 475026 459310
rect 475518 458149 475578 460330
rect 476126 459370 476186 460020
rect 476070 459310 476186 459370
rect 475515 458148 475581 458149
rect 475515 458084 475516 458148
rect 475580 458084 475581 458148
rect 475515 458083 475581 458084
rect 476070 457197 476130 459310
rect 476990 458149 477050 460330
rect 477294 459370 477354 460020
rect 478338 459370 478398 460020
rect 477174 459310 477354 459370
rect 478278 459310 478398 459370
rect 476987 458148 477053 458149
rect 476987 458084 476988 458148
rect 477052 458084 477053 458148
rect 476987 458083 477053 458084
rect 477174 457333 477234 459310
rect 478278 458149 478338 459310
rect 478275 458148 478341 458149
rect 478275 458084 478276 458148
rect 478340 458084 478341 458148
rect 478275 458083 478341 458084
rect 478462 457333 478522 460020
rect 479382 458149 479442 460330
rect 479630 459370 479690 460020
rect 480674 459370 480734 460020
rect 479566 459310 479690 459370
rect 480670 459310 480734 459370
rect 480798 459370 480858 460020
rect 480798 459310 480914 459370
rect 479379 458148 479445 458149
rect 479379 458084 479380 458148
rect 479444 458084 479445 458148
rect 479379 458083 479445 458084
rect 479566 457877 479626 459310
rect 480670 458013 480730 459310
rect 480667 458012 480733 458013
rect 480667 457948 480668 458012
rect 480732 457948 480733 458012
rect 480667 457947 480733 457948
rect 480854 457877 480914 459310
rect 479563 457876 479629 457877
rect 479563 457812 479564 457876
rect 479628 457812 479629 457876
rect 479563 457811 479629 457812
rect 480851 457876 480917 457877
rect 480851 457812 480852 457876
rect 480916 457812 480917 457876
rect 480851 457811 480917 457812
rect 481590 457741 481650 460670
rect 483614 460330 484208 460390
rect 484718 460330 485376 460390
rect 486006 460330 486544 460390
rect 488582 460330 488880 460390
rect 481966 459370 482026 460020
rect 483010 459509 483070 460020
rect 483007 459508 483073 459509
rect 483007 459444 483008 459508
rect 483072 459444 483073 459508
rect 483007 459443 483073 459444
rect 483134 459370 483194 460020
rect 481958 459310 482026 459370
rect 483062 459310 483194 459370
rect 481587 457740 481653 457741
rect 481587 457676 481588 457740
rect 481652 457676 481653 457740
rect 481587 457675 481653 457676
rect 477171 457332 477237 457333
rect 477171 457268 477172 457332
rect 477236 457268 477237 457332
rect 477171 457267 477237 457268
rect 478459 457332 478525 457333
rect 478459 457268 478460 457332
rect 478524 457268 478525 457332
rect 478459 457267 478525 457268
rect 481958 457197 482018 459310
rect 483062 458149 483122 459310
rect 483059 458148 483125 458149
rect 483059 458084 483060 458148
rect 483124 458084 483125 458148
rect 483059 458083 483125 458084
rect 483614 457469 483674 460330
rect 484302 459370 484362 460020
rect 484166 459310 484362 459370
rect 484166 458149 484226 459310
rect 484163 458148 484229 458149
rect 484163 458084 484164 458148
rect 484228 458084 484229 458148
rect 484163 458083 484229 458084
rect 484718 457877 484778 460330
rect 485470 459370 485530 460020
rect 485454 459310 485530 459370
rect 485454 458149 485514 459310
rect 485451 458148 485517 458149
rect 485451 458084 485452 458148
rect 485516 458084 485517 458148
rect 485451 458083 485517 458084
rect 484715 457876 484781 457877
rect 484715 457812 484716 457876
rect 484780 457812 484781 457876
rect 484715 457811 484781 457812
rect 486006 457741 486066 460330
rect 486638 459370 486698 460020
rect 487682 459370 487742 460020
rect 486558 459310 486698 459370
rect 487662 459310 487742 459370
rect 487806 459370 487866 460020
rect 487806 459310 487906 459370
rect 486003 457740 486069 457741
rect 486003 457676 486004 457740
rect 486068 457676 486069 457740
rect 486003 457675 486069 457676
rect 486558 457469 486618 459310
rect 487662 458013 487722 459310
rect 487659 458012 487725 458013
rect 487659 457948 487660 458012
rect 487724 457948 487725 458012
rect 487659 457947 487725 457948
rect 487846 457605 487906 459310
rect 488582 457741 488642 460330
rect 488974 459370 489034 460020
rect 488950 459310 489034 459370
rect 488579 457740 488645 457741
rect 488579 457676 488580 457740
rect 488644 457676 488645 457740
rect 488579 457675 488645 457676
rect 487843 457604 487909 457605
rect 487843 457540 487844 457604
rect 487908 457540 487909 457604
rect 487843 457539 487909 457540
rect 488950 457469 489010 459310
rect 483611 457468 483677 457469
rect 483611 457404 483612 457468
rect 483676 457404 483677 457468
rect 483611 457403 483677 457404
rect 486555 457468 486621 457469
rect 486555 457404 486556 457468
rect 486620 457404 486621 457468
rect 486555 457403 486621 457404
rect 488947 457468 489013 457469
rect 488947 457404 488948 457468
rect 489012 457404 489013 457468
rect 488947 457403 489013 457404
rect 476067 457196 476133 457197
rect 476067 457132 476068 457196
rect 476132 457132 476133 457196
rect 476067 457131 476133 457132
rect 481955 457196 482021 457197
rect 481955 457132 481956 457196
rect 482020 457132 482021 457196
rect 481955 457131 482021 457132
rect 473675 456924 473741 456925
rect 473675 456860 473676 456924
rect 473740 456860 473741 456924
rect 473675 456859 473741 456860
rect 474963 456924 475029 456925
rect 474963 456860 474964 456924
rect 475028 456860 475029 456924
rect 474963 456859 475029 456860
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 441654 476604 457000
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 445254 480204 457000
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 452454 487404 457000
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 456054 491004 457000
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 423654 494604 457000
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 427254 498204 457000
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 434454 505404 457000
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 438054 509004 457000
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 441654 512604 457000
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 445254 516204 457000
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 550587 673980 550653 673981
rect 550587 673916 550588 673980
rect 550652 673916 550653 673980
rect 550587 673915 550653 673916
rect 550590 673573 550650 673915
rect 550587 673572 550653 673573
rect 550587 673508 550588 673572
rect 550652 673508 550653 673572
rect 550587 673507 550653 673508
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 550587 650452 550653 650453
rect 550587 650388 550588 650452
rect 550652 650388 550653 650452
rect 550587 650387 550653 650388
rect 550590 650045 550650 650387
rect 550587 650044 550653 650045
rect 550587 649980 550588 650044
rect 550652 649980 550653 650044
rect 550587 649979 550653 649980
rect 550587 627060 550653 627061
rect 550587 626996 550588 627060
rect 550652 626996 550653 627060
rect 550587 626995 550653 626996
rect 550590 626653 550650 626995
rect 550587 626652 550653 626653
rect 550587 626588 550588 626652
rect 550652 626588 550653 626652
rect 550587 626587 550653 626588
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 136536 545818 136772 546054
rect 136536 545498 136772 545734
rect 136536 542218 136772 542454
rect 136536 541898 136772 542134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 136982 535018 137218 535254
rect 136982 534698 137218 534934
rect 136982 531418 137218 531654
rect 136982 531098 137218 531334
rect 136982 527818 137218 528054
rect 136982 527498 137218 527734
rect 136982 524218 137218 524454
rect 136982 523898 137218 524134
rect 136536 517018 136772 517254
rect 136536 516698 136772 516934
rect 136536 513418 136772 513654
rect 136536 513098 136772 513334
rect 136536 509818 136772 510054
rect 136536 509498 136772 509734
rect 136536 506218 136772 506454
rect 136536 505898 136772 506134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 136982 499018 137218 499254
rect 136982 498698 137218 498934
rect 136982 495418 137218 495654
rect 136982 495098 137218 495334
rect 136982 491818 137218 492054
rect 136982 491498 137218 491734
rect 136982 488218 137218 488454
rect 136982 487898 137218 488134
rect 136536 481018 136772 481254
rect 136536 480698 136772 480934
rect 136536 477418 136772 477654
rect 136536 477098 136772 477334
rect 136536 473818 136772 474054
rect 136536 473498 136772 473734
rect 136536 470218 136772 470454
rect 136536 469898 136772 470134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 136982 463018 137218 463254
rect 136982 462698 137218 462934
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 266536 545818 266772 546054
rect 266536 545498 266772 545734
rect 266536 542218 266772 542454
rect 266536 541898 266772 542134
rect 266982 535018 267218 535254
rect 266982 534698 267218 534934
rect 266982 531418 267218 531654
rect 266982 531098 267218 531334
rect 266982 527818 267218 528054
rect 266982 527498 267218 527734
rect 266982 524218 267218 524454
rect 266982 523898 267218 524134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 266536 517018 266772 517254
rect 266536 516698 266772 516934
rect 266536 513418 266772 513654
rect 266536 513098 266772 513334
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 266536 509818 266772 510054
rect 266536 509498 266772 509734
rect 266536 506218 266772 506454
rect 266536 505898 266772 506134
rect 266982 499018 267218 499254
rect 266982 498698 267218 498934
rect 266982 495418 267218 495654
rect 266982 495098 267218 495334
rect 266982 491818 267218 492054
rect 266982 491498 267218 491734
rect 266982 488218 267218 488454
rect 266982 487898 267218 488134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 266536 481018 266772 481254
rect 266536 480698 266772 480934
rect 266536 477418 266772 477654
rect 266536 477098 266772 477334
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 266536 473818 266772 474054
rect 266536 473498 266772 473734
rect 266536 470218 266772 470454
rect 266536 469898 266772 470134
rect 266982 463018 267218 463254
rect 266982 462698 267218 462934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 386536 545818 386772 546054
rect 386536 545498 386772 545734
rect 386536 542218 386772 542454
rect 386536 541898 386772 542134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 386982 535018 387218 535254
rect 386982 534698 387218 534934
rect 386982 531418 387218 531654
rect 386982 531098 387218 531334
rect 386982 527818 387218 528054
rect 386982 527498 387218 527734
rect 386982 524218 387218 524454
rect 386982 523898 387218 524134
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 386536 517018 386772 517254
rect 386536 516698 386772 516934
rect 386536 513418 386772 513654
rect 386536 513098 386772 513334
rect 386536 509818 386772 510054
rect 386536 509498 386772 509734
rect 386536 506218 386772 506454
rect 386536 505898 386772 506134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 386982 499018 387218 499254
rect 386982 498698 387218 498934
rect 386982 495418 387218 495654
rect 386982 495098 387218 495334
rect 386982 491818 387218 492054
rect 386982 491498 387218 491734
rect 386982 488218 387218 488454
rect 386982 487898 387218 488134
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 386536 481018 386772 481254
rect 386536 480698 386772 480934
rect 386536 477418 386772 477654
rect 386536 477098 386772 477334
rect 386536 473818 386772 474054
rect 386536 473498 386772 473734
rect 386536 470218 386772 470454
rect 386536 469898 386772 470134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 386982 463018 387218 463254
rect 386982 462698 387218 462934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 64250 434218 64486 434454
rect 64250 433898 64486 434134
rect 79610 427018 79846 427254
rect 79610 426698 79846 426934
rect 79610 423418 79846 423654
rect 79610 423098 79846 423334
rect 79610 419818 79846 420054
rect 79610 419498 79846 419734
rect 79610 416218 79846 416454
rect 79610 415898 79846 416134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 64250 409018 64486 409254
rect 64250 408698 64486 408934
rect 64250 405418 64486 405654
rect 64250 405098 64486 405334
rect 64250 401818 64486 402054
rect 64250 401498 64486 401734
rect 64250 398218 64486 398454
rect 64250 397898 64486 398134
rect 79610 391018 79846 391254
rect 79610 390698 79846 390934
rect 79610 387418 79846 387654
rect 79610 387098 79846 387334
rect 79610 383818 79846 384054
rect 79610 383498 79846 383734
rect 79610 380218 79846 380454
rect 79610 379898 79846 380134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 64250 373018 64486 373254
rect 64250 372698 64486 372934
rect 64250 369418 64486 369654
rect 64250 369098 64486 369334
rect 64250 365818 64486 366054
rect 64250 365498 64486 365734
rect 64250 362218 64486 362454
rect 64250 361898 64486 362134
rect 79610 355018 79846 355254
rect 79610 354698 79846 354934
rect 79610 351418 79846 351654
rect 79610 351098 79846 351334
rect 79610 347818 79846 348054
rect 79610 347498 79846 347734
rect 79610 344218 79846 344454
rect 79610 343898 79846 344134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 64250 337018 64486 337254
rect 64250 336698 64486 336934
rect 64250 333418 64486 333654
rect 64250 333098 64486 333334
rect 64250 329818 64486 330054
rect 64250 329498 64486 329734
rect 64250 326218 64486 326454
rect 64250 325898 64486 326134
rect 79610 319018 79846 319254
rect 79610 318698 79846 318934
rect 79610 315418 79846 315654
rect 79610 315098 79846 315334
rect 79610 311818 79846 312054
rect 79610 311498 79846 311734
rect 79610 308218 79846 308454
rect 79610 307898 79846 308134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 64250 301018 64486 301254
rect 64250 300698 64486 300934
rect 64250 297418 64486 297654
rect 64250 297098 64486 297334
rect 64250 293818 64486 294054
rect 64250 293498 64486 293734
rect 64250 290218 64486 290454
rect 64250 289898 64486 290134
rect 79610 283018 79846 283254
rect 79610 282698 79846 282934
rect 79610 279418 79846 279654
rect 79610 279098 79846 279334
rect 79610 275818 79846 276054
rect 79610 275498 79846 275734
rect 79610 272218 79846 272454
rect 79610 271898 79846 272134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 64250 265018 64486 265254
rect 64250 264698 64486 264934
rect 64250 261418 64486 261654
rect 64250 261098 64486 261334
rect 64250 257818 64486 258054
rect 64250 257498 64486 257734
rect 64250 254218 64486 254454
rect 64250 253898 64486 254134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 79610 247018 79846 247254
rect 79610 246698 79846 246934
rect 79610 243418 79846 243654
rect 79610 243098 79846 243334
rect 79610 239818 79846 240054
rect 79610 239498 79846 239734
rect 79610 236218 79846 236454
rect 79610 235898 79846 236134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 64250 229018 64486 229254
rect 64250 228698 64486 228934
rect 64250 225418 64486 225654
rect 64250 225098 64486 225334
rect 64250 221818 64486 222054
rect 64250 221498 64486 221734
rect 64250 218218 64486 218454
rect 64250 217898 64486 218134
rect 79610 211018 79846 211254
rect 79610 210698 79846 210934
rect 79610 207418 79846 207654
rect 79610 207098 79846 207334
rect 79610 203818 79846 204054
rect 79610 203498 79846 203734
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 516536 545818 516772 546054
rect 516536 545498 516772 545734
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 516536 542218 516772 542454
rect 516536 541898 516772 542134
rect 516982 535018 517218 535254
rect 516982 534698 517218 534934
rect 516982 531418 517218 531654
rect 516982 531098 517218 531334
rect 516982 527818 517218 528054
rect 516982 527498 517218 527734
rect 516982 524218 517218 524454
rect 516982 523898 517218 524134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 516536 517018 516772 517254
rect 516536 516698 516772 516934
rect 516536 513418 516772 513654
rect 516536 513098 516772 513334
rect 516536 509818 516772 510054
rect 516536 509498 516772 509734
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 516536 506218 516772 506454
rect 516536 505898 516772 506134
rect 516982 499018 517218 499254
rect 516982 498698 517218 498934
rect 516982 495418 517218 495654
rect 516982 495098 517218 495334
rect 516982 491818 517218 492054
rect 516982 491498 517218 491734
rect 516982 488218 517218 488454
rect 516982 487898 517218 488134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 516536 481018 516772 481254
rect 516536 480698 516772 480934
rect 516536 477418 516772 477654
rect 516536 477098 516772 477334
rect 516536 473818 516772 474054
rect 516536 473498 516772 473734
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 516536 470218 516772 470454
rect 516536 469898 516772 470134
rect 516982 463018 517218 463254
rect 516982 462698 517218 462934
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 155604 553276 156204 553278
rect 299604 553276 300204 553278
rect 407604 553276 408204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 155786 553254
rect 156022 553018 299786 553254
rect 300022 553018 407786 553254
rect 408022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 155786 552934
rect 156022 552698 299786 552934
rect 300022 552698 407786 552934
rect 408022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 155604 552674 156204 552676
rect 299604 552674 300204 552676
rect 407604 552674 408204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 152004 549676 152604 549678
rect 296004 549676 296604 549678
rect 404004 549676 404604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 152186 549654
rect 152422 549418 296186 549654
rect 296422 549418 404186 549654
rect 404422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 152186 549334
rect 152422 549098 296186 549334
rect 296422 549098 404186 549334
rect 404422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 152004 549074 152604 549076
rect 296004 549074 296604 549076
rect 404004 549074 404604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 136494 546076 136814 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 266494 546076 266814 546078
rect 292404 546076 293004 546078
rect 386494 546076 386814 546078
rect 400404 546076 401004 546078
rect 516494 546076 516814 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 136536 546054
rect 136772 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 266536 546054
rect 266772 545818 292586 546054
rect 292822 545818 386536 546054
rect 386772 545818 400586 546054
rect 400822 545818 516536 546054
rect 516772 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 136536 545734
rect 136772 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 266536 545734
rect 266772 545498 292586 545734
rect 292822 545498 386536 545734
rect 386772 545498 400586 545734
rect 400822 545498 516536 545734
rect 516772 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 136494 545474 136814 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 266494 545474 266814 545476
rect 292404 545474 293004 545476
rect 386494 545474 386814 545476
rect 400404 545474 401004 545476
rect 516494 545474 516814 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 136494 542476 136814 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 266494 542476 266814 542478
rect 288804 542476 289404 542478
rect 386494 542476 386814 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 516494 542476 516814 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 136536 542454
rect 136772 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 266536 542454
rect 266772 542218 288986 542454
rect 289222 542218 386536 542454
rect 386772 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 516536 542454
rect 516772 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 136536 542134
rect 136772 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 266536 542134
rect 266772 541898 288986 542134
rect 289222 541898 386536 542134
rect 386772 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 516536 542134
rect 516772 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 136494 541874 136814 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 266494 541874 266814 541876
rect 288804 541874 289404 541876
rect 386494 541874 386814 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 516494 541874 516814 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 136938 535276 137262 535278
rect 173604 535276 174204 535278
rect 266938 535276 267262 535278
rect 281604 535276 282204 535278
rect 386938 535276 387262 535278
rect 425604 535276 426204 535278
rect 516938 535276 517262 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 136982 535254
rect 137218 535018 173786 535254
rect 174022 535018 266982 535254
rect 267218 535018 281786 535254
rect 282022 535018 386982 535254
rect 387218 535018 425786 535254
rect 426022 535018 516982 535254
rect 517218 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 136982 534934
rect 137218 534698 173786 534934
rect 174022 534698 266982 534934
rect 267218 534698 281786 534934
rect 282022 534698 386982 534934
rect 387218 534698 425786 534934
rect 426022 534698 516982 534934
rect 517218 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 136938 534674 137262 534676
rect 173604 534674 174204 534676
rect 266938 534674 267262 534676
rect 281604 534674 282204 534676
rect 386938 534674 387262 534676
rect 425604 534674 426204 534676
rect 516938 534674 517262 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 136938 531676 137262 531678
rect 170004 531676 170604 531678
rect 266938 531676 267262 531678
rect 278004 531676 278604 531678
rect 386938 531676 387262 531678
rect 422004 531676 422604 531678
rect 516938 531676 517262 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 136982 531654
rect 137218 531418 170186 531654
rect 170422 531418 266982 531654
rect 267218 531418 278186 531654
rect 278422 531418 386982 531654
rect 387218 531418 422186 531654
rect 422422 531418 516982 531654
rect 517218 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 136982 531334
rect 137218 531098 170186 531334
rect 170422 531098 266982 531334
rect 267218 531098 278186 531334
rect 278422 531098 386982 531334
rect 387218 531098 422186 531334
rect 422422 531098 516982 531334
rect 517218 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 136938 531074 137262 531076
rect 170004 531074 170604 531076
rect 266938 531074 267262 531076
rect 278004 531074 278604 531076
rect 386938 531074 387262 531076
rect 422004 531074 422604 531076
rect 516938 531074 517262 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 136938 528076 137262 528078
rect 166404 528076 167004 528078
rect 266938 528076 267262 528078
rect 274404 528076 275004 528078
rect 386938 528076 387262 528078
rect 418404 528076 419004 528078
rect 516938 528076 517262 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 136982 528054
rect 137218 527818 166586 528054
rect 166822 527818 266982 528054
rect 267218 527818 274586 528054
rect 274822 527818 386982 528054
rect 387218 527818 418586 528054
rect 418822 527818 516982 528054
rect 517218 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 136982 527734
rect 137218 527498 166586 527734
rect 166822 527498 266982 527734
rect 267218 527498 274586 527734
rect 274822 527498 386982 527734
rect 387218 527498 418586 527734
rect 418822 527498 516982 527734
rect 517218 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 136938 527474 137262 527476
rect 166404 527474 167004 527476
rect 266938 527474 267262 527476
rect 274404 527474 275004 527476
rect 386938 527474 387262 527476
rect 418404 527474 419004 527476
rect 516938 527474 517262 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 136938 524476 137262 524478
rect 162804 524476 163404 524478
rect 266938 524476 267262 524478
rect 270804 524476 271404 524478
rect 386938 524476 387262 524478
rect 414804 524476 415404 524478
rect 516938 524476 517262 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 136982 524454
rect 137218 524218 162986 524454
rect 163222 524218 266982 524454
rect 267218 524218 270986 524454
rect 271222 524218 386982 524454
rect 387218 524218 414986 524454
rect 415222 524218 516982 524454
rect 517218 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 136982 524134
rect 137218 523898 162986 524134
rect 163222 523898 266982 524134
rect 267218 523898 270986 524134
rect 271222 523898 386982 524134
rect 387218 523898 414986 524134
rect 415222 523898 516982 524134
rect 517218 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 136938 523874 137262 523876
rect 162804 523874 163404 523876
rect 266938 523874 267262 523876
rect 270804 523874 271404 523876
rect 386938 523874 387262 523876
rect 414804 523874 415404 523876
rect 516938 523874 517262 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 136494 517276 136814 517278
rect 155604 517276 156204 517278
rect 266494 517276 266814 517278
rect 299604 517276 300204 517278
rect 386494 517276 386814 517278
rect 407604 517276 408204 517278
rect 516494 517276 516814 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 136536 517254
rect 136772 517018 155786 517254
rect 156022 517018 266536 517254
rect 266772 517018 299786 517254
rect 300022 517018 386536 517254
rect 386772 517018 407786 517254
rect 408022 517018 516536 517254
rect 516772 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 136536 516934
rect 136772 516698 155786 516934
rect 156022 516698 266536 516934
rect 266772 516698 299786 516934
rect 300022 516698 386536 516934
rect 386772 516698 407786 516934
rect 408022 516698 516536 516934
rect 516772 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 136494 516674 136814 516676
rect 155604 516674 156204 516676
rect 266494 516674 266814 516676
rect 299604 516674 300204 516676
rect 386494 516674 386814 516676
rect 407604 516674 408204 516676
rect 516494 516674 516814 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 136494 513676 136814 513678
rect 152004 513676 152604 513678
rect 266494 513676 266814 513678
rect 296004 513676 296604 513678
rect 386494 513676 386814 513678
rect 404004 513676 404604 513678
rect 516494 513676 516814 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 136536 513654
rect 136772 513418 152186 513654
rect 152422 513418 266536 513654
rect 266772 513418 296186 513654
rect 296422 513418 386536 513654
rect 386772 513418 404186 513654
rect 404422 513418 516536 513654
rect 516772 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 136536 513334
rect 136772 513098 152186 513334
rect 152422 513098 266536 513334
rect 266772 513098 296186 513334
rect 296422 513098 386536 513334
rect 386772 513098 404186 513334
rect 404422 513098 516536 513334
rect 516772 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 136494 513074 136814 513076
rect 152004 513074 152604 513076
rect 266494 513074 266814 513076
rect 296004 513074 296604 513076
rect 386494 513074 386814 513076
rect 404004 513074 404604 513076
rect 516494 513074 516814 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 136494 510076 136814 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 266494 510076 266814 510078
rect 292404 510076 293004 510078
rect 386494 510076 386814 510078
rect 400404 510076 401004 510078
rect 516494 510076 516814 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 136536 510054
rect 136772 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 266536 510054
rect 266772 509818 292586 510054
rect 292822 509818 386536 510054
rect 386772 509818 400586 510054
rect 400822 509818 516536 510054
rect 516772 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 136536 509734
rect 136772 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 266536 509734
rect 266772 509498 292586 509734
rect 292822 509498 386536 509734
rect 386772 509498 400586 509734
rect 400822 509498 516536 509734
rect 516772 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 136494 509474 136814 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 266494 509474 266814 509476
rect 292404 509474 293004 509476
rect 386494 509474 386814 509476
rect 400404 509474 401004 509476
rect 516494 509474 516814 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 136494 506476 136814 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 266494 506476 266814 506478
rect 288804 506476 289404 506478
rect 386494 506476 386814 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 516494 506476 516814 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 136536 506454
rect 136772 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 266536 506454
rect 266772 506218 288986 506454
rect 289222 506218 386536 506454
rect 386772 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 516536 506454
rect 516772 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 136536 506134
rect 136772 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 266536 506134
rect 266772 505898 288986 506134
rect 289222 505898 386536 506134
rect 386772 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 516536 506134
rect 516772 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 136494 505874 136814 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 266494 505874 266814 505876
rect 288804 505874 289404 505876
rect 386494 505874 386814 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 516494 505874 516814 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 136938 499276 137262 499278
rect 173604 499276 174204 499278
rect 266938 499276 267262 499278
rect 281604 499276 282204 499278
rect 386938 499276 387262 499278
rect 425604 499276 426204 499278
rect 516938 499276 517262 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 136982 499254
rect 137218 499018 173786 499254
rect 174022 499018 266982 499254
rect 267218 499018 281786 499254
rect 282022 499018 386982 499254
rect 387218 499018 425786 499254
rect 426022 499018 516982 499254
rect 517218 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 136982 498934
rect 137218 498698 173786 498934
rect 174022 498698 266982 498934
rect 267218 498698 281786 498934
rect 282022 498698 386982 498934
rect 387218 498698 425786 498934
rect 426022 498698 516982 498934
rect 517218 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 136938 498674 137262 498676
rect 173604 498674 174204 498676
rect 266938 498674 267262 498676
rect 281604 498674 282204 498676
rect 386938 498674 387262 498676
rect 425604 498674 426204 498676
rect 516938 498674 517262 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 136938 495676 137262 495678
rect 170004 495676 170604 495678
rect 266938 495676 267262 495678
rect 278004 495676 278604 495678
rect 386938 495676 387262 495678
rect 422004 495676 422604 495678
rect 516938 495676 517262 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 136982 495654
rect 137218 495418 170186 495654
rect 170422 495418 266982 495654
rect 267218 495418 278186 495654
rect 278422 495418 386982 495654
rect 387218 495418 422186 495654
rect 422422 495418 516982 495654
rect 517218 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 136982 495334
rect 137218 495098 170186 495334
rect 170422 495098 266982 495334
rect 267218 495098 278186 495334
rect 278422 495098 386982 495334
rect 387218 495098 422186 495334
rect 422422 495098 516982 495334
rect 517218 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 136938 495074 137262 495076
rect 170004 495074 170604 495076
rect 266938 495074 267262 495076
rect 278004 495074 278604 495076
rect 386938 495074 387262 495076
rect 422004 495074 422604 495076
rect 516938 495074 517262 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 136938 492076 137262 492078
rect 166404 492076 167004 492078
rect 266938 492076 267262 492078
rect 274404 492076 275004 492078
rect 386938 492076 387262 492078
rect 418404 492076 419004 492078
rect 516938 492076 517262 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 136982 492054
rect 137218 491818 166586 492054
rect 166822 491818 266982 492054
rect 267218 491818 274586 492054
rect 274822 491818 386982 492054
rect 387218 491818 418586 492054
rect 418822 491818 516982 492054
rect 517218 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 136982 491734
rect 137218 491498 166586 491734
rect 166822 491498 266982 491734
rect 267218 491498 274586 491734
rect 274822 491498 386982 491734
rect 387218 491498 418586 491734
rect 418822 491498 516982 491734
rect 517218 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 136938 491474 137262 491476
rect 166404 491474 167004 491476
rect 266938 491474 267262 491476
rect 274404 491474 275004 491476
rect 386938 491474 387262 491476
rect 418404 491474 419004 491476
rect 516938 491474 517262 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 136938 488476 137262 488478
rect 162804 488476 163404 488478
rect 266938 488476 267262 488478
rect 270804 488476 271404 488478
rect 386938 488476 387262 488478
rect 414804 488476 415404 488478
rect 516938 488476 517262 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 136982 488454
rect 137218 488218 162986 488454
rect 163222 488218 266982 488454
rect 267218 488218 270986 488454
rect 271222 488218 386982 488454
rect 387218 488218 414986 488454
rect 415222 488218 516982 488454
rect 517218 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 136982 488134
rect 137218 487898 162986 488134
rect 163222 487898 266982 488134
rect 267218 487898 270986 488134
rect 271222 487898 386982 488134
rect 387218 487898 414986 488134
rect 415222 487898 516982 488134
rect 517218 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 136938 487874 137262 487876
rect 162804 487874 163404 487876
rect 266938 487874 267262 487876
rect 270804 487874 271404 487876
rect 386938 487874 387262 487876
rect 414804 487874 415404 487876
rect 516938 487874 517262 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 136494 481276 136814 481278
rect 155604 481276 156204 481278
rect 266494 481276 266814 481278
rect 299604 481276 300204 481278
rect 386494 481276 386814 481278
rect 407604 481276 408204 481278
rect 516494 481276 516814 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 136536 481254
rect 136772 481018 155786 481254
rect 156022 481018 266536 481254
rect 266772 481018 299786 481254
rect 300022 481018 386536 481254
rect 386772 481018 407786 481254
rect 408022 481018 516536 481254
rect 516772 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 136536 480934
rect 136772 480698 155786 480934
rect 156022 480698 266536 480934
rect 266772 480698 299786 480934
rect 300022 480698 386536 480934
rect 386772 480698 407786 480934
rect 408022 480698 516536 480934
rect 516772 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 136494 480674 136814 480676
rect 155604 480674 156204 480676
rect 266494 480674 266814 480676
rect 299604 480674 300204 480676
rect 386494 480674 386814 480676
rect 407604 480674 408204 480676
rect 516494 480674 516814 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 136494 477676 136814 477678
rect 152004 477676 152604 477678
rect 266494 477676 266814 477678
rect 296004 477676 296604 477678
rect 386494 477676 386814 477678
rect 404004 477676 404604 477678
rect 516494 477676 516814 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 136536 477654
rect 136772 477418 152186 477654
rect 152422 477418 266536 477654
rect 266772 477418 296186 477654
rect 296422 477418 386536 477654
rect 386772 477418 404186 477654
rect 404422 477418 516536 477654
rect 516772 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 136536 477334
rect 136772 477098 152186 477334
rect 152422 477098 266536 477334
rect 266772 477098 296186 477334
rect 296422 477098 386536 477334
rect 386772 477098 404186 477334
rect 404422 477098 516536 477334
rect 516772 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 136494 477074 136814 477076
rect 152004 477074 152604 477076
rect 266494 477074 266814 477076
rect 296004 477074 296604 477076
rect 386494 477074 386814 477076
rect 404004 477074 404604 477076
rect 516494 477074 516814 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 136494 474076 136814 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 266494 474076 266814 474078
rect 292404 474076 293004 474078
rect 386494 474076 386814 474078
rect 400404 474076 401004 474078
rect 516494 474076 516814 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 136536 474054
rect 136772 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 266536 474054
rect 266772 473818 292586 474054
rect 292822 473818 386536 474054
rect 386772 473818 400586 474054
rect 400822 473818 516536 474054
rect 516772 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 136536 473734
rect 136772 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 266536 473734
rect 266772 473498 292586 473734
rect 292822 473498 386536 473734
rect 386772 473498 400586 473734
rect 400822 473498 516536 473734
rect 516772 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 136494 473474 136814 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 266494 473474 266814 473476
rect 292404 473474 293004 473476
rect 386494 473474 386814 473476
rect 400404 473474 401004 473476
rect 516494 473474 516814 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 136494 470476 136814 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 266494 470476 266814 470478
rect 288804 470476 289404 470478
rect 386494 470476 386814 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 516494 470476 516814 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 136536 470454
rect 136772 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 266536 470454
rect 266772 470218 288986 470454
rect 289222 470218 386536 470454
rect 386772 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 516536 470454
rect 516772 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 136536 470134
rect 136772 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 266536 470134
rect 266772 469898 288986 470134
rect 289222 469898 386536 470134
rect 386772 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 516536 470134
rect 516772 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 136494 469874 136814 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 266494 469874 266814 469876
rect 288804 469874 289404 469876
rect 386494 469874 386814 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 516494 469874 516814 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 136938 463276 137262 463278
rect 173604 463276 174204 463278
rect 266938 463276 267262 463278
rect 281604 463276 282204 463278
rect 386938 463276 387262 463278
rect 425604 463276 426204 463278
rect 516938 463276 517262 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 136982 463254
rect 137218 463018 173786 463254
rect 174022 463018 266982 463254
rect 267218 463018 281786 463254
rect 282022 463018 386982 463254
rect 387218 463018 425786 463254
rect 426022 463018 516982 463254
rect 517218 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 136982 462934
rect 137218 462698 173786 462934
rect 174022 462698 266982 462934
rect 267218 462698 281786 462934
rect 282022 462698 386982 462934
rect 387218 462698 425786 462934
rect 426022 462698 516982 462934
rect 517218 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 136938 462674 137262 462676
rect 173604 462674 174204 462676
rect 266938 462674 267262 462676
rect 281604 462674 282204 462676
rect 386938 462674 387262 462676
rect 425604 462674 426204 462676
rect 516938 462674 517262 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 170004 459676 170604 459678
rect 278004 459676 278604 459678
rect 422004 459676 422604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 170186 459654
rect 170422 459418 278186 459654
rect 278422 459418 422186 459654
rect 422422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 170186 459334
rect 170422 459098 278186 459334
rect 278422 459098 422186 459334
rect 422422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 170004 459074 170604 459076
rect 278004 459074 278604 459076
rect 422004 459074 422604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 64208 434476 64528 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 64250 434454
rect 64486 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 64250 434134
rect 64486 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 64208 433874 64528 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 79568 427276 79888 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 79610 427254
rect 79846 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 79610 426934
rect 79846 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 79568 426674 79888 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 79568 423676 79888 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 79610 423654
rect 79846 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 79610 423334
rect 79846 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 79568 423074 79888 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 79568 420076 79888 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 79610 420054
rect 79846 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 79610 419734
rect 79846 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 79568 419474 79888 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 79568 416476 79888 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 79610 416454
rect 79846 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 79610 416134
rect 79846 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 79568 415874 79888 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 64208 409276 64528 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 64250 409254
rect 64486 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 64250 408934
rect 64486 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 64208 408674 64528 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 64208 405676 64528 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 64250 405654
rect 64486 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 64250 405334
rect 64486 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 64208 405074 64528 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 64208 402076 64528 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 64250 402054
rect 64486 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 64250 401734
rect 64486 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 64208 401474 64528 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 64208 398476 64528 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 64250 398454
rect 64486 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 64250 398134
rect 64486 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 64208 397874 64528 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 79568 391276 79888 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 79610 391254
rect 79846 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 79610 390934
rect 79846 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 79568 390674 79888 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 79568 387676 79888 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 79610 387654
rect 79846 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 79610 387334
rect 79846 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 79568 387074 79888 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 79568 384076 79888 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 79610 384054
rect 79846 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 79610 383734
rect 79846 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 79568 383474 79888 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 79568 380476 79888 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 79610 380454
rect 79846 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 79610 380134
rect 79846 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 79568 379874 79888 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 64208 373276 64528 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 64250 373254
rect 64486 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 64250 372934
rect 64486 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 64208 372674 64528 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 64208 369676 64528 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 64250 369654
rect 64486 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 64250 369334
rect 64486 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 64208 369074 64528 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 64208 366076 64528 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 64250 366054
rect 64486 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 64250 365734
rect 64486 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 64208 365474 64528 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 64208 362476 64528 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 64250 362454
rect 64486 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 64250 362134
rect 64486 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 64208 361874 64528 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 79568 355276 79888 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 79610 355254
rect 79846 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 79610 354934
rect 79846 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 79568 354674 79888 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 79568 351676 79888 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 79610 351654
rect 79846 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 79610 351334
rect 79846 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 79568 351074 79888 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 79568 348076 79888 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 79610 348054
rect 79846 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 79610 347734
rect 79846 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 79568 347474 79888 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 79568 344476 79888 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 79610 344454
rect 79846 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 79610 344134
rect 79846 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 79568 343874 79888 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 64208 337276 64528 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 64250 337254
rect 64486 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 64250 336934
rect 64486 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 64208 336674 64528 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 64208 333676 64528 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 64250 333654
rect 64486 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 64250 333334
rect 64486 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 64208 333074 64528 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 64208 330076 64528 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 64250 330054
rect 64486 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 64250 329734
rect 64486 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 64208 329474 64528 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 64208 326476 64528 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 64250 326454
rect 64486 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 64250 326134
rect 64486 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 64208 325874 64528 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 79568 319276 79888 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 79610 319254
rect 79846 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 79610 318934
rect 79846 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 79568 318674 79888 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 79568 315676 79888 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 79610 315654
rect 79846 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 79610 315334
rect 79846 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 79568 315074 79888 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 79568 312076 79888 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 79610 312054
rect 79846 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 79610 311734
rect 79846 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 79568 311474 79888 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 79568 308476 79888 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 79610 308454
rect 79846 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 79610 308134
rect 79846 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 79568 307874 79888 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 64208 301276 64528 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 64250 301254
rect 64486 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 64250 300934
rect 64486 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 64208 300674 64528 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 64208 297676 64528 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 64250 297654
rect 64486 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 64250 297334
rect 64486 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 64208 297074 64528 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 64208 294076 64528 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 64250 294054
rect 64486 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 64250 293734
rect 64486 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 64208 293474 64528 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 64208 290476 64528 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 64250 290454
rect 64486 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 64250 290134
rect 64486 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 64208 289874 64528 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 79568 283276 79888 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 79610 283254
rect 79846 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 79610 282934
rect 79846 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 79568 282674 79888 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 79568 279676 79888 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 79610 279654
rect 79846 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 79610 279334
rect 79846 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 79568 279074 79888 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 79568 276076 79888 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 79610 276054
rect 79846 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 79610 275734
rect 79846 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 79568 275474 79888 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 79568 272476 79888 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 79610 272454
rect 79846 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 79610 272134
rect 79846 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 79568 271874 79888 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 64208 265276 64528 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 64250 265254
rect 64486 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 64250 264934
rect 64486 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 64208 264674 64528 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 64208 261676 64528 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 64250 261654
rect 64486 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 64250 261334
rect 64486 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 64208 261074 64528 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 64208 258076 64528 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 64250 258054
rect 64486 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 64250 257734
rect 64486 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 64208 257474 64528 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 64208 254476 64528 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 64250 254454
rect 64486 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 64250 254134
rect 64486 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 64208 253874 64528 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 79568 247276 79888 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 79610 247254
rect 79846 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 79610 246934
rect 79846 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 79568 246674 79888 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 79568 243676 79888 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 79610 243654
rect 79846 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 79610 243334
rect 79846 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 79568 243074 79888 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 79568 240076 79888 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 79610 240054
rect 79846 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 79610 239734
rect 79846 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 79568 239474 79888 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 79568 236476 79888 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 79610 236454
rect 79846 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 79610 236134
rect 79846 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 79568 235874 79888 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 64208 229276 64528 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 64250 229254
rect 64486 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 64250 228934
rect 64486 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 64208 228674 64528 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 64208 225676 64528 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 64250 225654
rect 64486 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 64250 225334
rect 64486 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 64208 225074 64528 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 64208 222076 64528 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 64250 222054
rect 64486 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 64250 221734
rect 64486 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 64208 221474 64528 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 64208 218476 64528 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 64250 218454
rect 64486 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 64250 218134
rect 64486 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 64208 217874 64528 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 79568 211276 79888 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 79610 211254
rect 79846 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 79610 210934
rect 79846 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 79568 210674 79888 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 79568 207676 79888 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 79610 207654
rect 79846 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 79610 207334
rect 79846 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 79568 207074 79888 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 79568 204076 79888 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 79610 204054
rect 79846 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 79610 203734
rect 79846 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 79568 203474 79888 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use sram_1rw1r_32_256_8_sky130  sram3
timestamp 1608756459
transform 1 0 440000 0 1 460000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram2
timestamp 1608756459
transform 1 0 310000 0 1 460000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram1
timestamp 1608756459
transform 1 0 190000 0 1 460000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram0
timestamp 1608756459
transform 1 0 60000 0 1 460000
box 0 0 77296 91247
use hs32_core1  core1
timestamp 1608756459
transform 1 0 60000 0 1 200000
box 0 0 240000 240000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
