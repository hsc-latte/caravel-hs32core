VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2611.950 1200.780 2612.270 1200.840 ;
        RECT 2625.290 1200.780 2625.610 1200.840 ;
        RECT 2611.950 1200.640 2625.610 1200.780 ;
        RECT 2611.950 1200.580 2612.270 1200.640 ;
        RECT 2625.290 1200.580 2625.610 1200.640 ;
        RECT 2625.290 89.660 2625.610 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2625.290 89.520 2899.310 89.660 ;
        RECT 2625.290 89.460 2625.610 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2611.980 1200.580 2612.240 1200.840 ;
        RECT 2625.320 1200.580 2625.580 1200.840 ;
        RECT 2625.320 89.460 2625.580 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2611.970 1202.395 2612.250 1202.765 ;
        RECT 2612.040 1200.870 2612.180 1202.395 ;
        RECT 2611.980 1200.550 2612.240 1200.870 ;
        RECT 2625.320 1200.550 2625.580 1200.870 ;
        RECT 2625.380 89.750 2625.520 1200.550 ;
        RECT 2625.320 89.430 2625.580 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2611.970 1202.440 2612.250 1202.720 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2596.000 1204.800 2600.000 1205.400 ;
        RECT 2599.310 1202.730 2599.610 1204.800 ;
        RECT 2611.945 1202.730 2612.275 1202.745 ;
        RECT 2599.310 1202.430 2612.275 1202.730 ;
        RECT 2611.945 1202.415 2612.275 1202.430 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.310 2429.200 2619.630 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 2619.310 2429.060 2901.150 2429.200 ;
        RECT 2619.310 2429.000 2619.630 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 2608.270 1521.400 2608.590 1521.460 ;
        RECT 2619.310 1521.400 2619.630 1521.460 ;
        RECT 2608.270 1521.260 2619.630 1521.400 ;
        RECT 2608.270 1521.200 2608.590 1521.260 ;
        RECT 2619.310 1521.200 2619.630 1521.260 ;
      LAYER via ;
        RECT 2619.340 2429.000 2619.600 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 2608.300 1521.200 2608.560 1521.460 ;
        RECT 2619.340 1521.200 2619.600 1521.460 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 2619.340 2428.970 2619.600 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 2619.400 1521.490 2619.540 2428.970 ;
        RECT 2608.300 1521.170 2608.560 1521.490 ;
        RECT 2619.340 1521.170 2619.600 1521.490 ;
        RECT 2608.360 1521.005 2608.500 1521.170 ;
        RECT 2608.290 1520.635 2608.570 1521.005 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 2608.290 1520.680 2608.570 1520.960 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2608.265 1520.970 2608.595 1520.985 ;
        RECT 2599.460 1520.920 2608.595 1520.970 ;
        RECT 2596.000 1520.670 2608.595 1520.920 ;
        RECT 2596.000 1520.320 2600.000 1520.670 ;
        RECT 2608.265 1520.655 2608.595 1520.670 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.850 2663.800 2619.170 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 2618.850 2663.660 2901.150 2663.800 ;
        RECT 2618.850 2663.600 2619.170 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 2608.270 1552.340 2608.590 1552.400 ;
        RECT 2618.850 1552.340 2619.170 1552.400 ;
        RECT 2608.270 1552.200 2619.170 1552.340 ;
        RECT 2608.270 1552.140 2608.590 1552.200 ;
        RECT 2618.850 1552.140 2619.170 1552.200 ;
      LAYER via ;
        RECT 2618.880 2663.600 2619.140 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 2608.300 1552.140 2608.560 1552.400 ;
        RECT 2618.880 1552.140 2619.140 1552.400 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 2618.880 2663.570 2619.140 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 2618.940 1552.430 2619.080 2663.570 ;
        RECT 2608.300 1552.285 2608.560 1552.430 ;
        RECT 2608.290 1551.915 2608.570 1552.285 ;
        RECT 2618.880 1552.110 2619.140 1552.430 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
        RECT 2608.290 1551.960 2608.570 1552.240 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2608.265 1552.250 2608.595 1552.265 ;
        RECT 2599.460 1552.200 2608.595 1552.250 ;
        RECT 2596.000 1551.950 2608.595 1552.200 ;
        RECT 2596.000 1551.600 2600.000 1551.950 ;
        RECT 2608.265 1551.935 2608.595 1551.950 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 2898.400 2618.710 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2618.390 2898.260 2901.150 2898.400 ;
        RECT 2618.390 2898.200 2618.710 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2608.270 1584.300 2608.590 1584.360 ;
        RECT 2618.390 1584.300 2618.710 1584.360 ;
        RECT 2608.270 1584.160 2618.710 1584.300 ;
        RECT 2608.270 1584.100 2608.590 1584.160 ;
        RECT 2618.390 1584.100 2618.710 1584.160 ;
      LAYER via ;
        RECT 2618.420 2898.200 2618.680 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2608.300 1584.100 2608.560 1584.360 ;
        RECT 2618.420 1584.100 2618.680 1584.360 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2618.420 2898.170 2618.680 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2618.480 1584.390 2618.620 2898.170 ;
        RECT 2608.300 1584.245 2608.560 1584.390 ;
        RECT 2608.290 1583.875 2608.570 1584.245 ;
        RECT 2618.420 1584.070 2618.680 1584.390 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 2608.290 1583.920 2608.570 1584.200 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2608.265 1584.210 2608.595 1584.225 ;
        RECT 2599.460 1584.160 2608.595 1584.210 ;
        RECT 2596.000 1583.910 2608.595 1584.160 ;
        RECT 2596.000 1583.560 2600.000 1583.910 ;
        RECT 2608.265 1583.895 2608.595 1583.910 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2625.290 3133.000 2625.610 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2625.290 3132.860 2901.150 3133.000 ;
        RECT 2625.290 3132.800 2625.610 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 2612.870 1617.280 2613.190 1617.340 ;
        RECT 2625.290 1617.280 2625.610 1617.340 ;
        RECT 2612.870 1617.140 2625.610 1617.280 ;
        RECT 2612.870 1617.080 2613.190 1617.140 ;
        RECT 2625.290 1617.080 2625.610 1617.140 ;
      LAYER via ;
        RECT 2625.320 3132.800 2625.580 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 2612.900 1617.080 2613.160 1617.340 ;
        RECT 2625.320 1617.080 2625.580 1617.340 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2625.320 3132.770 2625.580 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 2625.380 1617.370 2625.520 3132.770 ;
        RECT 2612.900 1617.050 2613.160 1617.370 ;
        RECT 2625.320 1617.050 2625.580 1617.370 ;
        RECT 2612.960 1615.525 2613.100 1617.050 ;
        RECT 2612.890 1615.155 2613.170 1615.525 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 2612.890 1615.200 2613.170 1615.480 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2612.865 1615.490 2613.195 1615.505 ;
        RECT 2599.460 1615.440 2613.195 1615.490 ;
        RECT 2596.000 1615.190 2613.195 1615.440 ;
        RECT 2596.000 1614.840 2600.000 1615.190 ;
        RECT 2612.865 1615.175 2613.195 1615.190 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2645.990 3367.600 2646.310 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2645.990 3367.460 2901.150 3367.600 ;
        RECT 2645.990 3367.400 2646.310 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 2613.790 1642.780 2614.110 1642.840 ;
        RECT 2645.990 1642.780 2646.310 1642.840 ;
        RECT 2613.790 1642.640 2646.310 1642.780 ;
        RECT 2613.790 1642.580 2614.110 1642.640 ;
        RECT 2645.990 1642.580 2646.310 1642.640 ;
      LAYER via ;
        RECT 2646.020 3367.400 2646.280 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 2613.820 1642.580 2614.080 1642.840 ;
        RECT 2646.020 1642.580 2646.280 1642.840 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2646.020 3367.370 2646.280 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 2613.810 1647.115 2614.090 1647.485 ;
        RECT 2613.880 1642.870 2614.020 1647.115 ;
        RECT 2646.080 1642.870 2646.220 3367.370 ;
        RECT 2613.820 1642.550 2614.080 1642.870 ;
        RECT 2646.020 1642.550 2646.280 1642.870 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 2613.810 1647.160 2614.090 1647.440 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2613.785 1647.450 2614.115 1647.465 ;
        RECT 2599.460 1647.400 2614.115 1647.450 ;
        RECT 2596.000 1647.150 2614.115 1647.400 ;
        RECT 2596.000 1646.800 2600.000 1647.150 ;
        RECT 2613.785 1647.135 2614.115 1647.150 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2659.790 3501.560 2660.110 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 2659.790 3501.420 2798.570 3501.560 ;
        RECT 2659.790 3501.360 2660.110 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
        RECT 2614.250 1683.580 2614.570 1683.640 ;
        RECT 2659.790 1683.580 2660.110 1683.640 ;
        RECT 2614.250 1683.440 2660.110 1683.580 ;
        RECT 2614.250 1683.380 2614.570 1683.440 ;
        RECT 2659.790 1683.380 2660.110 1683.440 ;
      LAYER via ;
        RECT 2659.820 3501.360 2660.080 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
        RECT 2614.280 1683.380 2614.540 1683.640 ;
        RECT 2659.820 1683.380 2660.080 1683.640 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 2659.820 3501.330 2660.080 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 2659.880 1683.670 2660.020 3501.330 ;
        RECT 2614.280 1683.350 2614.540 1683.670 ;
        RECT 2659.820 1683.350 2660.080 1683.670 ;
        RECT 2614.340 1678.765 2614.480 1683.350 ;
        RECT 2614.270 1678.395 2614.550 1678.765 ;
      LAYER via2 ;
        RECT 2614.270 1678.440 2614.550 1678.720 ;
      LAYER met3 ;
        RECT 2614.245 1678.730 2614.575 1678.745 ;
        RECT 2599.460 1678.680 2614.575 1678.730 ;
        RECT 2596.000 1678.430 2614.575 1678.680 ;
        RECT 2596.000 1678.080 2600.000 1678.430 ;
        RECT 2614.245 1678.415 2614.575 1678.430 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2473.950 3498.500 2474.270 3498.560 ;
        RECT 2476.710 3498.500 2477.030 3498.560 ;
        RECT 2473.950 3498.360 2477.030 3498.500 ;
        RECT 2473.950 3498.300 2474.270 3498.360 ;
        RECT 2476.710 3498.300 2477.030 3498.360 ;
        RECT 2476.710 3054.120 2477.030 3054.180 ;
        RECT 2602.750 3054.120 2603.070 3054.180 ;
        RECT 2476.710 3053.980 2603.070 3054.120 ;
        RECT 2476.710 3053.920 2477.030 3053.980 ;
        RECT 2602.750 3053.920 2603.070 3053.980 ;
      LAYER via ;
        RECT 2473.980 3498.300 2474.240 3498.560 ;
        RECT 2476.740 3498.300 2477.000 3498.560 ;
        RECT 2476.740 3053.920 2477.000 3054.180 ;
        RECT 2602.780 3053.920 2603.040 3054.180 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3498.590 2474.180 3517.600 ;
        RECT 2473.980 3498.270 2474.240 3498.590 ;
        RECT 2476.740 3498.270 2477.000 3498.590 ;
        RECT 2476.800 3054.210 2476.940 3498.270 ;
        RECT 2476.740 3053.890 2477.000 3054.210 ;
        RECT 2602.780 3053.890 2603.040 3054.210 ;
        RECT 2602.840 1710.725 2602.980 3053.890 ;
        RECT 2602.770 1710.355 2603.050 1710.725 ;
      LAYER via2 ;
        RECT 2602.770 1710.400 2603.050 1710.680 ;
      LAYER met3 ;
        RECT 2602.745 1710.690 2603.075 1710.705 ;
        RECT 2599.460 1710.640 2603.075 1710.690 ;
        RECT 2596.000 1710.390 2603.075 1710.640 ;
        RECT 2596.000 1710.040 2600.000 1710.390 ;
        RECT 2602.745 1710.375 2603.075 1710.390 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2149.190 3498.500 2149.510 3498.560 ;
        RECT 2152.410 3498.500 2152.730 3498.560 ;
        RECT 2149.190 3498.360 2152.730 3498.500 ;
        RECT 2149.190 3498.300 2149.510 3498.360 ;
        RECT 2152.410 3498.300 2152.730 3498.360 ;
        RECT 2152.410 3053.440 2152.730 3053.500 ;
        RECT 2603.210 3053.440 2603.530 3053.500 ;
        RECT 2152.410 3053.300 2603.530 3053.440 ;
        RECT 2152.410 3053.240 2152.730 3053.300 ;
        RECT 2603.210 3053.240 2603.530 3053.300 ;
      LAYER via ;
        RECT 2149.220 3498.300 2149.480 3498.560 ;
        RECT 2152.440 3498.300 2152.700 3498.560 ;
        RECT 2152.440 3053.240 2152.700 3053.500 ;
        RECT 2603.240 3053.240 2603.500 3053.500 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3498.590 2149.420 3517.600 ;
        RECT 2149.220 3498.270 2149.480 3498.590 ;
        RECT 2152.440 3498.270 2152.700 3498.590 ;
        RECT 2152.500 3053.530 2152.640 3498.270 ;
        RECT 2152.440 3053.210 2152.700 3053.530 ;
        RECT 2603.240 3053.210 2603.500 3053.530 ;
        RECT 2603.300 1742.005 2603.440 3053.210 ;
        RECT 2603.230 1741.635 2603.510 1742.005 ;
      LAYER via2 ;
        RECT 2603.230 1741.680 2603.510 1741.960 ;
      LAYER met3 ;
        RECT 2603.205 1741.970 2603.535 1741.985 ;
        RECT 2599.460 1741.920 2603.535 1741.970 ;
        RECT 2596.000 1741.670 2603.535 1741.920 ;
        RECT 2596.000 1741.320 2600.000 1741.670 ;
        RECT 2603.205 1741.655 2603.535 1741.670 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3498.500 1825.210 3498.560 ;
        RECT 1828.110 3498.500 1828.430 3498.560 ;
        RECT 1824.890 3498.360 1828.430 3498.500 ;
        RECT 1824.890 3498.300 1825.210 3498.360 ;
        RECT 1828.110 3498.300 1828.430 3498.360 ;
        RECT 1828.110 3053.100 1828.430 3053.160 ;
        RECT 2603.670 3053.100 2603.990 3053.160 ;
        RECT 1828.110 3052.960 2603.990 3053.100 ;
        RECT 1828.110 3052.900 1828.430 3052.960 ;
        RECT 2603.670 3052.900 2603.990 3052.960 ;
      LAYER via ;
        RECT 1824.920 3498.300 1825.180 3498.560 ;
        RECT 1828.140 3498.300 1828.400 3498.560 ;
        RECT 1828.140 3052.900 1828.400 3053.160 ;
        RECT 2603.700 3052.900 2603.960 3053.160 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3498.590 1825.120 3517.600 ;
        RECT 1824.920 3498.270 1825.180 3498.590 ;
        RECT 1828.140 3498.270 1828.400 3498.590 ;
        RECT 1828.200 3053.190 1828.340 3498.270 ;
        RECT 1828.140 3052.870 1828.400 3053.190 ;
        RECT 2603.700 3052.870 2603.960 3053.190 ;
        RECT 2603.760 1773.965 2603.900 3052.870 ;
        RECT 2603.690 1773.595 2603.970 1773.965 ;
      LAYER via2 ;
        RECT 2603.690 1773.640 2603.970 1773.920 ;
      LAYER met3 ;
        RECT 2603.665 1773.930 2603.995 1773.945 ;
        RECT 2599.460 1773.880 2603.995 1773.930 ;
        RECT 2596.000 1773.630 2603.995 1773.880 ;
        RECT 2596.000 1773.280 2600.000 1773.630 ;
        RECT 2603.665 1773.615 2603.995 1773.630 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1502.890 3498.500 1503.210 3498.560 ;
        RECT 1500.590 3498.360 1503.210 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1502.890 3498.300 1503.210 3498.360 ;
        RECT 1502.890 2399.620 1503.210 2399.680 ;
        RECT 2605.050 2399.620 2605.370 2399.680 ;
        RECT 1502.890 2399.480 2605.370 2399.620 ;
        RECT 1502.890 2399.420 1503.210 2399.480 ;
        RECT 2605.050 2399.420 2605.370 2399.480 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1502.920 3498.300 1503.180 3498.560 ;
        RECT 1502.920 2399.420 1503.180 2399.680 ;
        RECT 2605.080 2399.420 2605.340 2399.680 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1502.920 3498.270 1503.180 3498.590 ;
        RECT 1502.980 2399.710 1503.120 3498.270 ;
        RECT 1502.920 2399.390 1503.180 2399.710 ;
        RECT 2605.080 2399.390 2605.340 2399.710 ;
        RECT 2605.140 1805.245 2605.280 2399.390 ;
        RECT 2605.070 1804.875 2605.350 1805.245 ;
      LAYER via2 ;
        RECT 2605.070 1804.920 2605.350 1805.200 ;
      LAYER met3 ;
        RECT 2605.045 1805.210 2605.375 1805.225 ;
        RECT 2599.460 1805.160 2605.375 1805.210 ;
        RECT 2596.000 1804.910 2605.375 1805.160 ;
        RECT 2596.000 1804.560 2600.000 1804.910 ;
        RECT 2605.045 1804.895 2605.375 1804.910 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2608.270 1235.460 2608.590 1235.520 ;
        RECT 2639.090 1235.460 2639.410 1235.520 ;
        RECT 2608.270 1235.320 2639.410 1235.460 ;
        RECT 2608.270 1235.260 2608.590 1235.320 ;
        RECT 2639.090 1235.260 2639.410 1235.320 ;
        RECT 2639.090 324.260 2639.410 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2639.090 324.120 2899.310 324.260 ;
        RECT 2639.090 324.060 2639.410 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2608.300 1235.260 2608.560 1235.520 ;
        RECT 2639.120 1235.260 2639.380 1235.520 ;
        RECT 2639.120 324.060 2639.380 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2608.290 1236.395 2608.570 1236.765 ;
        RECT 2608.360 1235.550 2608.500 1236.395 ;
        RECT 2608.300 1235.230 2608.560 1235.550 ;
        RECT 2639.120 1235.230 2639.380 1235.550 ;
        RECT 2639.180 324.350 2639.320 1235.230 ;
        RECT 2639.120 324.030 2639.380 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2608.290 1236.440 2608.570 1236.720 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2608.265 1236.730 2608.595 1236.745 ;
        RECT 2599.460 1236.680 2608.595 1236.730 ;
        RECT 2596.000 1236.430 2608.595 1236.680 ;
        RECT 2596.000 1236.080 2600.000 1236.430 ;
        RECT 2608.265 1236.415 2608.595 1236.430 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1179.510 2399.280 1179.830 2399.340 ;
        RECT 2605.510 2399.280 2605.830 2399.340 ;
        RECT 1179.510 2399.140 2605.830 2399.280 ;
        RECT 1179.510 2399.080 1179.830 2399.140 ;
        RECT 2605.510 2399.080 2605.830 2399.140 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1179.540 2399.080 1179.800 2399.340 ;
        RECT 2605.540 2399.080 2605.800 2399.340 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 2399.370 1179.740 3498.270 ;
        RECT 1179.540 2399.050 1179.800 2399.370 ;
        RECT 2605.540 2399.050 2605.800 2399.370 ;
        RECT 2605.600 1836.525 2605.740 2399.050 ;
        RECT 2605.530 1836.155 2605.810 1836.525 ;
      LAYER via2 ;
        RECT 2605.530 1836.200 2605.810 1836.480 ;
      LAYER met3 ;
        RECT 2605.505 1836.490 2605.835 1836.505 ;
        RECT 2599.460 1836.440 2605.835 1836.490 ;
        RECT 2596.000 1836.190 2605.835 1836.440 ;
        RECT 2596.000 1835.840 2600.000 1836.190 ;
        RECT 2605.505 1836.175 2605.835 1836.190 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3504.620 851.850 3504.680 ;
        RECT 855.210 3504.620 855.530 3504.680 ;
        RECT 851.530 3504.480 855.530 3504.620 ;
        RECT 851.530 3504.420 851.850 3504.480 ;
        RECT 855.210 3504.420 855.530 3504.480 ;
        RECT 855.210 2398.940 855.530 2399.000 ;
        RECT 2605.970 2398.940 2606.290 2399.000 ;
        RECT 855.210 2398.800 2606.290 2398.940 ;
        RECT 855.210 2398.740 855.530 2398.800 ;
        RECT 2605.970 2398.740 2606.290 2398.800 ;
      LAYER via ;
        RECT 851.560 3504.420 851.820 3504.680 ;
        RECT 855.240 3504.420 855.500 3504.680 ;
        RECT 855.240 2398.740 855.500 2399.000 ;
        RECT 2606.000 2398.740 2606.260 2399.000 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3504.710 851.760 3517.600 ;
        RECT 851.560 3504.390 851.820 3504.710 ;
        RECT 855.240 3504.390 855.500 3504.710 ;
        RECT 855.300 2399.030 855.440 3504.390 ;
        RECT 855.240 2398.710 855.500 2399.030 ;
        RECT 2606.000 2398.710 2606.260 2399.030 ;
        RECT 2606.060 1868.485 2606.200 2398.710 ;
        RECT 2605.990 1868.115 2606.270 1868.485 ;
      LAYER via2 ;
        RECT 2605.990 1868.160 2606.270 1868.440 ;
      LAYER met3 ;
        RECT 2605.965 1868.450 2606.295 1868.465 ;
        RECT 2599.460 1868.400 2606.295 1868.450 ;
        RECT 2596.000 1868.150 2606.295 1868.400 ;
        RECT 2596.000 1867.800 2600.000 1868.150 ;
        RECT 2605.965 1868.135 2606.295 1868.150 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 2125.730 2399.960 2126.050 2400.020 ;
        RECT 2172.190 2399.960 2172.510 2400.020 ;
        RECT 2125.730 2399.820 2172.510 2399.960 ;
        RECT 2125.730 2399.760 2126.050 2399.820 ;
        RECT 2172.190 2399.760 2172.510 2399.820 ;
        RECT 2363.550 2399.960 2363.870 2400.020 ;
        RECT 2414.610 2399.960 2414.930 2400.020 ;
        RECT 2363.550 2399.820 2414.930 2399.960 ;
        RECT 2363.550 2399.760 2363.870 2399.820 ;
        RECT 2414.610 2399.760 2414.930 2399.820 ;
        RECT 1220.910 2399.620 1221.230 2399.680 ;
        RECT 1255.410 2399.620 1255.730 2399.680 ;
        RECT 1220.910 2399.480 1255.730 2399.620 ;
        RECT 1220.910 2399.420 1221.230 2399.480 ;
        RECT 1255.410 2399.420 1255.730 2399.480 ;
        RECT 1317.510 2399.620 1317.830 2399.680 ;
        RECT 1352.010 2399.620 1352.330 2399.680 ;
        RECT 1317.510 2399.480 1352.330 2399.620 ;
        RECT 1317.510 2399.420 1317.830 2399.480 ;
        RECT 1352.010 2399.420 1352.330 2399.480 ;
        RECT 834.510 2399.280 834.830 2399.340 ;
        RECT 869.010 2399.280 869.330 2399.340 ;
        RECT 834.510 2399.140 869.330 2399.280 ;
        RECT 834.510 2399.080 834.830 2399.140 ;
        RECT 869.010 2399.080 869.330 2399.140 ;
        RECT 931.110 2399.280 931.430 2399.340 ;
        RECT 965.610 2399.280 965.930 2399.340 ;
        RECT 931.110 2399.140 965.930 2399.280 ;
        RECT 931.110 2399.080 931.430 2399.140 ;
        RECT 965.610 2399.080 965.930 2399.140 ;
        RECT 1027.710 2399.280 1028.030 2399.340 ;
        RECT 1062.210 2399.280 1062.530 2399.340 ;
        RECT 1027.710 2399.140 1062.530 2399.280 ;
        RECT 1027.710 2399.080 1028.030 2399.140 ;
        RECT 1062.210 2399.080 1062.530 2399.140 ;
        RECT 1124.310 2399.280 1124.630 2399.340 ;
        RECT 1158.810 2399.280 1159.130 2399.340 ;
        RECT 1124.310 2399.140 1159.130 2399.280 ;
        RECT 1124.310 2399.080 1124.630 2399.140 ;
        RECT 1158.810 2399.080 1159.130 2399.140 ;
        RECT 732.850 2398.940 733.170 2399.000 ;
        RECT 772.410 2398.940 772.730 2399.000 ;
        RECT 732.850 2398.800 772.730 2398.940 ;
        RECT 732.850 2398.740 733.170 2398.800 ;
        RECT 772.410 2398.740 772.730 2398.800 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 2125.760 2399.760 2126.020 2400.020 ;
        RECT 2172.220 2399.760 2172.480 2400.020 ;
        RECT 2363.580 2399.760 2363.840 2400.020 ;
        RECT 2414.640 2399.760 2414.900 2400.020 ;
        RECT 1220.940 2399.420 1221.200 2399.680 ;
        RECT 1255.440 2399.420 1255.700 2399.680 ;
        RECT 1317.540 2399.420 1317.800 2399.680 ;
        RECT 1352.040 2399.420 1352.300 2399.680 ;
        RECT 834.540 2399.080 834.800 2399.340 ;
        RECT 869.040 2399.080 869.300 2399.340 ;
        RECT 931.140 2399.080 931.400 2399.340 ;
        RECT 965.640 2399.080 965.900 2399.340 ;
        RECT 1027.740 2399.080 1028.000 2399.340 ;
        RECT 1062.240 2399.080 1062.500 2399.340 ;
        RECT 1124.340 2399.080 1124.600 2399.340 ;
        RECT 1158.840 2399.080 1159.100 2399.340 ;
        RECT 732.880 2398.740 733.140 2399.000 ;
        RECT 772.440 2398.740 772.700 2399.000 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 2398.205 531.140 3498.270 ;
        RECT 2124.830 2401.235 2125.110 2401.605 ;
        RECT 1738.430 2399.875 1738.710 2400.245 ;
        RECT 1220.940 2399.390 1221.200 2399.710 ;
        RECT 1255.440 2399.390 1255.700 2399.710 ;
        RECT 1317.540 2399.390 1317.800 2399.710 ;
        RECT 1352.040 2399.390 1352.300 2399.710 ;
        RECT 834.540 2399.050 834.800 2399.370 ;
        RECT 869.040 2399.050 869.300 2399.370 ;
        RECT 931.140 2399.050 931.400 2399.370 ;
        RECT 965.640 2399.050 965.900 2399.370 ;
        RECT 1027.740 2399.050 1028.000 2399.370 ;
        RECT 1062.240 2399.050 1062.500 2399.370 ;
        RECT 1124.340 2399.050 1124.600 2399.370 ;
        RECT 1158.840 2399.050 1159.100 2399.370 ;
        RECT 732.880 2398.885 733.140 2399.030 ;
        RECT 732.870 2398.515 733.150 2398.885 ;
        RECT 772.440 2398.710 772.700 2399.030 ;
        RECT 834.600 2398.885 834.740 2399.050 ;
        RECT 772.500 2398.205 772.640 2398.710 ;
        RECT 834.530 2398.515 834.810 2398.885 ;
        RECT 869.100 2398.205 869.240 2399.050 ;
        RECT 931.200 2398.885 931.340 2399.050 ;
        RECT 931.130 2398.515 931.410 2398.885 ;
        RECT 965.700 2398.205 965.840 2399.050 ;
        RECT 1027.800 2398.885 1027.940 2399.050 ;
        RECT 1027.730 2398.515 1028.010 2398.885 ;
        RECT 1062.300 2398.205 1062.440 2399.050 ;
        RECT 1124.400 2398.885 1124.540 2399.050 ;
        RECT 1124.330 2398.515 1124.610 2398.885 ;
        RECT 1158.900 2398.205 1159.040 2399.050 ;
        RECT 1221.000 2398.885 1221.140 2399.390 ;
        RECT 1220.930 2398.515 1221.210 2398.885 ;
        RECT 1255.500 2398.205 1255.640 2399.390 ;
        RECT 1317.600 2398.885 1317.740 2399.390 ;
        RECT 1317.530 2398.515 1317.810 2398.885 ;
        RECT 1352.100 2398.205 1352.240 2399.390 ;
        RECT 1738.500 2398.205 1738.640 2399.875 ;
        RECT 2124.900 2398.885 2125.040 2401.235 ;
        RECT 2125.760 2399.730 2126.020 2400.050 ;
        RECT 2172.220 2399.730 2172.480 2400.050 ;
        RECT 2363.580 2399.730 2363.840 2400.050 ;
        RECT 2414.640 2399.730 2414.900 2400.050 ;
        RECT 2125.820 2398.885 2125.960 2399.730 ;
        RECT 2124.830 2398.515 2125.110 2398.885 ;
        RECT 2125.750 2398.515 2126.030 2398.885 ;
        RECT 530.930 2397.835 531.210 2398.205 ;
        RECT 772.430 2397.835 772.710 2398.205 ;
        RECT 869.030 2397.835 869.310 2398.205 ;
        RECT 965.630 2397.835 965.910 2398.205 ;
        RECT 1062.230 2397.835 1062.510 2398.205 ;
        RECT 1158.830 2397.835 1159.110 2398.205 ;
        RECT 1255.430 2397.835 1255.710 2398.205 ;
        RECT 1352.030 2397.835 1352.310 2398.205 ;
        RECT 1738.430 2397.835 1738.710 2398.205 ;
        RECT 2172.280 2398.090 2172.420 2399.730 ;
        RECT 2269.270 2399.195 2269.550 2399.565 ;
        RECT 2269.340 2398.885 2269.480 2399.195 ;
        RECT 2269.270 2398.515 2269.550 2398.885 ;
        RECT 2172.670 2398.090 2172.950 2398.205 ;
        RECT 2172.280 2397.950 2172.950 2398.090 ;
        RECT 2172.670 2397.835 2172.950 2397.950 ;
        RECT 2363.640 2396.845 2363.780 2399.730 ;
        RECT 2414.700 2399.565 2414.840 2399.730 ;
        RECT 2414.630 2399.195 2414.910 2399.565 ;
        RECT 2363.570 2396.475 2363.850 2396.845 ;
      LAYER via2 ;
        RECT 2124.830 2401.280 2125.110 2401.560 ;
        RECT 1738.430 2399.920 1738.710 2400.200 ;
        RECT 732.870 2398.560 733.150 2398.840 ;
        RECT 834.530 2398.560 834.810 2398.840 ;
        RECT 931.130 2398.560 931.410 2398.840 ;
        RECT 1027.730 2398.560 1028.010 2398.840 ;
        RECT 1124.330 2398.560 1124.610 2398.840 ;
        RECT 1220.930 2398.560 1221.210 2398.840 ;
        RECT 1317.530 2398.560 1317.810 2398.840 ;
        RECT 2124.830 2398.560 2125.110 2398.840 ;
        RECT 2125.750 2398.560 2126.030 2398.840 ;
        RECT 530.930 2397.880 531.210 2398.160 ;
        RECT 772.430 2397.880 772.710 2398.160 ;
        RECT 869.030 2397.880 869.310 2398.160 ;
        RECT 965.630 2397.880 965.910 2398.160 ;
        RECT 1062.230 2397.880 1062.510 2398.160 ;
        RECT 1158.830 2397.880 1159.110 2398.160 ;
        RECT 1255.430 2397.880 1255.710 2398.160 ;
        RECT 1352.030 2397.880 1352.310 2398.160 ;
        RECT 1738.430 2397.880 1738.710 2398.160 ;
        RECT 2269.270 2399.240 2269.550 2399.520 ;
        RECT 2269.270 2398.560 2269.550 2398.840 ;
        RECT 2172.670 2397.880 2172.950 2398.160 ;
        RECT 2414.630 2399.240 2414.910 2399.520 ;
        RECT 2363.570 2396.520 2363.850 2396.800 ;
      LAYER met3 ;
        RECT 2076.710 2401.570 2077.090 2401.580 ;
        RECT 2124.805 2401.570 2125.135 2401.585 ;
        RECT 2076.710 2401.270 2125.135 2401.570 ;
        RECT 2076.710 2401.260 2077.090 2401.270 ;
        RECT 2124.805 2401.255 2125.135 2401.270 ;
        RECT 1738.405 2400.210 1738.735 2400.225 ;
        RECT 2076.710 2400.210 2077.090 2400.220 ;
        RECT 1703.230 2399.910 1738.735 2400.210 ;
        RECT 1441.910 2399.530 1442.290 2399.540 ;
        RECT 544.950 2399.230 641.850 2399.530 ;
        RECT 530.905 2398.170 531.235 2398.185 ;
        RECT 544.950 2398.170 545.250 2399.230 ;
        RECT 530.905 2397.870 545.250 2398.170 ;
        RECT 641.550 2398.170 641.850 2399.230 ;
        RECT 1414.350 2399.230 1442.290 2399.530 ;
        RECT 732.845 2398.850 733.175 2398.865 ;
        RECT 834.505 2398.850 834.835 2398.865 ;
        RECT 931.105 2398.850 931.435 2398.865 ;
        RECT 1027.705 2398.850 1028.035 2398.865 ;
        RECT 1124.305 2398.850 1124.635 2398.865 ;
        RECT 1220.905 2398.850 1221.235 2398.865 ;
        RECT 1317.505 2398.850 1317.835 2398.865 ;
        RECT 690.310 2398.550 733.175 2398.850 ;
        RECT 690.310 2398.170 690.610 2398.550 ;
        RECT 732.845 2398.535 733.175 2398.550 ;
        RECT 786.910 2398.550 834.835 2398.850 ;
        RECT 641.550 2397.870 690.610 2398.170 ;
        RECT 772.405 2398.170 772.735 2398.185 ;
        RECT 786.910 2398.170 787.210 2398.550 ;
        RECT 834.505 2398.535 834.835 2398.550 ;
        RECT 883.510 2398.550 931.435 2398.850 ;
        RECT 772.405 2397.870 787.210 2398.170 ;
        RECT 869.005 2398.170 869.335 2398.185 ;
        RECT 883.510 2398.170 883.810 2398.550 ;
        RECT 931.105 2398.535 931.435 2398.550 ;
        RECT 980.110 2398.550 1028.035 2398.850 ;
        RECT 869.005 2397.870 883.810 2398.170 ;
        RECT 965.605 2398.170 965.935 2398.185 ;
        RECT 980.110 2398.170 980.410 2398.550 ;
        RECT 1027.705 2398.535 1028.035 2398.550 ;
        RECT 1076.710 2398.550 1124.635 2398.850 ;
        RECT 965.605 2397.870 980.410 2398.170 ;
        RECT 1062.205 2398.170 1062.535 2398.185 ;
        RECT 1076.710 2398.170 1077.010 2398.550 ;
        RECT 1124.305 2398.535 1124.635 2398.550 ;
        RECT 1173.310 2398.550 1221.235 2398.850 ;
        RECT 1062.205 2397.870 1077.010 2398.170 ;
        RECT 1158.805 2398.170 1159.135 2398.185 ;
        RECT 1173.310 2398.170 1173.610 2398.550 ;
        RECT 1220.905 2398.535 1221.235 2398.550 ;
        RECT 1269.910 2398.550 1317.835 2398.850 ;
        RECT 1158.805 2397.870 1173.610 2398.170 ;
        RECT 1255.405 2398.170 1255.735 2398.185 ;
        RECT 1269.910 2398.170 1270.210 2398.550 ;
        RECT 1317.505 2398.535 1317.835 2398.550 ;
        RECT 1255.405 2397.870 1270.210 2398.170 ;
        RECT 1352.005 2398.170 1352.335 2398.185 ;
        RECT 1414.350 2398.170 1414.650 2399.230 ;
        RECT 1441.910 2399.220 1442.290 2399.230 ;
        RECT 1510.950 2399.230 1607.850 2399.530 ;
        RECT 1352.005 2397.870 1414.650 2398.170 ;
        RECT 1441.910 2398.170 1442.290 2398.180 ;
        RECT 1510.950 2398.170 1511.250 2399.230 ;
        RECT 1441.910 2397.870 1511.250 2398.170 ;
        RECT 1607.550 2398.170 1607.850 2399.230 ;
        RECT 1703.230 2398.850 1703.530 2399.910 ;
        RECT 1738.405 2399.895 1738.735 2399.910 ;
        RECT 1944.270 2399.910 1995.170 2400.210 ;
        RECT 1656.310 2398.550 1703.530 2398.850 ;
        RECT 1800.750 2399.230 1897.650 2399.530 ;
        RECT 1656.310 2398.170 1656.610 2398.550 ;
        RECT 1607.550 2397.870 1656.610 2398.170 ;
        RECT 1738.405 2398.170 1738.735 2398.185 ;
        RECT 1800.750 2398.170 1801.050 2399.230 ;
        RECT 1897.350 2398.850 1897.650 2399.230 ;
        RECT 1897.350 2398.550 1898.570 2398.850 ;
        RECT 1738.405 2397.870 1801.050 2398.170 ;
        RECT 1898.270 2398.170 1898.570 2398.550 ;
        RECT 1944.270 2398.170 1944.570 2399.910 ;
        RECT 1994.870 2398.850 1995.170 2399.910 ;
        RECT 2041.790 2399.910 2077.090 2400.210 ;
        RECT 2041.790 2398.850 2042.090 2399.910 ;
        RECT 2076.710 2399.900 2077.090 2399.910 ;
        RECT 2269.245 2399.530 2269.575 2399.545 ;
        RECT 2222.110 2399.230 2269.575 2399.530 ;
        RECT 1994.870 2398.550 2042.090 2398.850 ;
        RECT 2124.805 2398.850 2125.135 2398.865 ;
        RECT 2125.725 2398.850 2126.055 2398.865 ;
        RECT 2124.805 2398.550 2126.055 2398.850 ;
        RECT 2124.805 2398.535 2125.135 2398.550 ;
        RECT 2125.725 2398.535 2126.055 2398.550 ;
        RECT 2221.150 2398.850 2221.530 2398.860 ;
        RECT 2222.110 2398.850 2222.410 2399.230 ;
        RECT 2269.245 2399.215 2269.575 2399.230 ;
        RECT 2414.605 2399.530 2414.935 2399.545 ;
        RECT 2604.790 2399.530 2605.170 2399.540 ;
        RECT 2414.605 2399.230 2477.250 2399.530 ;
        RECT 2414.605 2399.215 2414.935 2399.230 ;
        RECT 2221.150 2398.550 2222.410 2398.850 ;
        RECT 2269.245 2398.850 2269.575 2398.865 ;
        RECT 2269.245 2398.550 2339.250 2398.850 ;
        RECT 2221.150 2398.540 2221.530 2398.550 ;
        RECT 2269.245 2398.535 2269.575 2398.550 ;
        RECT 1898.270 2397.870 1944.570 2398.170 ;
        RECT 2172.645 2398.170 2172.975 2398.185 ;
        RECT 2338.950 2398.180 2339.250 2398.550 ;
        RECT 2173.310 2398.170 2173.690 2398.180 ;
        RECT 2172.645 2397.870 2173.690 2398.170 ;
        RECT 530.905 2397.855 531.235 2397.870 ;
        RECT 772.405 2397.855 772.735 2397.870 ;
        RECT 869.005 2397.855 869.335 2397.870 ;
        RECT 965.605 2397.855 965.935 2397.870 ;
        RECT 1062.205 2397.855 1062.535 2397.870 ;
        RECT 1158.805 2397.855 1159.135 2397.870 ;
        RECT 1255.405 2397.855 1255.735 2397.870 ;
        RECT 1352.005 2397.855 1352.335 2397.870 ;
        RECT 1441.910 2397.860 1442.290 2397.870 ;
        RECT 1738.405 2397.855 1738.735 2397.870 ;
        RECT 2172.645 2397.855 2172.975 2397.870 ;
        RECT 2173.310 2397.860 2173.690 2397.870 ;
        RECT 2338.910 2397.860 2339.290 2398.180 ;
        RECT 2476.950 2398.170 2477.250 2399.230 ;
        RECT 2589.190 2399.230 2605.170 2399.530 ;
        RECT 2589.190 2398.170 2589.490 2399.230 ;
        RECT 2604.790 2399.220 2605.170 2399.230 ;
        RECT 2476.950 2397.870 2589.490 2398.170 ;
        RECT 2173.310 2396.810 2173.690 2396.820 ;
        RECT 2221.150 2396.810 2221.530 2396.820 ;
        RECT 2173.310 2396.510 2221.530 2396.810 ;
        RECT 2173.310 2396.500 2173.690 2396.510 ;
        RECT 2221.150 2396.500 2221.530 2396.510 ;
        RECT 2338.910 2396.810 2339.290 2396.820 ;
        RECT 2363.545 2396.810 2363.875 2396.825 ;
        RECT 2338.910 2396.510 2363.875 2396.810 ;
        RECT 2338.910 2396.500 2339.290 2396.510 ;
        RECT 2363.545 2396.495 2363.875 2396.510 ;
        RECT 2604.790 1899.730 2605.170 1899.740 ;
        RECT 2599.460 1899.680 2605.170 1899.730 ;
        RECT 2596.000 1899.430 2605.170 1899.680 ;
        RECT 2596.000 1899.080 2600.000 1899.430 ;
        RECT 2604.790 1899.420 2605.170 1899.430 ;
      LAYER via3 ;
        RECT 2076.740 2401.260 2077.060 2401.580 ;
        RECT 1441.940 2399.220 1442.260 2399.540 ;
        RECT 1441.940 2397.860 1442.260 2398.180 ;
        RECT 2076.740 2399.900 2077.060 2400.220 ;
        RECT 2221.180 2398.540 2221.500 2398.860 ;
        RECT 2173.340 2397.860 2173.660 2398.180 ;
        RECT 2338.940 2397.860 2339.260 2398.180 ;
        RECT 2604.820 2399.220 2605.140 2399.540 ;
        RECT 2173.340 2396.500 2173.660 2396.820 ;
        RECT 2221.180 2396.500 2221.500 2396.820 ;
        RECT 2338.940 2396.500 2339.260 2396.820 ;
        RECT 2604.820 1899.420 2605.140 1899.740 ;
      LAYER met4 ;
        RECT 2076.735 2401.255 2077.065 2401.585 ;
        RECT 2076.750 2400.225 2077.050 2401.255 ;
        RECT 2076.735 2399.895 2077.065 2400.225 ;
        RECT 1441.935 2399.215 1442.265 2399.545 ;
        RECT 2604.815 2399.215 2605.145 2399.545 ;
        RECT 1441.950 2398.185 1442.250 2399.215 ;
        RECT 2221.175 2398.535 2221.505 2398.865 ;
        RECT 1441.935 2397.855 1442.265 2398.185 ;
        RECT 2173.335 2397.855 2173.665 2398.185 ;
        RECT 2173.350 2396.825 2173.650 2397.855 ;
        RECT 2221.190 2396.825 2221.490 2398.535 ;
        RECT 2338.935 2397.855 2339.265 2398.185 ;
        RECT 2338.950 2396.825 2339.250 2397.855 ;
        RECT 2173.335 2396.495 2173.665 2396.825 ;
        RECT 2221.175 2396.495 2221.505 2396.825 ;
        RECT 2338.935 2396.495 2339.265 2396.825 ;
        RECT 2604.830 1899.745 2605.130 2399.215 ;
        RECT 2604.815 1899.415 2605.145 1899.745 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 2397.525 206.840 3501.670 ;
        RECT 206.630 2397.155 206.910 2397.525 ;
      LAYER via2 ;
        RECT 206.630 2397.200 206.910 2397.480 ;
      LAYER met3 ;
        RECT 2598.350 2397.860 2598.730 2398.180 ;
        RECT 206.605 2397.490 206.935 2397.505 ;
        RECT 2598.390 2397.490 2598.690 2397.860 ;
        RECT 206.605 2397.190 2598.690 2397.490 ;
        RECT 206.605 2397.175 206.935 2397.190 ;
        RECT 2598.350 1932.060 2598.730 1932.380 ;
        RECT 2598.390 1931.640 2598.690 1932.060 ;
        RECT 2596.000 1931.040 2600.000 1931.640 ;
      LAYER via3 ;
        RECT 2598.380 2397.860 2598.700 2398.180 ;
        RECT 2598.380 1932.060 2598.700 1932.380 ;
      LAYER met4 ;
        RECT 2598.375 2397.855 2598.705 2398.185 ;
        RECT 2598.390 1932.385 2598.690 2397.855 ;
        RECT 2598.375 1932.055 2598.705 1932.385 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT -4.800 3411.070 3.370 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 3.070 3409.330 3.370 3411.070 ;
        RECT 2596.510 3409.330 2596.890 3409.340 ;
        RECT 3.070 3409.030 2596.890 3409.330 ;
        RECT 2596.510 3409.020 2596.890 3409.030 ;
        RECT 2596.510 1965.380 2596.890 1965.700 ;
        RECT 2596.550 1962.920 2596.850 1965.380 ;
        RECT 2596.000 1962.320 2600.000 1962.920 ;
      LAYER via3 ;
        RECT 2596.540 3409.020 2596.860 3409.340 ;
        RECT 2596.540 1965.380 2596.860 1965.700 ;
      LAYER met4 ;
        RECT 2596.535 3409.015 2596.865 3409.345 ;
        RECT 2596.550 1965.705 2596.850 3409.015 ;
        RECT 2596.535 1965.375 2596.865 1965.705 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3119.060 17.410 3119.120 ;
        RECT 2598.610 3119.060 2598.930 3119.120 ;
        RECT 17.090 3118.920 2598.930 3119.060 ;
        RECT 17.090 3118.860 17.410 3118.920 ;
        RECT 2598.610 3118.860 2598.930 3118.920 ;
      LAYER via ;
        RECT 17.120 3118.860 17.380 3119.120 ;
        RECT 2598.640 3118.860 2598.900 3119.120 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.150 17.320 3124.075 ;
        RECT 17.120 3118.830 17.380 3119.150 ;
        RECT 2598.640 3118.830 2598.900 3119.150 ;
        RECT 2598.700 1997.685 2598.840 3118.830 ;
        RECT 2598.630 1997.315 2598.910 1997.685 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
        RECT 2598.630 1997.360 2598.910 1997.640 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
        RECT 2598.605 1997.650 2598.935 1997.665 ;
        RECT 2598.390 1997.335 2598.935 1997.650 ;
        RECT 2598.390 1994.880 2598.690 1997.335 ;
        RECT 2596.000 1994.280 2600.000 1994.880 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 2398.600 18.330 2398.660 ;
        RECT 2606.890 2398.600 2607.210 2398.660 ;
        RECT 18.010 2398.460 2607.210 2398.600 ;
        RECT 18.010 2398.400 18.330 2398.460 ;
        RECT 2606.890 2398.400 2607.210 2398.460 ;
      LAYER via ;
        RECT 18.040 2398.400 18.300 2398.660 ;
        RECT 2606.920 2398.400 2607.180 2398.660 ;
      LAYER met2 ;
        RECT 18.030 2836.435 18.310 2836.805 ;
        RECT 18.100 2398.690 18.240 2836.435 ;
        RECT 18.040 2398.370 18.300 2398.690 ;
        RECT 2606.920 2398.370 2607.180 2398.690 ;
        RECT 2606.980 2026.245 2607.120 2398.370 ;
        RECT 2606.910 2025.875 2607.190 2026.245 ;
      LAYER via2 ;
        RECT 18.030 2836.480 18.310 2836.760 ;
        RECT 2606.910 2025.920 2607.190 2026.200 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 18.005 2836.770 18.335 2836.785 ;
        RECT -4.800 2836.470 18.335 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 18.005 2836.455 18.335 2836.470 ;
        RECT 2606.885 2026.210 2607.215 2026.225 ;
        RECT 2599.460 2026.160 2607.215 2026.210 ;
        RECT 2596.000 2025.910 2607.215 2026.160 ;
        RECT 2596.000 2025.560 2600.000 2025.910 ;
        RECT 2606.885 2025.895 2607.215 2025.910 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 2546.500 16.950 2546.560 ;
        RECT 2599.990 2546.500 2600.310 2546.560 ;
        RECT 16.630 2546.360 2600.310 2546.500 ;
        RECT 16.630 2546.300 16.950 2546.360 ;
        RECT 2599.990 2546.300 2600.310 2546.360 ;
      LAYER via ;
        RECT 16.660 2546.300 16.920 2546.560 ;
        RECT 2600.020 2546.300 2600.280 2546.560 ;
      LAYER met2 ;
        RECT 16.650 2549.475 16.930 2549.845 ;
        RECT 16.720 2546.590 16.860 2549.475 ;
        RECT 16.660 2546.270 16.920 2546.590 ;
        RECT 2600.020 2546.270 2600.280 2546.590 ;
        RECT 2600.080 2060.925 2600.220 2546.270 ;
        RECT 2600.010 2060.555 2600.290 2060.925 ;
      LAYER via2 ;
        RECT 16.650 2549.520 16.930 2549.800 ;
        RECT 2600.010 2060.600 2600.290 2060.880 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 16.625 2549.810 16.955 2549.825 ;
        RECT -4.800 2549.510 16.955 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 16.625 2549.495 16.955 2549.510 ;
        RECT 2599.985 2060.890 2600.315 2060.905 ;
        RECT 2599.310 2060.590 2600.315 2060.890 ;
        RECT 2599.310 2058.120 2599.610 2060.590 ;
        RECT 2599.985 2060.575 2600.315 2060.590 ;
        RECT 2596.000 2057.520 2600.000 2058.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1395.710 2396.220 1396.030 2396.280 ;
        RECT 2599.530 2396.220 2599.850 2396.280 ;
        RECT 1395.710 2396.080 2599.850 2396.220 ;
        RECT 1395.710 2396.020 1396.030 2396.080 ;
        RECT 2599.530 2396.020 2599.850 2396.080 ;
        RECT 17.550 2262.940 17.870 2263.000 ;
        RECT 1395.710 2262.940 1396.030 2263.000 ;
        RECT 17.550 2262.800 1396.030 2262.940 ;
        RECT 17.550 2262.740 17.870 2262.800 ;
        RECT 1395.710 2262.740 1396.030 2262.800 ;
      LAYER via ;
        RECT 1395.740 2396.020 1396.000 2396.280 ;
        RECT 2599.560 2396.020 2599.820 2396.280 ;
        RECT 17.580 2262.740 17.840 2263.000 ;
        RECT 1395.740 2262.740 1396.000 2263.000 ;
      LAYER met2 ;
        RECT 1395.740 2395.990 1396.000 2396.310 ;
        RECT 2599.560 2395.990 2599.820 2396.310 ;
        RECT 1395.800 2263.030 1395.940 2395.990 ;
        RECT 2599.620 2381.205 2599.760 2395.990 ;
        RECT 2599.550 2380.835 2599.830 2381.205 ;
        RECT 2600.930 2379.475 2601.210 2379.845 ;
        RECT 17.580 2262.710 17.840 2263.030 ;
        RECT 1395.740 2262.710 1396.000 2263.030 ;
        RECT 17.640 2262.205 17.780 2262.710 ;
        RECT 17.570 2261.835 17.850 2262.205 ;
        RECT 2601.000 2089.485 2601.140 2379.475 ;
        RECT 2600.930 2089.115 2601.210 2089.485 ;
      LAYER via2 ;
        RECT 2599.550 2380.880 2599.830 2381.160 ;
        RECT 2600.930 2379.520 2601.210 2379.800 ;
        RECT 17.570 2261.880 17.850 2262.160 ;
        RECT 2600.930 2089.160 2601.210 2089.440 ;
      LAYER met3 ;
        RECT 2599.525 2381.170 2599.855 2381.185 ;
        RECT 2600.190 2381.170 2600.570 2381.180 ;
        RECT 2599.525 2380.870 2600.570 2381.170 ;
        RECT 2599.525 2380.855 2599.855 2380.870 ;
        RECT 2600.190 2380.860 2600.570 2380.870 ;
        RECT 2600.190 2379.810 2600.570 2379.820 ;
        RECT 2600.905 2379.810 2601.235 2379.825 ;
        RECT 2600.190 2379.510 2601.235 2379.810 ;
        RECT 2600.190 2379.500 2600.570 2379.510 ;
        RECT 2600.905 2379.495 2601.235 2379.510 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.545 2262.170 17.875 2262.185 ;
        RECT -4.800 2261.870 17.875 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.545 2261.855 17.875 2261.870 ;
        RECT 2600.905 2089.450 2601.235 2089.465 ;
        RECT 2599.460 2089.400 2601.235 2089.450 ;
        RECT 2596.000 2089.150 2601.235 2089.400 ;
        RECT 2596.000 2088.800 2600.000 2089.150 ;
        RECT 2600.905 2089.135 2601.235 2089.150 ;
      LAYER via3 ;
        RECT 2600.220 2380.860 2600.540 2381.180 ;
        RECT 2600.220 2379.500 2600.540 2379.820 ;
      LAYER met4 ;
        RECT 2600.215 2380.855 2600.545 2381.185 ;
        RECT 2600.230 2379.825 2600.530 2380.855 ;
        RECT 2600.215 2379.495 2600.545 2379.825 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 2396.560 1400.630 2396.620 ;
        RECT 2604.590 2396.560 2604.910 2396.620 ;
        RECT 1400.310 2396.420 2604.910 2396.560 ;
        RECT 1400.310 2396.360 1400.630 2396.420 ;
        RECT 2604.590 2396.360 2604.910 2396.420 ;
        RECT 15.710 1980.060 16.030 1980.120 ;
        RECT 1400.310 1980.060 1400.630 1980.120 ;
        RECT 15.710 1979.920 1400.630 1980.060 ;
        RECT 15.710 1979.860 16.030 1979.920 ;
        RECT 1400.310 1979.860 1400.630 1979.920 ;
      LAYER via ;
        RECT 1400.340 2396.360 1400.600 2396.620 ;
        RECT 2604.620 2396.360 2604.880 2396.620 ;
        RECT 15.740 1979.860 16.000 1980.120 ;
        RECT 1400.340 1979.860 1400.600 1980.120 ;
      LAYER met2 ;
        RECT 1400.340 2396.330 1400.600 2396.650 ;
        RECT 2604.620 2396.330 2604.880 2396.650 ;
        RECT 1400.400 1980.150 1400.540 2396.330 ;
        RECT 2604.680 2120.765 2604.820 2396.330 ;
        RECT 2604.610 2120.395 2604.890 2120.765 ;
        RECT 15.740 1979.830 16.000 1980.150 ;
        RECT 1400.340 1979.830 1400.600 1980.150 ;
        RECT 15.800 1975.245 15.940 1979.830 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 2604.610 2120.440 2604.890 2120.720 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT 2604.585 2120.730 2604.915 2120.745 ;
        RECT 2599.460 2120.680 2604.915 2120.730 ;
        RECT 2596.000 2120.430 2604.915 2120.680 ;
        RECT 2596.000 2120.080 2600.000 2120.430 ;
        RECT 2604.585 2120.415 2604.915 2120.430 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2618.390 558.860 2618.710 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2618.390 558.720 2899.310 558.860 ;
        RECT 2618.390 558.660 2618.710 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2618.420 558.660 2618.680 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2618.410 1267.675 2618.690 1268.045 ;
        RECT 2618.480 558.950 2618.620 1267.675 ;
        RECT 2618.420 558.630 2618.680 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2618.410 1267.720 2618.690 1268.000 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2618.385 1268.010 2618.715 1268.025 ;
        RECT 2599.460 1267.960 2618.715 1268.010 ;
        RECT 2596.000 1267.710 2618.715 1267.960 ;
        RECT 2596.000 1267.360 2600.000 1267.710 ;
        RECT 2618.385 1267.695 2618.715 1267.710 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1398.930 2393.160 1399.250 2393.220 ;
        RECT 2608.270 2393.160 2608.590 2393.220 ;
        RECT 1398.930 2393.020 2608.590 2393.160 ;
        RECT 1398.930 2392.960 1399.250 2393.020 ;
        RECT 2608.270 2392.960 2608.590 2393.020 ;
        RECT 2608.270 2331.760 2608.590 2332.020 ;
        RECT 2608.360 2331.000 2608.500 2331.760 ;
        RECT 2608.270 2330.740 2608.590 2331.000 ;
        RECT 17.550 1690.380 17.870 1690.440 ;
        RECT 1398.930 1690.380 1399.250 1690.440 ;
        RECT 17.550 1690.240 1399.250 1690.380 ;
        RECT 17.550 1690.180 17.870 1690.240 ;
        RECT 1398.930 1690.180 1399.250 1690.240 ;
      LAYER via ;
        RECT 1398.960 2392.960 1399.220 2393.220 ;
        RECT 2608.300 2392.960 2608.560 2393.220 ;
        RECT 2608.300 2331.760 2608.560 2332.020 ;
        RECT 2608.300 2330.740 2608.560 2331.000 ;
        RECT 17.580 1690.180 17.840 1690.440 ;
        RECT 1398.960 1690.180 1399.220 1690.440 ;
      LAYER met2 ;
        RECT 1398.960 2392.930 1399.220 2393.250 ;
        RECT 2608.300 2392.930 2608.560 2393.250 ;
        RECT 1399.020 1690.470 1399.160 2392.930 ;
        RECT 2608.360 2332.050 2608.500 2392.930 ;
        RECT 2608.300 2331.730 2608.560 2332.050 ;
        RECT 2608.300 2330.710 2608.560 2331.030 ;
        RECT 2608.360 2152.725 2608.500 2330.710 ;
        RECT 2608.290 2152.355 2608.570 2152.725 ;
        RECT 17.580 1690.150 17.840 1690.470 ;
        RECT 1398.960 1690.150 1399.220 1690.470 ;
        RECT 17.640 1687.605 17.780 1690.150 ;
        RECT 17.570 1687.235 17.850 1687.605 ;
      LAYER via2 ;
        RECT 2608.290 2152.400 2608.570 2152.680 ;
        RECT 17.570 1687.280 17.850 1687.560 ;
      LAYER met3 ;
        RECT 2608.265 2152.690 2608.595 2152.705 ;
        RECT 2599.460 2152.640 2608.595 2152.690 ;
        RECT 2596.000 2152.390 2608.595 2152.640 ;
        RECT 2596.000 2152.040 2600.000 2152.390 ;
        RECT 2608.265 2152.375 2608.595 2152.390 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.545 1687.570 17.875 1687.585 ;
        RECT -4.800 1687.270 17.875 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.545 1687.255 17.875 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1397.550 2392.820 1397.870 2392.880 ;
        RECT 2614.250 2392.820 2614.570 2392.880 ;
        RECT 1397.550 2392.680 2614.570 2392.820 ;
        RECT 1397.550 2392.620 1397.870 2392.680 ;
        RECT 2614.250 2392.620 2614.570 2392.680 ;
        RECT 15.250 1476.520 15.570 1476.580 ;
        RECT 1397.550 1476.520 1397.870 1476.580 ;
        RECT 15.250 1476.380 1397.870 1476.520 ;
        RECT 15.250 1476.320 15.570 1476.380 ;
        RECT 1397.550 1476.320 1397.870 1476.380 ;
      LAYER via ;
        RECT 1397.580 2392.620 1397.840 2392.880 ;
        RECT 2614.280 2392.620 2614.540 2392.880 ;
        RECT 15.280 1476.320 15.540 1476.580 ;
        RECT 1397.580 1476.320 1397.840 1476.580 ;
      LAYER met2 ;
        RECT 1397.580 2392.590 1397.840 2392.910 ;
        RECT 2614.280 2392.590 2614.540 2392.910 ;
        RECT 1397.640 1476.610 1397.780 2392.590 ;
        RECT 2614.340 2184.005 2614.480 2392.590 ;
        RECT 2614.270 2183.635 2614.550 2184.005 ;
        RECT 15.280 1476.290 15.540 1476.610 ;
        RECT 1397.580 1476.290 1397.840 1476.610 ;
        RECT 15.340 1472.045 15.480 1476.290 ;
        RECT 15.270 1471.675 15.550 1472.045 ;
      LAYER via2 ;
        RECT 2614.270 2183.680 2614.550 2183.960 ;
        RECT 15.270 1471.720 15.550 1472.000 ;
      LAYER met3 ;
        RECT 2614.245 2183.970 2614.575 2183.985 ;
        RECT 2599.460 2183.920 2614.575 2183.970 ;
        RECT 2596.000 2183.670 2614.575 2183.920 ;
        RECT 2596.000 2183.320 2600.000 2183.670 ;
        RECT 2614.245 2183.655 2614.575 2183.670 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 15.245 1472.010 15.575 1472.025 ;
        RECT -4.800 1471.710 15.575 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 15.245 1471.695 15.575 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 1203.840 18.330 1203.900 ;
        RECT 2607.810 1203.840 2608.130 1203.900 ;
        RECT 18.010 1203.700 2608.130 1203.840 ;
        RECT 18.010 1203.640 18.330 1203.700 ;
        RECT 2607.810 1203.640 2608.130 1203.700 ;
      LAYER via ;
        RECT 18.040 1203.640 18.300 1203.900 ;
        RECT 2607.840 1203.640 2608.100 1203.900 ;
      LAYER met2 ;
        RECT 2607.830 2208.115 2608.110 2208.485 ;
        RECT 18.030 1256.115 18.310 1256.485 ;
        RECT 18.100 1203.930 18.240 1256.115 ;
        RECT 2607.900 1203.930 2608.040 2208.115 ;
        RECT 18.040 1203.610 18.300 1203.930 ;
        RECT 2607.840 1203.610 2608.100 1203.930 ;
      LAYER via2 ;
        RECT 2607.830 2208.160 2608.110 2208.440 ;
        RECT 18.030 1256.160 18.310 1256.440 ;
      LAYER met3 ;
        RECT 2606.630 2215.930 2607.010 2215.940 ;
        RECT 2599.460 2215.880 2607.010 2215.930 ;
        RECT 2596.000 2215.630 2607.010 2215.880 ;
        RECT 2596.000 2215.280 2600.000 2215.630 ;
        RECT 2606.630 2215.620 2607.010 2215.630 ;
        RECT 2606.630 2208.450 2607.010 2208.460 ;
        RECT 2607.805 2208.450 2608.135 2208.465 ;
        RECT 2606.630 2208.150 2608.135 2208.450 ;
        RECT 2606.630 2208.140 2607.010 2208.150 ;
        RECT 2607.805 2208.135 2608.135 2208.150 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 18.005 1256.450 18.335 1256.465 ;
        RECT -4.800 1256.150 18.335 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 18.005 1256.135 18.335 1256.150 ;
      LAYER via3 ;
        RECT 2606.660 2215.620 2606.980 2215.940 ;
        RECT 2606.660 2208.140 2606.980 2208.460 ;
      LAYER met4 ;
        RECT 2606.655 2215.615 2606.985 2215.945 ;
        RECT 2606.670 2208.465 2606.970 2215.615 ;
        RECT 2606.655 2208.135 2606.985 2208.465 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 1041.660 17.870 1041.720 ;
        RECT 2611.030 1041.660 2611.350 1041.720 ;
        RECT 17.550 1041.520 2611.350 1041.660 ;
        RECT 17.550 1041.460 17.870 1041.520 ;
        RECT 2611.030 1041.460 2611.350 1041.520 ;
      LAYER via ;
        RECT 17.580 1041.460 17.840 1041.720 ;
        RECT 2611.060 1041.460 2611.320 1041.720 ;
      LAYER met2 ;
        RECT 2611.050 2246.875 2611.330 2247.245 ;
        RECT 2611.120 1041.750 2611.260 2246.875 ;
        RECT 17.580 1041.430 17.840 1041.750 ;
        RECT 2611.060 1041.430 2611.320 1041.750 ;
        RECT 17.640 1040.925 17.780 1041.430 ;
        RECT 17.570 1040.555 17.850 1040.925 ;
      LAYER via2 ;
        RECT 2611.050 2246.920 2611.330 2247.200 ;
        RECT 17.570 1040.600 17.850 1040.880 ;
      LAYER met3 ;
        RECT 2611.025 2247.210 2611.355 2247.225 ;
        RECT 2599.460 2247.160 2611.355 2247.210 ;
        RECT 2596.000 2246.910 2611.355 2247.160 ;
        RECT 2596.000 2246.560 2600.000 2246.910 ;
        RECT 2611.025 2246.895 2611.355 2246.910 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.545 1040.890 17.875 1040.905 ;
        RECT -4.800 1040.590 17.875 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.545 1040.575 17.875 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.930 1004.940 19.250 1005.000 ;
        RECT 2609.650 1004.940 2609.970 1005.000 ;
        RECT 18.930 1004.800 2609.970 1004.940 ;
        RECT 18.930 1004.740 19.250 1004.800 ;
        RECT 2609.650 1004.740 2609.970 1004.800 ;
      LAYER via ;
        RECT 18.960 1004.740 19.220 1005.000 ;
        RECT 2609.680 1004.740 2609.940 1005.000 ;
      LAYER met2 ;
        RECT 2609.670 2278.835 2609.950 2279.205 ;
        RECT 2609.740 1005.030 2609.880 2278.835 ;
        RECT 18.960 1004.710 19.220 1005.030 ;
        RECT 2609.680 1004.710 2609.940 1005.030 ;
        RECT 19.020 825.365 19.160 1004.710 ;
        RECT 18.950 824.995 19.230 825.365 ;
      LAYER via2 ;
        RECT 2609.670 2278.880 2609.950 2279.160 ;
        RECT 18.950 825.040 19.230 825.320 ;
      LAYER met3 ;
        RECT 2609.645 2279.170 2609.975 2279.185 ;
        RECT 2599.460 2279.120 2609.975 2279.170 ;
        RECT 2596.000 2278.870 2609.975 2279.120 ;
        RECT 2596.000 2278.520 2600.000 2278.870 ;
        RECT 2609.645 2278.855 2609.975 2278.870 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 18.925 825.330 19.255 825.345 ;
        RECT -4.800 825.030 19.255 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 18.925 825.015 19.255 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 1004.600 17.870 1004.660 ;
        RECT 2614.710 1004.600 2615.030 1004.660 ;
        RECT 17.550 1004.460 2615.030 1004.600 ;
        RECT 17.550 1004.400 17.870 1004.460 ;
        RECT 2614.710 1004.400 2615.030 1004.460 ;
      LAYER via ;
        RECT 17.580 1004.400 17.840 1004.660 ;
        RECT 2614.740 1004.400 2615.000 1004.660 ;
      LAYER met2 ;
        RECT 2614.730 2310.115 2615.010 2310.485 ;
        RECT 2614.800 1004.690 2614.940 2310.115 ;
        RECT 17.580 1004.370 17.840 1004.690 ;
        RECT 2614.740 1004.370 2615.000 1004.690 ;
        RECT 17.640 610.485 17.780 1004.370 ;
        RECT 17.570 610.115 17.850 610.485 ;
      LAYER via2 ;
        RECT 2614.730 2310.160 2615.010 2310.440 ;
        RECT 17.570 610.160 17.850 610.440 ;
      LAYER met3 ;
        RECT 2614.705 2310.450 2615.035 2310.465 ;
        RECT 2599.460 2310.400 2615.035 2310.450 ;
        RECT 2596.000 2310.150 2615.035 2310.400 ;
        RECT 2596.000 2309.800 2600.000 2310.150 ;
        RECT 2614.705 2310.135 2615.035 2310.150 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.545 610.450 17.875 610.465 ;
        RECT -4.800 610.150 17.875 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.545 610.135 17.875 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 399.995 17.850 400.365 ;
        RECT 17.640 394.925 17.780 399.995 ;
        RECT 17.570 394.555 17.850 394.925 ;
      LAYER via2 ;
        RECT 17.570 400.040 17.850 400.320 ;
        RECT 17.570 394.600 17.850 394.880 ;
      LAYER met3 ;
        RECT 2611.230 2342.410 2611.610 2342.420 ;
        RECT 2599.460 2342.360 2611.610 2342.410 ;
        RECT 2596.000 2342.110 2611.610 2342.360 ;
        RECT 2596.000 2341.760 2600.000 2342.110 ;
        RECT 2611.230 2342.100 2611.610 2342.110 ;
        RECT 17.545 400.330 17.875 400.345 ;
        RECT 2611.230 400.330 2611.610 400.340 ;
        RECT 17.545 400.030 2611.610 400.330 ;
        RECT 17.545 400.015 17.875 400.030 ;
        RECT 2611.230 400.020 2611.610 400.030 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.545 394.890 17.875 394.905 ;
        RECT -4.800 394.590 17.875 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.545 394.575 17.875 394.590 ;
      LAYER via3 ;
        RECT 2611.260 2342.100 2611.580 2342.420 ;
        RECT 2611.260 400.020 2611.580 400.340 ;
      LAYER met4 ;
        RECT 2611.255 2342.095 2611.585 2342.425 ;
        RECT 2611.270 400.345 2611.570 2342.095 ;
        RECT 2611.255 400.015 2611.585 400.345 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2609.390 2373.690 2609.770 2373.700 ;
        RECT 2599.460 2373.640 2609.770 2373.690 ;
        RECT 2596.000 2373.390 2609.770 2373.640 ;
        RECT 2596.000 2373.040 2600.000 2373.390 ;
        RECT 2609.390 2373.380 2609.770 2373.390 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 2609.390 179.330 2609.770 179.340 ;
        RECT -4.800 179.030 2609.770 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 2609.390 179.020 2609.770 179.030 ;
      LAYER via3 ;
        RECT 2609.420 2373.380 2609.740 2373.700 ;
        RECT 2609.420 179.020 2609.740 179.340 ;
      LAYER met4 ;
        RECT 2609.415 2373.375 2609.745 2373.705 ;
        RECT 2609.430 179.345 2609.730 2373.375 ;
        RECT 2609.415 179.015 2609.745 179.345 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2613.790 1297.340 2614.110 1297.400 ;
        RECT 2618.850 1297.340 2619.170 1297.400 ;
        RECT 2613.790 1297.200 2619.170 1297.340 ;
        RECT 2613.790 1297.140 2614.110 1297.200 ;
        RECT 2618.850 1297.140 2619.170 1297.200 ;
        RECT 2618.850 793.460 2619.170 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2618.850 793.320 2899.310 793.460 ;
        RECT 2618.850 793.260 2619.170 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2613.820 1297.140 2614.080 1297.400 ;
        RECT 2618.880 1297.140 2619.140 1297.400 ;
        RECT 2618.880 793.260 2619.140 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2613.810 1299.635 2614.090 1300.005 ;
        RECT 2613.880 1297.430 2614.020 1299.635 ;
        RECT 2613.820 1297.110 2614.080 1297.430 ;
        RECT 2618.880 1297.110 2619.140 1297.430 ;
        RECT 2618.940 793.550 2619.080 1297.110 ;
        RECT 2618.880 793.230 2619.140 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2613.810 1299.680 2614.090 1299.960 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2613.785 1299.970 2614.115 1299.985 ;
        RECT 2599.460 1299.920 2614.115 1299.970 ;
        RECT 2596.000 1299.670 2614.115 1299.920 ;
        RECT 2596.000 1299.320 2600.000 1299.670 ;
        RECT 2613.785 1299.655 2614.115 1299.670 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2613.790 1324.880 2614.110 1324.940 ;
        RECT 2620.230 1324.880 2620.550 1324.940 ;
        RECT 2613.790 1324.740 2620.550 1324.880 ;
        RECT 2613.790 1324.680 2614.110 1324.740 ;
        RECT 2620.230 1324.680 2620.550 1324.740 ;
        RECT 2620.230 1028.060 2620.550 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 2620.230 1027.920 2899.310 1028.060 ;
        RECT 2620.230 1027.860 2620.550 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 2613.820 1324.680 2614.080 1324.940 ;
        RECT 2620.260 1324.680 2620.520 1324.940 ;
        RECT 2620.260 1027.860 2620.520 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 2613.810 1330.915 2614.090 1331.285 ;
        RECT 2613.880 1324.970 2614.020 1330.915 ;
        RECT 2613.820 1324.650 2614.080 1324.970 ;
        RECT 2620.260 1324.650 2620.520 1324.970 ;
        RECT 2620.320 1028.150 2620.460 1324.650 ;
        RECT 2620.260 1027.830 2620.520 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2613.810 1330.960 2614.090 1331.240 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 2613.785 1331.250 2614.115 1331.265 ;
        RECT 2599.460 1331.200 2614.115 1331.250 ;
        RECT 2596.000 1330.950 2614.115 1331.200 ;
        RECT 2596.000 1330.600 2600.000 1330.950 ;
        RECT 2613.785 1330.935 2614.115 1330.950 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2608.270 1262.660 2608.590 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 2608.270 1262.520 2899.310 1262.660 ;
        RECT 2608.270 1262.460 2608.590 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 2608.300 1262.460 2608.560 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 2608.290 1362.875 2608.570 1363.245 ;
        RECT 2608.360 1262.750 2608.500 1362.875 ;
        RECT 2608.300 1262.430 2608.560 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 2608.290 1362.920 2608.570 1363.200 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 2608.265 1363.210 2608.595 1363.225 ;
        RECT 2599.460 1363.160 2608.595 1363.210 ;
        RECT 2596.000 1362.910 2608.595 1363.160 ;
        RECT 2596.000 1362.560 2600.000 1362.910 ;
        RECT 2608.265 1362.895 2608.595 1362.910 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2612.870 1473.120 2613.190 1473.180 ;
        RECT 2899.910 1473.120 2900.230 1473.180 ;
        RECT 2612.870 1472.980 2900.230 1473.120 ;
        RECT 2612.870 1472.920 2613.190 1472.980 ;
        RECT 2899.910 1472.920 2900.230 1472.980 ;
      LAYER via ;
        RECT 2612.900 1472.920 2613.160 1473.180 ;
        RECT 2899.940 1472.920 2900.200 1473.180 ;
      LAYER met2 ;
        RECT 2899.930 1495.475 2900.210 1495.845 ;
        RECT 2900.000 1473.210 2900.140 1495.475 ;
        RECT 2612.900 1472.890 2613.160 1473.210 ;
        RECT 2899.940 1472.890 2900.200 1473.210 ;
        RECT 2612.960 1394.525 2613.100 1472.890 ;
        RECT 2612.890 1394.155 2613.170 1394.525 ;
      LAYER via2 ;
        RECT 2899.930 1495.520 2900.210 1495.800 ;
        RECT 2612.890 1394.200 2613.170 1394.480 ;
      LAYER met3 ;
        RECT 2899.905 1495.810 2900.235 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2899.905 1495.510 2924.800 1495.810 ;
        RECT 2899.905 1495.495 2900.235 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2612.865 1394.490 2613.195 1394.505 ;
        RECT 2599.460 1394.440 2613.195 1394.490 ;
        RECT 2596.000 1394.190 2613.195 1394.440 ;
        RECT 2596.000 1393.840 2600.000 1394.190 ;
        RECT 2612.865 1394.175 2613.195 1394.190 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2614.250 1428.240 2614.570 1428.300 ;
        RECT 2902.670 1428.240 2902.990 1428.300 ;
        RECT 2614.250 1428.100 2902.990 1428.240 ;
        RECT 2614.250 1428.040 2614.570 1428.100 ;
        RECT 2902.670 1428.040 2902.990 1428.100 ;
      LAYER via ;
        RECT 2614.280 1428.040 2614.540 1428.300 ;
        RECT 2902.700 1428.040 2902.960 1428.300 ;
      LAYER met2 ;
        RECT 2902.690 1730.075 2902.970 1730.445 ;
        RECT 2902.760 1428.330 2902.900 1730.075 ;
        RECT 2614.280 1428.010 2614.540 1428.330 ;
        RECT 2902.700 1428.010 2902.960 1428.330 ;
        RECT 2614.340 1426.485 2614.480 1428.010 ;
        RECT 2614.270 1426.115 2614.550 1426.485 ;
      LAYER via2 ;
        RECT 2902.690 1730.120 2902.970 1730.400 ;
        RECT 2614.270 1426.160 2614.550 1426.440 ;
      LAYER met3 ;
        RECT 2902.665 1730.410 2902.995 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2902.665 1730.110 2924.800 1730.410 ;
        RECT 2902.665 1730.095 2902.995 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2614.245 1426.450 2614.575 1426.465 ;
        RECT 2599.460 1426.400 2614.575 1426.450 ;
        RECT 2596.000 1426.150 2614.575 1426.400 ;
        RECT 2596.000 1425.800 2600.000 1426.150 ;
        RECT 2614.245 1426.135 2614.575 1426.150 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2619.770 1960.000 2620.090 1960.060 ;
        RECT 2899.450 1960.000 2899.770 1960.060 ;
        RECT 2619.770 1959.860 2899.770 1960.000 ;
        RECT 2619.770 1959.800 2620.090 1959.860 ;
        RECT 2899.450 1959.800 2899.770 1959.860 ;
        RECT 2608.270 1457.820 2608.590 1457.880 ;
        RECT 2619.770 1457.820 2620.090 1457.880 ;
        RECT 2608.270 1457.680 2620.090 1457.820 ;
        RECT 2608.270 1457.620 2608.590 1457.680 ;
        RECT 2619.770 1457.620 2620.090 1457.680 ;
      LAYER via ;
        RECT 2619.800 1959.800 2620.060 1960.060 ;
        RECT 2899.480 1959.800 2899.740 1960.060 ;
        RECT 2608.300 1457.620 2608.560 1457.880 ;
        RECT 2619.800 1457.620 2620.060 1457.880 ;
      LAYER met2 ;
        RECT 2899.470 1964.675 2899.750 1965.045 ;
        RECT 2899.540 1960.090 2899.680 1964.675 ;
        RECT 2619.800 1959.770 2620.060 1960.090 ;
        RECT 2899.480 1959.770 2899.740 1960.090 ;
        RECT 2619.860 1457.910 2620.000 1959.770 ;
        RECT 2608.300 1457.765 2608.560 1457.910 ;
        RECT 2608.290 1457.395 2608.570 1457.765 ;
        RECT 2619.800 1457.590 2620.060 1457.910 ;
      LAYER via2 ;
        RECT 2899.470 1964.720 2899.750 1965.000 ;
        RECT 2608.290 1457.440 2608.570 1457.720 ;
      LAYER met3 ;
        RECT 2899.445 1965.010 2899.775 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2899.445 1964.710 2924.800 1965.010 ;
        RECT 2899.445 1964.695 2899.775 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2608.265 1457.730 2608.595 1457.745 ;
        RECT 2599.460 1457.680 2608.595 1457.730 ;
        RECT 2596.000 1457.430 2608.595 1457.680 ;
        RECT 2596.000 1457.080 2600.000 1457.430 ;
        RECT 2608.265 1457.415 2608.595 1457.430 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2673.590 2194.600 2673.910 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2673.590 2194.460 2901.150 2194.600 ;
        RECT 2673.590 2194.400 2673.910 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
        RECT 2614.250 1490.460 2614.570 1490.520 ;
        RECT 2673.590 1490.460 2673.910 1490.520 ;
        RECT 2614.250 1490.320 2673.910 1490.460 ;
        RECT 2614.250 1490.260 2614.570 1490.320 ;
        RECT 2673.590 1490.260 2673.910 1490.320 ;
      LAYER via ;
        RECT 2673.620 2194.400 2673.880 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
        RECT 2614.280 1490.260 2614.540 1490.520 ;
        RECT 2673.620 1490.260 2673.880 1490.520 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2673.620 2194.370 2673.880 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2673.680 1490.550 2673.820 2194.370 ;
        RECT 2614.280 1490.230 2614.540 1490.550 ;
        RECT 2673.620 1490.230 2673.880 1490.550 ;
        RECT 2614.340 1489.725 2614.480 1490.230 ;
        RECT 2614.270 1489.355 2614.550 1489.725 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2614.270 1489.400 2614.550 1489.680 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2614.245 1489.690 2614.575 1489.705 ;
        RECT 2599.460 1489.640 2614.575 1489.690 ;
        RECT 2596.000 1489.390 2614.575 1489.640 ;
        RECT 2596.000 1489.040 2600.000 1489.390 ;
        RECT 2614.245 1489.375 2614.575 1489.390 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2611.950 1214.720 2612.270 1214.780 ;
        RECT 2645.990 1214.720 2646.310 1214.780 ;
        RECT 2611.950 1214.580 2646.310 1214.720 ;
        RECT 2611.950 1214.520 2612.270 1214.580 ;
        RECT 2645.990 1214.520 2646.310 1214.580 ;
        RECT 2645.990 206.960 2646.310 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2645.990 206.820 2901.150 206.960 ;
        RECT 2645.990 206.760 2646.310 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2611.980 1214.520 2612.240 1214.780 ;
        RECT 2646.020 1214.520 2646.280 1214.780 ;
        RECT 2646.020 206.760 2646.280 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2611.970 1215.315 2612.250 1215.685 ;
        RECT 2612.040 1214.810 2612.180 1215.315 ;
        RECT 2611.980 1214.490 2612.240 1214.810 ;
        RECT 2646.020 1214.490 2646.280 1214.810 ;
        RECT 2646.080 207.050 2646.220 1214.490 ;
        RECT 2646.020 206.730 2646.280 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2611.970 1215.360 2612.250 1215.640 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2611.945 1215.650 2612.275 1215.665 ;
        RECT 2599.460 1215.600 2612.275 1215.650 ;
        RECT 2596.000 1215.350 2612.275 1215.600 ;
        RECT 2596.000 1215.000 2600.000 1215.350 ;
        RECT 2611.945 1215.335 2612.275 1215.350 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2680.490 2546.500 2680.810 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 2680.490 2546.360 2901.150 2546.500 ;
        RECT 2680.490 2546.300 2680.810 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
        RECT 2614.250 1531.600 2614.570 1531.660 ;
        RECT 2680.490 1531.600 2680.810 1531.660 ;
        RECT 2614.250 1531.460 2680.810 1531.600 ;
        RECT 2614.250 1531.400 2614.570 1531.460 ;
        RECT 2680.490 1531.400 2680.810 1531.460 ;
      LAYER via ;
        RECT 2680.520 2546.300 2680.780 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
        RECT 2614.280 1531.400 2614.540 1531.660 ;
        RECT 2680.520 1531.400 2680.780 1531.660 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 2680.520 2546.270 2680.780 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 2680.580 1531.690 2680.720 2546.270 ;
        RECT 2614.280 1531.370 2614.540 1531.690 ;
        RECT 2680.520 1531.370 2680.780 1531.690 ;
        RECT 2614.340 1531.205 2614.480 1531.370 ;
        RECT 2614.270 1530.835 2614.550 1531.205 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
        RECT 2614.270 1530.880 2614.550 1531.160 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2614.245 1531.170 2614.575 1531.185 ;
        RECT 2599.460 1531.120 2614.575 1531.170 ;
        RECT 2596.000 1530.870 2614.575 1531.120 ;
        RECT 2596.000 1530.520 2600.000 1530.870 ;
        RECT 2614.245 1530.855 2614.575 1530.870 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2687.390 2781.100 2687.710 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2687.390 2780.960 2901.150 2781.100 ;
        RECT 2687.390 2780.900 2687.710 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
        RECT 2614.250 1566.280 2614.570 1566.340 ;
        RECT 2687.390 1566.280 2687.710 1566.340 ;
        RECT 2614.250 1566.140 2687.710 1566.280 ;
        RECT 2614.250 1566.080 2614.570 1566.140 ;
        RECT 2687.390 1566.080 2687.710 1566.140 ;
      LAYER via ;
        RECT 2687.420 2780.900 2687.680 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
        RECT 2614.280 1566.080 2614.540 1566.340 ;
        RECT 2687.420 1566.080 2687.680 1566.340 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2687.420 2780.870 2687.680 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2687.480 1566.370 2687.620 2780.870 ;
        RECT 2614.280 1566.050 2614.540 1566.370 ;
        RECT 2687.420 1566.050 2687.680 1566.370 ;
        RECT 2614.340 1563.165 2614.480 1566.050 ;
        RECT 2614.270 1562.795 2614.550 1563.165 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2614.270 1562.840 2614.550 1563.120 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2614.245 1563.130 2614.575 1563.145 ;
        RECT 2599.460 1563.080 2614.575 1563.130 ;
        RECT 2596.000 1562.830 2614.575 1563.080 ;
        RECT 2596.000 1562.480 2600.000 1562.830 ;
        RECT 2614.245 1562.815 2614.575 1562.830 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2694.290 3015.700 2694.610 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 2694.290 3015.560 2901.150 3015.700 ;
        RECT 2694.290 3015.500 2694.610 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
        RECT 2614.250 1600.620 2614.570 1600.680 ;
        RECT 2694.290 1600.620 2694.610 1600.680 ;
        RECT 2614.250 1600.480 2694.610 1600.620 ;
        RECT 2614.250 1600.420 2614.570 1600.480 ;
        RECT 2694.290 1600.420 2694.610 1600.480 ;
      LAYER via ;
        RECT 2694.320 3015.500 2694.580 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
        RECT 2614.280 1600.420 2614.540 1600.680 ;
        RECT 2694.320 1600.420 2694.580 1600.680 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 2694.320 3015.470 2694.580 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 2694.380 1600.710 2694.520 3015.470 ;
        RECT 2614.280 1600.390 2614.540 1600.710 ;
        RECT 2694.320 1600.390 2694.580 1600.710 ;
        RECT 2614.340 1594.445 2614.480 1600.390 ;
        RECT 2614.270 1594.075 2614.550 1594.445 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 2614.270 1594.120 2614.550 1594.400 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2614.245 1594.410 2614.575 1594.425 ;
        RECT 2599.460 1594.360 2614.575 1594.410 ;
        RECT 2596.000 1594.110 2614.575 1594.360 ;
        RECT 2596.000 1593.760 2600.000 1594.110 ;
        RECT 2614.245 1594.095 2614.575 1594.110 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2701.190 3250.300 2701.510 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 2701.190 3250.160 2901.150 3250.300 ;
        RECT 2701.190 3250.100 2701.510 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 2614.250 1628.160 2614.570 1628.220 ;
        RECT 2701.190 1628.160 2701.510 1628.220 ;
        RECT 2614.250 1628.020 2701.510 1628.160 ;
        RECT 2614.250 1627.960 2614.570 1628.020 ;
        RECT 2701.190 1627.960 2701.510 1628.020 ;
      LAYER via ;
        RECT 2701.220 3250.100 2701.480 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 2614.280 1627.960 2614.540 1628.220 ;
        RECT 2701.220 1627.960 2701.480 1628.220 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 2701.220 3250.070 2701.480 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 2701.280 1628.250 2701.420 3250.070 ;
        RECT 2614.280 1627.930 2614.540 1628.250 ;
        RECT 2701.220 1627.930 2701.480 1628.250 ;
        RECT 2614.340 1626.405 2614.480 1627.930 ;
        RECT 2614.270 1626.035 2614.550 1626.405 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 2614.270 1626.080 2614.550 1626.360 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2614.245 1626.370 2614.575 1626.385 ;
        RECT 2599.460 1626.320 2614.575 1626.370 ;
        RECT 2596.000 1626.070 2614.575 1626.320 ;
        RECT 2596.000 1625.720 2600.000 1626.070 ;
        RECT 2614.245 1626.055 2614.575 1626.070 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2728.790 3484.900 2729.110 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2728.790 3484.760 2901.150 3484.900 ;
        RECT 2728.790 3484.700 2729.110 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 2614.250 1662.840 2614.570 1662.900 ;
        RECT 2728.790 1662.840 2729.110 1662.900 ;
        RECT 2614.250 1662.700 2729.110 1662.840 ;
        RECT 2614.250 1662.640 2614.570 1662.700 ;
        RECT 2728.790 1662.640 2729.110 1662.700 ;
      LAYER via ;
        RECT 2728.820 3484.700 2729.080 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 2614.280 1662.640 2614.540 1662.900 ;
        RECT 2728.820 1662.640 2729.080 1662.900 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2728.820 3484.670 2729.080 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2728.880 1662.930 2729.020 3484.670 ;
        RECT 2614.280 1662.610 2614.540 1662.930 ;
        RECT 2728.820 1662.610 2729.080 1662.930 ;
        RECT 2614.340 1657.685 2614.480 1662.610 ;
        RECT 2614.270 1657.315 2614.550 1657.685 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 2614.270 1657.360 2614.550 1657.640 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2614.245 1657.650 2614.575 1657.665 ;
        RECT 2599.460 1657.600 2614.575 1657.650 ;
        RECT 2596.000 1657.350 2614.575 1657.600 ;
        RECT 2596.000 1657.000 2600.000 1657.350 ;
        RECT 2614.245 1657.335 2614.575 1657.350 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2614.250 1689.700 2614.570 1689.760 ;
        RECT 2635.870 1689.700 2636.190 1689.760 ;
        RECT 2614.250 1689.560 2636.190 1689.700 ;
        RECT 2614.250 1689.500 2614.570 1689.560 ;
        RECT 2635.870 1689.500 2636.190 1689.560 ;
      LAYER via ;
        RECT 2614.280 1689.500 2614.540 1689.760 ;
        RECT 2635.900 1689.500 2636.160 1689.760 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 1689.790 2636.100 3517.600 ;
        RECT 2614.280 1689.645 2614.540 1689.790 ;
        RECT 2614.270 1689.275 2614.550 1689.645 ;
        RECT 2635.900 1689.470 2636.160 1689.790 ;
      LAYER via2 ;
        RECT 2614.270 1689.320 2614.550 1689.600 ;
      LAYER met3 ;
        RECT 2614.245 1689.610 2614.575 1689.625 ;
        RECT 2599.460 1689.560 2614.575 1689.610 ;
        RECT 2596.000 1689.310 2614.575 1689.560 ;
        RECT 2596.000 1688.960 2600.000 1689.310 ;
        RECT 2614.245 1689.295 2614.575 1689.310 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2311.570 3500.540 2311.890 3500.600 ;
        RECT 2318.010 3500.540 2318.330 3500.600 ;
        RECT 2311.570 3500.400 2318.330 3500.540 ;
        RECT 2311.570 3500.340 2311.890 3500.400 ;
        RECT 2318.010 3500.340 2318.330 3500.400 ;
        RECT 2318.010 3053.780 2318.330 3053.840 ;
        RECT 2597.690 3053.780 2598.010 3053.840 ;
        RECT 2318.010 3053.640 2598.010 3053.780 ;
        RECT 2318.010 3053.580 2318.330 3053.640 ;
        RECT 2597.690 3053.580 2598.010 3053.640 ;
      LAYER via ;
        RECT 2311.600 3500.340 2311.860 3500.600 ;
        RECT 2318.040 3500.340 2318.300 3500.600 ;
        RECT 2318.040 3053.580 2318.300 3053.840 ;
        RECT 2597.720 3053.580 2597.980 3053.840 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3500.630 2311.800 3517.600 ;
        RECT 2311.600 3500.310 2311.860 3500.630 ;
        RECT 2318.040 3500.310 2318.300 3500.630 ;
        RECT 2318.100 3053.870 2318.240 3500.310 ;
        RECT 2318.040 3053.550 2318.300 3053.870 ;
        RECT 2597.720 3053.550 2597.980 3053.870 ;
        RECT 2597.780 1722.965 2597.920 3053.550 ;
        RECT 2597.710 1722.595 2597.990 1722.965 ;
      LAYER via2 ;
        RECT 2597.710 1722.640 2597.990 1722.920 ;
      LAYER met3 ;
        RECT 2597.685 1722.930 2598.015 1722.945 ;
        RECT 2597.470 1722.615 2598.015 1722.930 ;
        RECT 2597.470 1720.840 2597.770 1722.615 ;
        RECT 2596.000 1720.240 2600.000 1720.840 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1987.270 3499.860 1987.590 3499.920 ;
        RECT 1993.710 3499.860 1994.030 3499.920 ;
        RECT 1987.270 3499.720 1994.030 3499.860 ;
        RECT 1987.270 3499.660 1987.590 3499.720 ;
        RECT 1993.710 3499.660 1994.030 3499.720 ;
        RECT 1993.710 2404.720 1994.030 2404.780 ;
        RECT 1993.710 2404.580 2587.340 2404.720 ;
        RECT 1993.710 2404.520 1994.030 2404.580 ;
        RECT 2587.200 2404.040 2587.340 2404.580 ;
        RECT 2599.530 2404.040 2599.850 2404.100 ;
        RECT 2587.200 2403.900 2599.850 2404.040 ;
        RECT 2599.530 2403.840 2599.850 2403.900 ;
        RECT 2599.530 2396.900 2599.850 2396.960 ;
        RECT 2604.130 2396.900 2604.450 2396.960 ;
        RECT 2599.530 2396.760 2604.450 2396.900 ;
        RECT 2599.530 2396.700 2599.850 2396.760 ;
        RECT 2604.130 2396.700 2604.450 2396.760 ;
        RECT 2600.450 2380.580 2600.770 2380.640 ;
        RECT 2604.130 2380.580 2604.450 2380.640 ;
        RECT 2600.450 2380.440 2604.450 2380.580 ;
        RECT 2600.450 2380.380 2600.770 2380.440 ;
        RECT 2604.130 2380.380 2604.450 2380.440 ;
        RECT 2599.070 2342.500 2599.390 2342.560 ;
        RECT 2600.450 2342.500 2600.770 2342.560 ;
        RECT 2599.070 2342.360 2600.770 2342.500 ;
        RECT 2599.070 2342.300 2599.390 2342.360 ;
        RECT 2600.450 2342.300 2600.770 2342.360 ;
      LAYER via ;
        RECT 1987.300 3499.660 1987.560 3499.920 ;
        RECT 1993.740 3499.660 1994.000 3499.920 ;
        RECT 1993.740 2404.520 1994.000 2404.780 ;
        RECT 2599.560 2403.840 2599.820 2404.100 ;
        RECT 2599.560 2396.700 2599.820 2396.960 ;
        RECT 2604.160 2396.700 2604.420 2396.960 ;
        RECT 2600.480 2380.380 2600.740 2380.640 ;
        RECT 2604.160 2380.380 2604.420 2380.640 ;
        RECT 2599.100 2342.300 2599.360 2342.560 ;
        RECT 2600.480 2342.300 2600.740 2342.560 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3499.950 1987.500 3517.600 ;
        RECT 1987.300 3499.630 1987.560 3499.950 ;
        RECT 1993.740 3499.630 1994.000 3499.950 ;
        RECT 1993.800 2404.810 1993.940 3499.630 ;
        RECT 1993.740 2404.490 1994.000 2404.810 ;
        RECT 2599.560 2403.810 2599.820 2404.130 ;
        RECT 2599.620 2396.990 2599.760 2403.810 ;
        RECT 2599.560 2396.670 2599.820 2396.990 ;
        RECT 2604.160 2396.670 2604.420 2396.990 ;
        RECT 2604.220 2380.670 2604.360 2396.670 ;
        RECT 2600.480 2380.350 2600.740 2380.670 ;
        RECT 2604.160 2380.350 2604.420 2380.670 ;
        RECT 2600.540 2342.590 2600.680 2380.350 ;
        RECT 2599.100 2342.270 2599.360 2342.590 ;
        RECT 2600.480 2342.270 2600.740 2342.590 ;
        RECT 2599.160 1755.605 2599.300 2342.270 ;
        RECT 2599.090 1755.235 2599.370 1755.605 ;
      LAYER via2 ;
        RECT 2599.090 1755.280 2599.370 1755.560 ;
      LAYER met3 ;
        RECT 2599.065 1755.570 2599.395 1755.585 ;
        RECT 2599.065 1755.255 2599.610 1755.570 ;
        RECT 2599.310 1752.800 2599.610 1755.255 ;
        RECT 2596.000 1752.200 2600.000 1752.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 3503.600 1662.830 3503.660 ;
        RECT 2595.390 3503.600 2595.710 3503.660 ;
        RECT 1662.510 3503.460 2595.710 3503.600 ;
        RECT 1662.510 3503.400 1662.830 3503.460 ;
        RECT 2595.390 3503.400 2595.710 3503.460 ;
      LAYER via ;
        RECT 1662.540 3503.400 1662.800 3503.660 ;
        RECT 2595.420 3503.400 2595.680 3503.660 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3503.690 1662.740 3517.600 ;
        RECT 1662.540 3503.370 1662.800 3503.690 ;
        RECT 2595.420 3503.370 2595.680 3503.690 ;
        RECT 2595.480 1786.770 2595.620 3503.370 ;
        RECT 2596.790 1786.770 2597.070 1786.885 ;
        RECT 2595.480 1786.630 2597.070 1786.770 ;
        RECT 2596.790 1786.515 2597.070 1786.630 ;
      LAYER via2 ;
        RECT 2596.790 1786.560 2597.070 1786.840 ;
      LAYER met3 ;
        RECT 2596.765 1786.850 2597.095 1786.865 ;
        RECT 2596.550 1786.535 2597.095 1786.850 ;
        RECT 2596.550 1784.080 2596.850 1786.535 ;
        RECT 2596.000 1783.480 2600.000 1784.080 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3502.920 1338.530 3502.980 ;
        RECT 2595.850 3502.920 2596.170 3502.980 ;
        RECT 1338.210 3502.780 2596.170 3502.920 ;
        RECT 1338.210 3502.720 1338.530 3502.780 ;
        RECT 2595.850 3502.720 2596.170 3502.780 ;
      LAYER via ;
        RECT 1338.240 3502.720 1338.500 3502.980 ;
        RECT 2595.880 3502.720 2596.140 3502.980 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3503.010 1338.440 3517.600 ;
        RECT 1338.240 3502.690 1338.500 3503.010 ;
        RECT 2595.880 3502.690 2596.140 3503.010 ;
        RECT 2595.940 1818.050 2596.080 3502.690 ;
        RECT 2596.790 1818.050 2597.070 1818.165 ;
        RECT 2595.940 1817.910 2597.070 1818.050 ;
        RECT 2596.790 1817.795 2597.070 1817.910 ;
      LAYER via2 ;
        RECT 2596.790 1817.840 2597.070 1818.120 ;
      LAYER met3 ;
        RECT 2596.765 1818.130 2597.095 1818.145 ;
        RECT 2596.550 1817.815 2597.095 1818.130 ;
        RECT 2596.550 1815.360 2596.850 1817.815 ;
        RECT 2596.000 1814.760 2600.000 1815.360 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2608.270 1242.260 2608.590 1242.320 ;
        RECT 2659.790 1242.260 2660.110 1242.320 ;
        RECT 2608.270 1242.120 2660.110 1242.260 ;
        RECT 2608.270 1242.060 2608.590 1242.120 ;
        RECT 2659.790 1242.060 2660.110 1242.120 ;
        RECT 2659.790 441.560 2660.110 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2659.790 441.420 2901.150 441.560 ;
        RECT 2659.790 441.360 2660.110 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2608.300 1242.060 2608.560 1242.320 ;
        RECT 2659.820 1242.060 2660.080 1242.320 ;
        RECT 2659.820 441.360 2660.080 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2608.290 1246.595 2608.570 1246.965 ;
        RECT 2608.360 1242.350 2608.500 1246.595 ;
        RECT 2608.300 1242.030 2608.560 1242.350 ;
        RECT 2659.820 1242.030 2660.080 1242.350 ;
        RECT 2659.880 441.650 2660.020 1242.030 ;
        RECT 2659.820 441.330 2660.080 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2608.290 1246.640 2608.570 1246.920 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2608.265 1246.930 2608.595 1246.945 ;
        RECT 2599.460 1246.880 2608.595 1246.930 ;
        RECT 2596.000 1246.630 2608.595 1246.880 ;
        RECT 2596.000 1246.280 2600.000 1246.630 ;
        RECT 2608.265 1246.615 2608.595 1246.630 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3502.240 1014.230 3502.300 ;
        RECT 2596.310 3502.240 2596.630 3502.300 ;
        RECT 1013.910 3502.100 2596.630 3502.240 ;
        RECT 1013.910 3502.040 1014.230 3502.100 ;
        RECT 2596.310 3502.040 2596.630 3502.100 ;
      LAYER via ;
        RECT 1013.940 3502.040 1014.200 3502.300 ;
        RECT 2596.340 3502.040 2596.600 3502.300 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3502.330 1014.140 3517.600 ;
        RECT 1013.940 3502.010 1014.200 3502.330 ;
        RECT 2596.340 3502.010 2596.600 3502.330 ;
        RECT 2596.400 1848.650 2596.540 3502.010 ;
        RECT 2596.790 1848.650 2597.070 1848.765 ;
        RECT 2596.400 1848.510 2597.070 1848.650 ;
        RECT 2596.790 1848.395 2597.070 1848.510 ;
      LAYER via2 ;
        RECT 2596.790 1848.440 2597.070 1848.720 ;
      LAYER met3 ;
        RECT 2596.765 1848.730 2597.095 1848.745 ;
        RECT 2596.550 1848.415 2597.095 1848.730 ;
        RECT 2596.550 1847.320 2596.850 1848.415 ;
        RECT 2596.000 1846.720 2600.000 1847.320 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3501.560 689.470 3501.620 ;
        RECT 2597.230 3501.560 2597.550 3501.620 ;
        RECT 689.150 3501.420 2597.550 3501.560 ;
        RECT 689.150 3501.360 689.470 3501.420 ;
        RECT 2597.230 3501.360 2597.550 3501.420 ;
      LAYER via ;
        RECT 689.180 3501.360 689.440 3501.620 ;
        RECT 2597.260 3501.360 2597.520 3501.620 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3501.650 689.380 3517.600 ;
        RECT 689.180 3501.330 689.440 3501.650 ;
        RECT 2597.260 3501.330 2597.520 3501.650 ;
        RECT 2597.320 1881.405 2597.460 3501.330 ;
        RECT 2597.250 1881.035 2597.530 1881.405 ;
      LAYER via2 ;
        RECT 2597.250 1881.080 2597.530 1881.360 ;
      LAYER met3 ;
        RECT 2597.225 1881.370 2597.555 1881.385 ;
        RECT 2597.225 1881.055 2597.770 1881.370 ;
        RECT 2597.470 1878.600 2597.770 1881.055 ;
        RECT 2596.000 1878.000 2600.000 1878.600 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3503.205 365.080 3517.600 ;
        RECT 364.870 3502.835 365.150 3503.205 ;
      LAYER via2 ;
        RECT 364.870 3502.880 365.150 3503.160 ;
      LAYER met3 ;
        RECT 364.845 3503.170 365.175 3503.185 ;
        RECT 2594.670 3503.170 2595.050 3503.180 ;
        RECT 364.845 3502.870 2595.050 3503.170 ;
        RECT 364.845 3502.855 365.175 3502.870 ;
        RECT 2594.670 3502.860 2595.050 3502.870 ;
        RECT 2596.510 1910.980 2596.890 1911.300 ;
        RECT 2596.550 1910.560 2596.850 1910.980 ;
        RECT 2596.000 1909.960 2600.000 1910.560 ;
      LAYER via3 ;
        RECT 2594.700 3502.860 2595.020 3503.180 ;
        RECT 2596.540 1910.980 2596.860 1911.300 ;
      LAYER met4 ;
        RECT 2594.695 3502.855 2595.025 3503.185 ;
        RECT 2594.710 1940.530 2595.010 3502.855 ;
        RECT 2594.710 1940.230 2596.850 1940.530 ;
        RECT 2596.550 1911.305 2596.850 1940.230 ;
        RECT 2596.535 1910.975 2596.865 1911.305 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 2595.590 3501.810 2595.970 3501.820 ;
        RECT 40.545 3501.510 2595.970 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 2595.590 3501.500 2595.970 3501.510 ;
        RECT 2596.510 1942.940 2596.890 1943.260 ;
        RECT 2596.550 1941.840 2596.850 1942.940 ;
        RECT 2596.000 1941.240 2600.000 1941.840 ;
      LAYER via3 ;
        RECT 2595.620 3501.500 2595.940 3501.820 ;
        RECT 2596.540 1942.940 2596.860 1943.260 ;
      LAYER met4 ;
        RECT 2595.615 3501.495 2595.945 3501.825 ;
        RECT 2595.630 1943.250 2595.930 3501.495 ;
        RECT 2596.535 1943.250 2596.865 1943.265 ;
        RECT 2595.630 1942.950 2596.865 1943.250 ;
        RECT 2596.535 1942.935 2596.865 1942.950 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.650 3267.555 16.930 3267.925 ;
        RECT 16.720 3264.525 16.860 3267.555 ;
        RECT 16.650 3264.155 16.930 3264.525 ;
      LAYER via2 ;
        RECT 16.650 3267.600 16.930 3267.880 ;
        RECT 16.650 3264.200 16.930 3264.480 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 16.625 3267.890 16.955 3267.905 ;
        RECT -4.800 3267.590 16.955 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 16.625 3267.575 16.955 3267.590 ;
        RECT 16.625 3264.490 16.955 3264.505 ;
        RECT 2597.430 3264.490 2597.810 3264.500 ;
        RECT 16.625 3264.190 2597.810 3264.490 ;
        RECT 16.625 3264.175 16.955 3264.190 ;
        RECT 2597.430 3264.180 2597.810 3264.190 ;
        RECT 2597.430 1976.260 2597.810 1976.580 ;
        RECT 2597.470 1973.800 2597.770 1976.260 ;
        RECT 2596.000 1973.200 2600.000 1973.800 ;
      LAYER via3 ;
        RECT 2597.460 3264.180 2597.780 3264.500 ;
        RECT 2597.460 1976.260 2597.780 1976.580 ;
      LAYER met4 ;
        RECT 2597.455 3264.175 2597.785 3264.505 ;
        RECT 2597.470 1976.585 2597.770 3264.175 ;
        RECT 2597.455 1976.255 2597.785 1976.585 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2397.920 17.870 2397.980 ;
        RECT 2612.870 2397.920 2613.190 2397.980 ;
        RECT 17.550 2397.780 2613.190 2397.920 ;
        RECT 17.550 2397.720 17.870 2397.780 ;
        RECT 2612.870 2397.720 2613.190 2397.780 ;
      LAYER via ;
        RECT 17.580 2397.720 17.840 2397.980 ;
        RECT 2612.900 2397.720 2613.160 2397.980 ;
      LAYER met2 ;
        RECT 17.570 2979.915 17.850 2980.285 ;
        RECT 17.640 2398.010 17.780 2979.915 ;
        RECT 17.580 2397.690 17.840 2398.010 ;
        RECT 2612.900 2397.690 2613.160 2398.010 ;
        RECT 2612.960 2005.165 2613.100 2397.690 ;
        RECT 2612.890 2004.795 2613.170 2005.165 ;
      LAYER via2 ;
        RECT 17.570 2979.960 17.850 2980.240 ;
        RECT 2612.890 2004.840 2613.170 2005.120 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 17.545 2980.250 17.875 2980.265 ;
        RECT -4.800 2979.950 17.875 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 17.545 2979.935 17.875 2979.950 ;
        RECT 2612.865 2005.130 2613.195 2005.145 ;
        RECT 2599.460 2005.080 2613.195 2005.130 ;
        RECT 2596.000 2004.830 2613.195 2005.080 ;
        RECT 2596.000 2004.480 2600.000 2004.830 ;
        RECT 2612.865 2004.815 2613.195 2004.830 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 2398.260 19.250 2398.320 ;
        RECT 2613.330 2398.260 2613.650 2398.320 ;
        RECT 18.930 2398.120 2613.650 2398.260 ;
        RECT 18.930 2398.060 19.250 2398.120 ;
        RECT 2613.330 2398.060 2613.650 2398.120 ;
      LAYER via ;
        RECT 18.960 2398.060 19.220 2398.320 ;
        RECT 2613.360 2398.060 2613.620 2398.320 ;
      LAYER met2 ;
        RECT 18.950 2692.955 19.230 2693.325 ;
        RECT 19.020 2398.350 19.160 2692.955 ;
        RECT 18.960 2398.030 19.220 2398.350 ;
        RECT 2613.360 2398.030 2613.620 2398.350 ;
        RECT 2613.420 2037.125 2613.560 2398.030 ;
        RECT 2613.350 2036.755 2613.630 2037.125 ;
      LAYER via2 ;
        RECT 18.950 2693.000 19.230 2693.280 ;
        RECT 2613.350 2036.800 2613.630 2037.080 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 18.925 2693.290 19.255 2693.305 ;
        RECT -4.800 2692.990 19.255 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 18.925 2692.975 19.255 2692.990 ;
        RECT 2613.325 2037.090 2613.655 2037.105 ;
        RECT 2599.460 2037.040 2613.655 2037.090 ;
        RECT 2596.000 2036.790 2613.655 2037.040 ;
        RECT 2596.000 2036.440 2600.000 2036.790 ;
        RECT 2613.325 2036.775 2613.655 2036.790 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 2401.320 15.110 2401.380 ;
        RECT 2599.070 2401.320 2599.390 2401.380 ;
        RECT 14.790 2401.180 2599.390 2401.320 ;
        RECT 14.790 2401.120 15.110 2401.180 ;
        RECT 2599.070 2401.120 2599.390 2401.180 ;
        RECT 2599.070 2343.180 2599.390 2343.240 ;
        RECT 2599.070 2343.040 2601.140 2343.180 ;
        RECT 2599.070 2342.980 2599.390 2343.040 ;
        RECT 2600.450 2341.820 2600.770 2341.880 ;
        RECT 2601.000 2341.820 2601.140 2343.040 ;
        RECT 2600.450 2341.680 2601.140 2341.820 ;
        RECT 2600.450 2341.620 2600.770 2341.680 ;
      LAYER via ;
        RECT 14.820 2401.120 15.080 2401.380 ;
        RECT 2599.100 2401.120 2599.360 2401.380 ;
        RECT 2599.100 2342.980 2599.360 2343.240 ;
        RECT 2600.480 2341.620 2600.740 2341.880 ;
      LAYER met2 ;
        RECT 14.810 2405.315 15.090 2405.685 ;
        RECT 14.880 2401.410 15.020 2405.315 ;
        RECT 14.820 2401.090 15.080 2401.410 ;
        RECT 2599.100 2401.090 2599.360 2401.410 ;
        RECT 2599.160 2343.270 2599.300 2401.090 ;
        RECT 2599.100 2342.950 2599.360 2343.270 ;
        RECT 2600.480 2341.590 2600.740 2341.910 ;
        RECT 2600.540 2068.405 2600.680 2341.590 ;
        RECT 2600.470 2068.035 2600.750 2068.405 ;
      LAYER via2 ;
        RECT 14.810 2405.360 15.090 2405.640 ;
        RECT 2600.470 2068.080 2600.750 2068.360 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 14.785 2405.650 15.115 2405.665 ;
        RECT -4.800 2405.350 15.115 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 14.785 2405.335 15.115 2405.350 ;
        RECT 2600.445 2068.370 2600.775 2068.385 ;
        RECT 2599.460 2068.320 2600.775 2068.370 ;
        RECT 2596.000 2068.070 2600.775 2068.320 ;
        RECT 2596.000 2067.720 2600.000 2068.070 ;
        RECT 2600.445 2068.055 2600.775 2068.070 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1396.630 2394.860 1396.950 2394.920 ;
        RECT 2615.170 2394.860 2615.490 2394.920 ;
        RECT 1396.630 2394.720 2615.490 2394.860 ;
        RECT 1396.630 2394.660 1396.950 2394.720 ;
        RECT 2615.170 2394.660 2615.490 2394.720 ;
        RECT 16.170 2125.240 16.490 2125.300 ;
        RECT 1396.630 2125.240 1396.950 2125.300 ;
        RECT 16.170 2125.100 1396.950 2125.240 ;
        RECT 16.170 2125.040 16.490 2125.100 ;
        RECT 1396.630 2125.040 1396.950 2125.100 ;
      LAYER via ;
        RECT 1396.660 2394.660 1396.920 2394.920 ;
        RECT 2615.200 2394.660 2615.460 2394.920 ;
        RECT 16.200 2125.040 16.460 2125.300 ;
        RECT 1396.660 2125.040 1396.920 2125.300 ;
      LAYER met2 ;
        RECT 1396.660 2394.630 1396.920 2394.950 ;
        RECT 2615.200 2394.630 2615.460 2394.950 ;
        RECT 1396.720 2125.330 1396.860 2394.630 ;
        RECT 16.200 2125.010 16.460 2125.330 ;
        RECT 1396.660 2125.010 1396.920 2125.330 ;
        RECT 16.260 2118.725 16.400 2125.010 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
        RECT 2615.260 2100.365 2615.400 2394.630 ;
        RECT 2615.190 2099.995 2615.470 2100.365 ;
      LAYER via2 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
        RECT 2615.190 2100.040 2615.470 2100.320 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
        RECT 2615.165 2100.330 2615.495 2100.345 ;
        RECT 2599.460 2100.280 2615.495 2100.330 ;
        RECT 2596.000 2100.030 2615.495 2100.280 ;
        RECT 2596.000 2099.680 2600.000 2100.030 ;
        RECT 2615.165 2100.015 2615.495 2100.030 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1399.390 2395.200 1399.710 2395.260 ;
        RECT 2616.090 2395.200 2616.410 2395.260 ;
        RECT 1399.390 2395.060 2616.410 2395.200 ;
        RECT 1399.390 2395.000 1399.710 2395.060 ;
        RECT 2616.090 2395.000 2616.410 2395.060 ;
        RECT 2608.270 2131.700 2608.590 2131.760 ;
        RECT 2616.090 2131.700 2616.410 2131.760 ;
        RECT 2608.270 2131.560 2616.410 2131.700 ;
        RECT 2608.270 2131.500 2608.590 2131.560 ;
        RECT 2616.090 2131.500 2616.410 2131.560 ;
        RECT 17.550 1835.220 17.870 1835.280 ;
        RECT 1399.390 1835.220 1399.710 1835.280 ;
        RECT 17.550 1835.080 1399.710 1835.220 ;
        RECT 17.550 1835.020 17.870 1835.080 ;
        RECT 1399.390 1835.020 1399.710 1835.080 ;
      LAYER via ;
        RECT 1399.420 2395.000 1399.680 2395.260 ;
        RECT 2616.120 2395.000 2616.380 2395.260 ;
        RECT 2608.300 2131.500 2608.560 2131.760 ;
        RECT 2616.120 2131.500 2616.380 2131.760 ;
        RECT 17.580 1835.020 17.840 1835.280 ;
        RECT 1399.420 1835.020 1399.680 1835.280 ;
      LAYER met2 ;
        RECT 1399.420 2394.970 1399.680 2395.290 ;
        RECT 2616.120 2394.970 2616.380 2395.290 ;
        RECT 1399.480 1835.310 1399.620 2394.970 ;
        RECT 2616.180 2131.790 2616.320 2394.970 ;
        RECT 2608.300 2131.645 2608.560 2131.790 ;
        RECT 2608.290 2131.275 2608.570 2131.645 ;
        RECT 2616.120 2131.470 2616.380 2131.790 ;
        RECT 17.580 1834.990 17.840 1835.310 ;
        RECT 1399.420 1834.990 1399.680 1835.310 ;
        RECT 17.640 1831.085 17.780 1834.990 ;
        RECT 17.570 1830.715 17.850 1831.085 ;
      LAYER via2 ;
        RECT 2608.290 2131.320 2608.570 2131.600 ;
        RECT 17.570 1830.760 17.850 1831.040 ;
      LAYER met3 ;
        RECT 2608.265 2131.610 2608.595 2131.625 ;
        RECT 2599.460 2131.560 2608.595 2131.610 ;
        RECT 2596.000 2131.310 2608.595 2131.560 ;
        RECT 2596.000 2130.960 2600.000 2131.310 ;
        RECT 2608.265 2131.295 2608.595 2131.310 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 17.545 1831.050 17.875 1831.065 ;
        RECT -4.800 1830.750 17.875 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 17.545 1830.735 17.875 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2613.790 676.160 2614.110 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2613.790 676.020 2901.150 676.160 ;
        RECT 2613.790 675.960 2614.110 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2613.820 675.960 2614.080 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2613.810 1278.555 2614.090 1278.925 ;
        RECT 2613.880 676.250 2614.020 1278.555 ;
        RECT 2613.820 675.930 2614.080 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2613.810 1278.600 2614.090 1278.880 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2613.785 1278.890 2614.115 1278.905 ;
        RECT 2599.460 1278.840 2614.115 1278.890 ;
        RECT 2596.000 1278.590 2614.115 1278.840 ;
        RECT 2596.000 1278.240 2600.000 1278.590 ;
        RECT 2613.785 1278.575 2614.115 1278.590 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1398.010 2397.240 1398.330 2397.300 ;
        RECT 2596.770 2397.240 2597.090 2397.300 ;
        RECT 1398.010 2397.100 2597.090 2397.240 ;
        RECT 1398.010 2397.040 1398.330 2397.100 ;
        RECT 2596.770 2397.040 2597.090 2397.100 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 1398.010 1545.540 1398.330 1545.600 ;
        RECT 16.630 1545.400 1398.330 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 1398.010 1545.340 1398.330 1545.400 ;
      LAYER via ;
        RECT 1398.040 2397.040 1398.300 2397.300 ;
        RECT 2596.800 2397.040 2597.060 2397.300 ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 1398.040 1545.340 1398.300 1545.600 ;
      LAYER met2 ;
        RECT 1398.040 2397.010 1398.300 2397.330 ;
        RECT 2596.800 2397.010 2597.060 2397.330 ;
        RECT 1398.100 1545.630 1398.240 2397.010 ;
        RECT 2596.860 2380.525 2597.000 2397.010 ;
        RECT 2596.790 2380.155 2597.070 2380.525 ;
        RECT 2596.790 2284.275 2597.070 2284.645 ;
        RECT 2596.860 2256.085 2597.000 2284.275 ;
        RECT 2596.790 2255.715 2597.070 2256.085 ;
        RECT 2596.790 2208.115 2597.070 2208.485 ;
        RECT 2596.860 2165.645 2597.000 2208.115 ;
        RECT 2596.790 2165.275 2597.070 2165.645 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 1398.040 1545.310 1398.300 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 2596.790 2380.200 2597.070 2380.480 ;
        RECT 2596.790 2284.320 2597.070 2284.600 ;
        RECT 2596.790 2255.760 2597.070 2256.040 ;
        RECT 2596.790 2208.160 2597.070 2208.440 ;
        RECT 2596.790 2165.320 2597.070 2165.600 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 2596.765 2380.490 2597.095 2380.505 ;
        RECT 2599.270 2380.490 2599.650 2380.500 ;
        RECT 2596.765 2380.190 2599.650 2380.490 ;
        RECT 2596.765 2380.175 2597.095 2380.190 ;
        RECT 2599.270 2380.180 2599.650 2380.190 ;
        RECT 2596.765 2284.610 2597.095 2284.625 ;
        RECT 2600.190 2284.610 2600.570 2284.620 ;
        RECT 2596.765 2284.310 2600.570 2284.610 ;
        RECT 2596.765 2284.295 2597.095 2284.310 ;
        RECT 2600.190 2284.300 2600.570 2284.310 ;
        RECT 2596.765 2256.050 2597.095 2256.065 ;
        RECT 2599.270 2256.050 2599.650 2256.060 ;
        RECT 2596.765 2255.750 2599.650 2256.050 ;
        RECT 2596.765 2255.735 2597.095 2255.750 ;
        RECT 2599.270 2255.740 2599.650 2255.750 ;
        RECT 2596.765 2208.450 2597.095 2208.465 ;
        RECT 2599.270 2208.450 2599.650 2208.460 ;
        RECT 2596.765 2208.150 2599.650 2208.450 ;
        RECT 2596.765 2208.135 2597.095 2208.150 ;
        RECT 2599.270 2208.140 2599.650 2208.150 ;
        RECT 2596.765 2165.610 2597.095 2165.625 ;
        RECT 2596.550 2165.295 2597.095 2165.610 ;
        RECT 2596.550 2162.840 2596.850 2165.295 ;
        RECT 2596.000 2162.240 2600.000 2162.840 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
      LAYER via3 ;
        RECT 2599.300 2380.180 2599.620 2380.500 ;
        RECT 2600.220 2284.300 2600.540 2284.620 ;
        RECT 2599.300 2255.740 2599.620 2256.060 ;
        RECT 2599.300 2208.140 2599.620 2208.460 ;
      LAYER met4 ;
        RECT 2599.295 2380.175 2599.625 2380.505 ;
        RECT 2599.310 2368.250 2599.610 2380.175 ;
        RECT 2599.310 2367.950 2600.530 2368.250 ;
        RECT 2600.230 2284.625 2600.530 2367.950 ;
        RECT 2600.215 2284.295 2600.545 2284.625 ;
        RECT 2599.295 2255.735 2599.625 2256.065 ;
        RECT 2599.310 2208.465 2599.610 2255.735 ;
        RECT 2599.295 2208.135 2599.625 2208.465 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2611.950 1215.880 2612.270 1216.140 ;
        RECT 2612.040 1215.060 2612.180 1215.880 ;
        RECT 2611.580 1214.920 2612.180 1215.060 ;
        RECT 2611.580 1214.040 2611.720 1214.920 ;
        RECT 2611.950 1214.040 2612.270 1214.100 ;
        RECT 2611.580 1213.900 2612.270 1214.040 ;
        RECT 2611.950 1213.840 2612.270 1213.900 ;
        RECT 17.550 1204.180 17.870 1204.240 ;
        RECT 2611.950 1204.180 2612.270 1204.240 ;
        RECT 17.550 1204.040 2612.270 1204.180 ;
        RECT 17.550 1203.980 17.870 1204.040 ;
        RECT 2611.950 1203.980 2612.270 1204.040 ;
      LAYER via ;
        RECT 2611.980 1215.880 2612.240 1216.140 ;
        RECT 2611.980 1213.840 2612.240 1214.100 ;
        RECT 17.580 1203.980 17.840 1204.240 ;
        RECT 2611.980 1203.980 2612.240 1204.240 ;
      LAYER met2 ;
        RECT 2611.970 2194.515 2612.250 2194.885 ;
        RECT 17.570 1328.195 17.850 1328.565 ;
        RECT 17.640 1204.270 17.780 1328.195 ;
        RECT 2612.040 1216.170 2612.180 2194.515 ;
        RECT 2611.980 1215.850 2612.240 1216.170 ;
        RECT 2611.980 1213.810 2612.240 1214.130 ;
        RECT 2612.040 1204.270 2612.180 1213.810 ;
        RECT 17.580 1203.950 17.840 1204.270 ;
        RECT 2611.980 1203.950 2612.240 1204.270 ;
      LAYER via2 ;
        RECT 2611.970 2194.560 2612.250 2194.840 ;
        RECT 17.570 1328.240 17.850 1328.520 ;
      LAYER met3 ;
        RECT 2611.945 2194.850 2612.275 2194.865 ;
        RECT 2599.460 2194.800 2612.275 2194.850 ;
        RECT 2596.000 2194.550 2612.275 2194.800 ;
        RECT 2596.000 2194.200 2600.000 2194.550 ;
        RECT 2611.945 2194.535 2612.275 2194.550 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 17.545 1328.530 17.875 1328.545 ;
        RECT -4.800 1328.230 17.875 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 17.545 1328.215 17.875 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 2611.490 1117.820 2611.810 1117.880 ;
        RECT 15.710 1117.680 2611.810 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 2611.490 1117.620 2611.810 1117.680 ;
      LAYER via ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 2611.520 1117.620 2611.780 1117.880 ;
      LAYER met2 ;
        RECT 2611.510 2225.795 2611.790 2226.165 ;
        RECT 2611.580 1117.910 2611.720 2225.795 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 2611.520 1117.590 2611.780 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 2611.510 2225.840 2611.790 2226.120 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT 2611.485 2226.130 2611.815 2226.145 ;
        RECT 2599.460 2226.080 2611.815 2226.130 ;
        RECT 2596.000 2225.830 2611.815 2226.080 ;
        RECT 2596.000 2225.480 2600.000 2225.830 ;
        RECT 2611.485 2225.815 2611.815 2225.830 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.390 1003.920 19.710 1003.980 ;
        RECT 2610.570 1003.920 2610.890 1003.980 ;
        RECT 19.390 1003.780 2610.890 1003.920 ;
        RECT 19.390 1003.720 19.710 1003.780 ;
        RECT 2610.570 1003.720 2610.890 1003.780 ;
      LAYER via ;
        RECT 19.420 1003.720 19.680 1003.980 ;
        RECT 2610.600 1003.720 2610.860 1003.980 ;
      LAYER met2 ;
        RECT 2610.590 2257.755 2610.870 2258.125 ;
        RECT 2610.660 1004.010 2610.800 2257.755 ;
        RECT 19.420 1003.690 19.680 1004.010 ;
        RECT 2610.600 1003.690 2610.860 1004.010 ;
        RECT 19.480 897.445 19.620 1003.690 ;
        RECT 19.410 897.075 19.690 897.445 ;
      LAYER via2 ;
        RECT 2610.590 2257.800 2610.870 2258.080 ;
        RECT 19.410 897.120 19.690 897.400 ;
      LAYER met3 ;
        RECT 2610.565 2258.090 2610.895 2258.105 ;
        RECT 2599.460 2258.040 2610.895 2258.090 ;
        RECT 2596.000 2257.790 2610.895 2258.040 ;
        RECT 2596.000 2257.440 2600.000 2257.790 ;
        RECT 2610.565 2257.775 2610.895 2257.790 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 19.385 897.410 19.715 897.425 ;
        RECT -4.800 897.110 19.715 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 19.385 897.095 19.715 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 1004.260 18.330 1004.320 ;
        RECT 2609.190 1004.260 2609.510 1004.320 ;
        RECT 18.010 1004.120 2609.510 1004.260 ;
        RECT 18.010 1004.060 18.330 1004.120 ;
        RECT 2609.190 1004.060 2609.510 1004.120 ;
      LAYER via ;
        RECT 18.040 1004.060 18.300 1004.320 ;
        RECT 2609.220 1004.060 2609.480 1004.320 ;
      LAYER met2 ;
        RECT 2609.210 2289.035 2609.490 2289.405 ;
        RECT 2609.280 1004.350 2609.420 2289.035 ;
        RECT 18.040 1004.030 18.300 1004.350 ;
        RECT 2609.220 1004.030 2609.480 1004.350 ;
        RECT 18.100 681.885 18.240 1004.030 ;
        RECT 18.030 681.515 18.310 681.885 ;
      LAYER via2 ;
        RECT 2609.210 2289.080 2609.490 2289.360 ;
        RECT 18.030 681.560 18.310 681.840 ;
      LAYER met3 ;
        RECT 2609.185 2289.370 2609.515 2289.385 ;
        RECT 2599.460 2289.320 2609.515 2289.370 ;
        RECT 2596.000 2289.070 2609.515 2289.320 ;
        RECT 2596.000 2288.720 2600.000 2289.070 ;
        RECT 2609.185 2289.055 2609.515 2289.070 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 18.005 681.850 18.335 681.865 ;
        RECT -4.800 681.550 18.335 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 18.005 681.535 18.335 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2612.150 2321.330 2612.530 2321.340 ;
        RECT 2599.460 2321.280 2612.530 2321.330 ;
        RECT 2596.000 2321.030 2612.530 2321.280 ;
        RECT 2596.000 2320.680 2600.000 2321.030 ;
        RECT 2612.150 2321.020 2612.530 2321.030 ;
        RECT 2612.150 469.010 2612.530 469.020 ;
        RECT 3.070 468.710 2612.530 469.010 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 3.070 466.290 3.370 468.710 ;
        RECT 2612.150 468.700 2612.530 468.710 ;
        RECT -4.800 465.990 3.370 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
      LAYER via3 ;
        RECT 2612.180 2321.020 2612.500 2321.340 ;
        RECT 2612.180 468.700 2612.500 469.020 ;
      LAYER met4 ;
        RECT 2612.175 2321.015 2612.505 2321.345 ;
        RECT 2612.190 469.025 2612.490 2321.015 ;
        RECT 2612.175 468.695 2612.505 469.025 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.650 254.475 16.930 254.845 ;
        RECT 16.720 250.765 16.860 254.475 ;
        RECT 16.650 250.395 16.930 250.765 ;
      LAYER via2 ;
        RECT 16.650 254.520 16.930 254.800 ;
        RECT 16.650 250.440 16.930 250.720 ;
      LAYER met3 ;
        RECT 2610.310 2352.610 2610.690 2352.620 ;
        RECT 2599.460 2352.560 2610.690 2352.610 ;
        RECT 2596.000 2352.310 2610.690 2352.560 ;
        RECT 2596.000 2351.960 2600.000 2352.310 ;
        RECT 2610.310 2352.300 2610.690 2352.310 ;
        RECT 16.625 254.810 16.955 254.825 ;
        RECT 2610.310 254.810 2610.690 254.820 ;
        RECT 16.625 254.510 2610.690 254.810 ;
        RECT 16.625 254.495 16.955 254.510 ;
        RECT 2610.310 254.500 2610.690 254.510 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 16.625 250.730 16.955 250.745 ;
        RECT -4.800 250.430 16.955 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 16.625 250.415 16.955 250.430 ;
      LAYER via3 ;
        RECT 2610.340 2352.300 2610.660 2352.620 ;
        RECT 2610.340 254.500 2610.660 254.820 ;
      LAYER met4 ;
        RECT 2610.335 2352.295 2610.665 2352.625 ;
        RECT 2610.350 254.825 2610.650 2352.295 ;
        RECT 2610.335 254.495 2610.665 254.825 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 40.955 17.390 41.325 ;
        RECT 17.180 35.885 17.320 40.955 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 17.110 41.000 17.390 41.280 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 2608.470 2384.570 2608.850 2384.580 ;
        RECT 2599.460 2384.520 2608.850 2384.570 ;
        RECT 2596.000 2384.270 2608.850 2384.520 ;
        RECT 2596.000 2383.920 2600.000 2384.270 ;
        RECT 2608.470 2384.260 2608.850 2384.270 ;
        RECT 17.085 41.290 17.415 41.305 ;
        RECT 2608.470 41.290 2608.850 41.300 ;
        RECT 17.085 40.990 2608.850 41.290 ;
        RECT 17.085 40.975 17.415 40.990 ;
        RECT 2608.470 40.980 2608.850 40.990 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
      LAYER via3 ;
        RECT 2608.500 2384.260 2608.820 2384.580 ;
        RECT 2608.500 40.980 2608.820 41.300 ;
      LAYER met4 ;
        RECT 2608.495 2384.255 2608.825 2384.585 ;
        RECT 2608.510 41.305 2608.810 2384.255 ;
        RECT 2608.495 40.975 2608.825 41.305 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2613.790 1304.480 2614.110 1304.540 ;
        RECT 2619.770 1304.480 2620.090 1304.540 ;
        RECT 2613.790 1304.340 2620.090 1304.480 ;
        RECT 2613.790 1304.280 2614.110 1304.340 ;
        RECT 2619.770 1304.280 2620.090 1304.340 ;
        RECT 2619.770 910.760 2620.090 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2619.770 910.620 2901.150 910.760 ;
        RECT 2619.770 910.560 2620.090 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 2613.820 1304.280 2614.080 1304.540 ;
        RECT 2619.800 1304.280 2620.060 1304.540 ;
        RECT 2619.800 910.560 2620.060 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 2613.810 1309.835 2614.090 1310.205 ;
        RECT 2613.880 1304.570 2614.020 1309.835 ;
        RECT 2613.820 1304.250 2614.080 1304.570 ;
        RECT 2619.800 1304.250 2620.060 1304.570 ;
        RECT 2619.860 910.850 2620.000 1304.250 ;
        RECT 2619.800 910.530 2620.060 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2613.810 1309.880 2614.090 1310.160 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2613.785 1310.170 2614.115 1310.185 ;
        RECT 2599.460 1310.120 2614.115 1310.170 ;
        RECT 2596.000 1309.870 2614.115 1310.120 ;
        RECT 2596.000 1309.520 2600.000 1309.870 ;
        RECT 2613.785 1309.855 2614.115 1309.870 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2614.250 1145.360 2614.570 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2614.250 1145.220 2901.150 1145.360 ;
        RECT 2614.250 1145.160 2614.570 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2614.280 1145.160 2614.540 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 2614.270 1341.795 2614.550 1342.165 ;
        RECT 2614.340 1145.450 2614.480 1341.795 ;
        RECT 2614.280 1145.130 2614.540 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2614.270 1341.840 2614.550 1342.120 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2614.245 1342.130 2614.575 1342.145 ;
        RECT 2599.460 1342.080 2614.575 1342.130 ;
        RECT 2596.000 1341.830 2614.575 1342.080 ;
        RECT 2596.000 1341.480 2600.000 1341.830 ;
        RECT 2614.245 1341.815 2614.575 1341.830 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2614.250 1376.560 2614.570 1376.620 ;
        RECT 2900.830 1376.560 2901.150 1376.620 ;
        RECT 2614.250 1376.420 2901.150 1376.560 ;
        RECT 2614.250 1376.360 2614.570 1376.420 ;
        RECT 2900.830 1376.360 2901.150 1376.420 ;
      LAYER via ;
        RECT 2614.280 1376.360 2614.540 1376.620 ;
        RECT 2900.860 1376.360 2901.120 1376.620 ;
      LAYER met2 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
        RECT 2900.920 1376.650 2901.060 1378.515 ;
        RECT 2614.280 1376.330 2614.540 1376.650 ;
        RECT 2900.860 1376.330 2901.120 1376.650 ;
        RECT 2614.340 1373.445 2614.480 1376.330 ;
        RECT 2614.270 1373.075 2614.550 1373.445 ;
      LAYER via2 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
        RECT 2614.270 1373.120 2614.550 1373.400 ;
      LAYER met3 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 2614.245 1373.410 2614.575 1373.425 ;
        RECT 2599.460 1373.360 2614.575 1373.410 ;
        RECT 2596.000 1373.110 2614.575 1373.360 ;
        RECT 2596.000 1372.760 2600.000 1373.110 ;
        RECT 2614.245 1373.095 2614.575 1373.110 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2614.250 1407.500 2614.570 1407.560 ;
        RECT 2903.130 1407.500 2903.450 1407.560 ;
        RECT 2614.250 1407.360 2903.450 1407.500 ;
        RECT 2614.250 1407.300 2614.570 1407.360 ;
        RECT 2903.130 1407.300 2903.450 1407.360 ;
      LAYER via ;
        RECT 2614.280 1407.300 2614.540 1407.560 ;
        RECT 2903.160 1407.300 2903.420 1407.560 ;
      LAYER met2 ;
        RECT 2903.150 1613.115 2903.430 1613.485 ;
        RECT 2903.220 1407.590 2903.360 1613.115 ;
        RECT 2614.280 1407.270 2614.540 1407.590 ;
        RECT 2903.160 1407.270 2903.420 1407.590 ;
        RECT 2614.340 1405.405 2614.480 1407.270 ;
        RECT 2614.270 1405.035 2614.550 1405.405 ;
      LAYER via2 ;
        RECT 2903.150 1613.160 2903.430 1613.440 ;
        RECT 2614.270 1405.080 2614.550 1405.360 ;
      LAYER met3 ;
        RECT 2903.125 1613.450 2903.455 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2903.125 1613.150 2924.800 1613.450 ;
        RECT 2903.125 1613.135 2903.455 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 2614.245 1405.370 2614.575 1405.385 ;
        RECT 2599.460 1405.320 2614.575 1405.370 ;
        RECT 2596.000 1405.070 2614.575 1405.320 ;
        RECT 2596.000 1404.720 2600.000 1405.070 ;
        RECT 2614.245 1405.055 2614.575 1405.070 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2614.250 1441.840 2614.570 1441.900 ;
        RECT 2901.750 1441.840 2902.070 1441.900 ;
        RECT 2614.250 1441.700 2902.070 1441.840 ;
        RECT 2614.250 1441.640 2614.570 1441.700 ;
        RECT 2901.750 1441.640 2902.070 1441.700 ;
      LAYER via ;
        RECT 2614.280 1441.640 2614.540 1441.900 ;
        RECT 2901.780 1441.640 2902.040 1441.900 ;
      LAYER met2 ;
        RECT 2901.770 1847.715 2902.050 1848.085 ;
        RECT 2901.840 1441.930 2901.980 1847.715 ;
        RECT 2614.280 1441.610 2614.540 1441.930 ;
        RECT 2901.780 1441.610 2902.040 1441.930 ;
        RECT 2614.340 1436.685 2614.480 1441.610 ;
        RECT 2614.270 1436.315 2614.550 1436.685 ;
      LAYER via2 ;
        RECT 2901.770 1847.760 2902.050 1848.040 ;
        RECT 2614.270 1436.360 2614.550 1436.640 ;
      LAYER met3 ;
        RECT 2901.745 1848.050 2902.075 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2901.745 1847.750 2924.800 1848.050 ;
        RECT 2901.745 1847.735 2902.075 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 2614.245 1436.650 2614.575 1436.665 ;
        RECT 2599.460 1436.600 2614.575 1436.650 ;
        RECT 2596.000 1436.350 2614.575 1436.600 ;
        RECT 2596.000 1436.000 2600.000 1436.350 ;
        RECT 2614.245 1436.335 2614.575 1436.350 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2735.690 2077.300 2736.010 2077.360 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 2735.690 2077.160 2901.150 2077.300 ;
        RECT 2735.690 2077.100 2736.010 2077.160 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
        RECT 2614.250 1469.720 2614.570 1469.780 ;
        RECT 2735.690 1469.720 2736.010 1469.780 ;
        RECT 2614.250 1469.580 2736.010 1469.720 ;
        RECT 2614.250 1469.520 2614.570 1469.580 ;
        RECT 2735.690 1469.520 2736.010 1469.580 ;
      LAYER via ;
        RECT 2735.720 2077.100 2735.980 2077.360 ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
        RECT 2614.280 1469.520 2614.540 1469.780 ;
        RECT 2735.720 1469.520 2735.980 1469.780 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 2735.720 2077.070 2735.980 2077.390 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
        RECT 2735.780 1469.810 2735.920 2077.070 ;
        RECT 2614.280 1469.490 2614.540 1469.810 ;
        RECT 2735.720 1469.490 2735.980 1469.810 ;
        RECT 2614.340 1468.645 2614.480 1469.490 ;
        RECT 2614.270 1468.275 2614.550 1468.645 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
        RECT 2614.270 1468.320 2614.550 1468.600 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 2614.245 1468.610 2614.575 1468.625 ;
        RECT 2599.460 1468.560 2614.575 1468.610 ;
        RECT 2596.000 1468.310 2614.575 1468.560 ;
        RECT 2596.000 1467.960 2600.000 1468.310 ;
        RECT 2614.245 1468.295 2614.575 1468.310 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2749.490 2311.900 2749.810 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2749.490 2311.760 2901.150 2311.900 ;
        RECT 2749.490 2311.700 2749.810 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
        RECT 2614.250 1504.060 2614.570 1504.120 ;
        RECT 2749.490 1504.060 2749.810 1504.120 ;
        RECT 2614.250 1503.920 2749.810 1504.060 ;
        RECT 2614.250 1503.860 2614.570 1503.920 ;
        RECT 2749.490 1503.860 2749.810 1503.920 ;
      LAYER via ;
        RECT 2749.520 2311.700 2749.780 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
        RECT 2614.280 1503.860 2614.540 1504.120 ;
        RECT 2749.520 1503.860 2749.780 1504.120 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2749.520 2311.670 2749.780 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 2749.580 1504.150 2749.720 2311.670 ;
        RECT 2614.280 1503.830 2614.540 1504.150 ;
        RECT 2749.520 1503.830 2749.780 1504.150 ;
        RECT 2614.340 1499.925 2614.480 1503.830 ;
        RECT 2614.270 1499.555 2614.550 1499.925 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 2614.270 1499.600 2614.550 1499.880 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2614.245 1499.890 2614.575 1499.905 ;
        RECT 2599.460 1499.840 2614.575 1499.890 ;
        RECT 2596.000 1499.590 2614.575 1499.840 ;
        RECT 2596.000 1499.240 2600.000 1499.590 ;
        RECT 2614.245 1499.575 2614.575 1499.590 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2608.270 151.540 2608.590 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2608.270 151.400 2901.150 151.540 ;
        RECT 2608.270 151.340 2608.590 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 2608.300 151.340 2608.560 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 2608.290 1225.515 2608.570 1225.885 ;
        RECT 2608.360 151.630 2608.500 1225.515 ;
        RECT 2608.300 151.310 2608.560 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2608.290 1225.560 2608.570 1225.840 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 2608.265 1225.850 2608.595 1225.865 ;
        RECT 2599.460 1225.800 2608.595 1225.850 ;
        RECT 2596.000 1225.550 2608.595 1225.800 ;
        RECT 2596.000 1225.200 2600.000 1225.550 ;
        RECT 2608.265 1225.535 2608.595 1225.550 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2770.190 2491.080 2770.510 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 2770.190 2490.940 2901.150 2491.080 ;
        RECT 2770.190 2490.880 2770.510 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
        RECT 2614.250 1545.540 2614.570 1545.600 ;
        RECT 2770.190 1545.540 2770.510 1545.600 ;
        RECT 2614.250 1545.400 2770.510 1545.540 ;
        RECT 2614.250 1545.340 2614.570 1545.400 ;
        RECT 2770.190 1545.340 2770.510 1545.400 ;
      LAYER via ;
        RECT 2770.220 2490.880 2770.480 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
        RECT 2614.280 1545.340 2614.540 1545.600 ;
        RECT 2770.220 1545.340 2770.480 1545.600 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 2770.220 2490.850 2770.480 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 2770.280 1545.630 2770.420 2490.850 ;
        RECT 2614.280 1545.310 2614.540 1545.630 ;
        RECT 2770.220 1545.310 2770.480 1545.630 ;
        RECT 2614.340 1542.085 2614.480 1545.310 ;
        RECT 2614.270 1541.715 2614.550 1542.085 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
        RECT 2614.270 1541.760 2614.550 1542.040 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 2614.245 1542.050 2614.575 1542.065 ;
        RECT 2599.460 1542.000 2614.575 1542.050 ;
        RECT 2596.000 1541.750 2614.575 1542.000 ;
        RECT 2596.000 1541.400 2600.000 1541.750 ;
        RECT 2614.245 1541.735 2614.575 1541.750 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2777.090 2725.680 2777.410 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 2777.090 2725.540 2901.150 2725.680 ;
        RECT 2777.090 2725.480 2777.410 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
        RECT 2614.250 1573.080 2614.570 1573.140 ;
        RECT 2777.090 1573.080 2777.410 1573.140 ;
        RECT 2614.250 1572.940 2777.410 1573.080 ;
        RECT 2614.250 1572.880 2614.570 1572.940 ;
        RECT 2777.090 1572.880 2777.410 1572.940 ;
      LAYER via ;
        RECT 2777.120 2725.480 2777.380 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
        RECT 2614.280 1572.880 2614.540 1573.140 ;
        RECT 2777.120 1572.880 2777.380 1573.140 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 2777.120 2725.450 2777.380 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 2614.270 1572.995 2614.550 1573.365 ;
        RECT 2777.180 1573.170 2777.320 2725.450 ;
        RECT 2614.280 1572.850 2614.540 1572.995 ;
        RECT 2777.120 1572.850 2777.380 1573.170 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
        RECT 2614.270 1573.040 2614.550 1573.320 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2614.245 1573.330 2614.575 1573.345 ;
        RECT 2599.460 1573.280 2614.575 1573.330 ;
        RECT 2596.000 1573.030 2614.575 1573.280 ;
        RECT 2596.000 1572.680 2600.000 1573.030 ;
        RECT 2614.245 1573.015 2614.575 1573.030 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2783.990 2960.280 2784.310 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 2783.990 2960.140 2901.150 2960.280 ;
        RECT 2783.990 2960.080 2784.310 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
        RECT 2614.250 1607.760 2614.570 1607.820 ;
        RECT 2783.990 1607.760 2784.310 1607.820 ;
        RECT 2614.250 1607.620 2784.310 1607.760 ;
        RECT 2614.250 1607.560 2614.570 1607.620 ;
        RECT 2783.990 1607.560 2784.310 1607.620 ;
      LAYER via ;
        RECT 2784.020 2960.080 2784.280 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
        RECT 2614.280 1607.560 2614.540 1607.820 ;
        RECT 2784.020 1607.560 2784.280 1607.820 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 2784.020 2960.050 2784.280 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 2784.080 1607.850 2784.220 2960.050 ;
        RECT 2614.280 1607.530 2614.540 1607.850 ;
        RECT 2784.020 1607.530 2784.280 1607.850 ;
        RECT 2614.340 1605.325 2614.480 1607.530 ;
        RECT 2614.270 1604.955 2614.550 1605.325 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
        RECT 2614.270 1605.000 2614.550 1605.280 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 2614.245 1605.290 2614.575 1605.305 ;
        RECT 2599.460 1605.240 2614.575 1605.290 ;
        RECT 2596.000 1604.990 2614.575 1605.240 ;
        RECT 2596.000 1604.640 2600.000 1604.990 ;
        RECT 2614.245 1604.975 2614.575 1604.990 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2790.890 3194.880 2791.210 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 2790.890 3194.740 2901.150 3194.880 ;
        RECT 2790.890 3194.680 2791.210 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
        RECT 2614.250 1642.100 2614.570 1642.160 ;
        RECT 2790.890 1642.100 2791.210 1642.160 ;
        RECT 2614.250 1641.960 2791.210 1642.100 ;
        RECT 2614.250 1641.900 2614.570 1641.960 ;
        RECT 2790.890 1641.900 2791.210 1641.960 ;
      LAYER via ;
        RECT 2790.920 3194.680 2791.180 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
        RECT 2614.280 1641.900 2614.540 1642.160 ;
        RECT 2790.920 1641.900 2791.180 1642.160 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 2790.920 3194.650 2791.180 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 2790.980 1642.190 2791.120 3194.650 ;
        RECT 2614.280 1641.870 2614.540 1642.190 ;
        RECT 2790.920 1641.870 2791.180 1642.190 ;
        RECT 2614.340 1636.605 2614.480 1641.870 ;
        RECT 2614.270 1636.235 2614.550 1636.605 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 2614.270 1636.280 2614.550 1636.560 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 2614.245 1636.570 2614.575 1636.585 ;
        RECT 2599.460 1636.520 2614.575 1636.570 ;
        RECT 2596.000 1636.270 2614.575 1636.520 ;
        RECT 2596.000 1635.920 2600.000 1636.270 ;
        RECT 2614.245 1636.255 2614.575 1636.270 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2804.690 3429.480 2805.010 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2804.690 3429.340 2901.150 3429.480 ;
        RECT 2804.690 3429.280 2805.010 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
        RECT 2614.250 1669.640 2614.570 1669.700 ;
        RECT 2804.690 1669.640 2805.010 1669.700 ;
        RECT 2614.250 1669.500 2805.010 1669.640 ;
        RECT 2614.250 1669.440 2614.570 1669.500 ;
        RECT 2804.690 1669.440 2805.010 1669.500 ;
      LAYER via ;
        RECT 2804.720 3429.280 2804.980 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
        RECT 2614.280 1669.440 2614.540 1669.700 ;
        RECT 2804.720 1669.440 2804.980 1669.700 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 2804.720 3429.250 2804.980 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 2804.780 1669.730 2804.920 3429.250 ;
        RECT 2614.280 1669.410 2614.540 1669.730 ;
        RECT 2804.720 1669.410 2804.980 1669.730 ;
        RECT 2614.340 1668.565 2614.480 1669.410 ;
        RECT 2614.270 1668.195 2614.550 1668.565 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 2614.270 1668.240 2614.550 1668.520 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2614.245 1668.530 2614.575 1668.545 ;
        RECT 2599.460 1668.480 2614.575 1668.530 ;
        RECT 2596.000 1668.230 2614.575 1668.480 ;
        RECT 2596.000 1667.880 2600.000 1668.230 ;
        RECT 2614.245 1668.215 2614.575 1668.230 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2713.610 3491.360 2713.930 3491.420 ;
        RECT 2717.750 3491.360 2718.070 3491.420 ;
        RECT 2713.610 3491.220 2718.070 3491.360 ;
        RECT 2713.610 3491.160 2713.930 3491.220 ;
        RECT 2717.750 3491.160 2718.070 3491.220 ;
        RECT 2712.690 3470.620 2713.010 3470.680 ;
        RECT 2713.610 3470.620 2713.930 3470.680 ;
        RECT 2712.690 3470.480 2713.930 3470.620 ;
        RECT 2712.690 3470.420 2713.010 3470.480 ;
        RECT 2713.610 3470.420 2713.930 3470.480 ;
        RECT 2712.230 3422.680 2712.550 3422.740 ;
        RECT 2712.690 3422.680 2713.010 3422.740 ;
        RECT 2712.230 3422.540 2713.010 3422.680 ;
        RECT 2712.230 3422.480 2712.550 3422.540 ;
        RECT 2712.690 3422.480 2713.010 3422.540 ;
        RECT 2712.690 3332.920 2713.010 3332.980 ;
        RECT 2714.070 3332.920 2714.390 3332.980 ;
        RECT 2712.690 3332.780 2714.390 3332.920 ;
        RECT 2712.690 3332.720 2713.010 3332.780 ;
        RECT 2714.070 3332.720 2714.390 3332.780 ;
        RECT 2712.690 3308.780 2713.010 3308.840 ;
        RECT 2714.070 3308.780 2714.390 3308.840 ;
        RECT 2712.690 3308.640 2714.390 3308.780 ;
        RECT 2712.690 3308.580 2713.010 3308.640 ;
        RECT 2714.070 3308.580 2714.390 3308.640 ;
        RECT 2712.690 3284.640 2713.010 3284.700 ;
        RECT 2713.150 3284.640 2713.470 3284.700 ;
        RECT 2712.690 3284.500 2713.470 3284.640 ;
        RECT 2712.690 3284.440 2713.010 3284.500 ;
        RECT 2713.150 3284.440 2713.470 3284.500 ;
        RECT 2712.690 3236.360 2713.010 3236.420 ;
        RECT 2713.150 3236.360 2713.470 3236.420 ;
        RECT 2712.690 3236.220 2713.470 3236.360 ;
        RECT 2712.690 3236.160 2713.010 3236.220 ;
        RECT 2713.150 3236.160 2713.470 3236.220 ;
        RECT 2712.690 3202.020 2713.010 3202.080 ;
        RECT 2713.150 3202.020 2713.470 3202.080 ;
        RECT 2712.690 3201.880 2713.470 3202.020 ;
        RECT 2712.690 3201.820 2713.010 3201.880 ;
        RECT 2713.150 3201.820 2713.470 3201.880 ;
        RECT 2712.230 3153.400 2712.550 3153.460 ;
        RECT 2713.150 3153.400 2713.470 3153.460 ;
        RECT 2712.230 3153.260 2713.470 3153.400 ;
        RECT 2712.230 3153.200 2712.550 3153.260 ;
        RECT 2713.150 3153.200 2713.470 3153.260 ;
        RECT 2712.230 3056.840 2712.550 3056.900 ;
        RECT 2713.150 3056.840 2713.470 3056.900 ;
        RECT 2712.230 3056.700 2713.470 3056.840 ;
        RECT 2712.230 3056.640 2712.550 3056.700 ;
        RECT 2713.150 3056.640 2713.470 3056.700 ;
        RECT 2712.230 3042.900 2712.550 3042.960 ;
        RECT 2712.690 3042.900 2713.010 3042.960 ;
        RECT 2712.230 3042.760 2713.010 3042.900 ;
        RECT 2712.230 3042.700 2712.550 3042.760 ;
        RECT 2712.690 3042.700 2713.010 3042.760 ;
        RECT 2712.230 3008.560 2712.550 3008.620 ;
        RECT 2713.610 3008.560 2713.930 3008.620 ;
        RECT 2712.230 3008.420 2713.930 3008.560 ;
        RECT 2712.230 3008.360 2712.550 3008.420 ;
        RECT 2713.610 3008.360 2713.930 3008.420 ;
        RECT 2712.690 2994.620 2713.010 2994.680 ;
        RECT 2713.610 2994.620 2713.930 2994.680 ;
        RECT 2712.690 2994.480 2713.930 2994.620 ;
        RECT 2712.690 2994.420 2713.010 2994.480 ;
        RECT 2713.610 2994.420 2713.930 2994.480 ;
        RECT 2712.690 2946.680 2713.010 2946.740 ;
        RECT 2714.070 2946.680 2714.390 2946.740 ;
        RECT 2712.690 2946.540 2714.390 2946.680 ;
        RECT 2712.690 2946.480 2713.010 2946.540 ;
        RECT 2714.070 2946.480 2714.390 2946.540 ;
        RECT 2714.070 2912.340 2714.390 2912.400 ;
        RECT 2713.700 2912.200 2714.390 2912.340 ;
        RECT 2713.700 2911.720 2713.840 2912.200 ;
        RECT 2714.070 2912.140 2714.390 2912.200 ;
        RECT 2713.610 2911.460 2713.930 2911.720 ;
        RECT 2712.230 2815.580 2712.550 2815.840 ;
        RECT 2712.320 2815.160 2712.460 2815.580 ;
        RECT 2712.230 2814.900 2712.550 2815.160 ;
        RECT 2711.770 2767.160 2712.090 2767.220 ;
        RECT 2711.770 2767.020 2712.460 2767.160 ;
        RECT 2711.770 2766.960 2712.090 2767.020 ;
        RECT 2712.320 2766.880 2712.460 2767.020 ;
        RECT 2712.230 2766.620 2712.550 2766.880 ;
        RECT 2711.770 2753.220 2712.090 2753.280 ;
        RECT 2712.230 2753.220 2712.550 2753.280 ;
        RECT 2711.770 2753.080 2712.550 2753.220 ;
        RECT 2711.770 2753.020 2712.090 2753.080 ;
        RECT 2712.230 2753.020 2712.550 2753.080 ;
        RECT 2711.770 2718.680 2712.090 2718.940 ;
        RECT 2711.860 2718.200 2712.000 2718.680 ;
        RECT 2712.230 2718.200 2712.550 2718.260 ;
        RECT 2711.860 2718.060 2712.550 2718.200 ;
        RECT 2712.230 2718.000 2712.550 2718.060 ;
        RECT 2712.230 2670.260 2712.550 2670.320 ;
        RECT 2713.150 2670.260 2713.470 2670.320 ;
        RECT 2712.230 2670.120 2713.470 2670.260 ;
        RECT 2712.230 2670.060 2712.550 2670.120 ;
        RECT 2713.150 2670.060 2713.470 2670.120 ;
        RECT 2713.150 2622.120 2713.470 2622.380 ;
        RECT 2713.240 2621.980 2713.380 2622.120 ;
        RECT 2713.610 2621.980 2713.930 2622.040 ;
        RECT 2713.240 2621.840 2713.930 2621.980 ;
        RECT 2713.610 2621.780 2713.930 2621.840 ;
        RECT 2712.690 2560.100 2713.010 2560.160 ;
        RECT 2714.070 2560.100 2714.390 2560.160 ;
        RECT 2712.690 2559.960 2714.390 2560.100 ;
        RECT 2712.690 2559.900 2713.010 2559.960 ;
        RECT 2714.070 2559.900 2714.390 2559.960 ;
        RECT 2713.150 2511.820 2713.470 2511.880 ;
        RECT 2714.070 2511.820 2714.390 2511.880 ;
        RECT 2713.150 2511.680 2714.390 2511.820 ;
        RECT 2713.150 2511.620 2713.470 2511.680 ;
        RECT 2714.070 2511.620 2714.390 2511.680 ;
        RECT 2712.690 2463.200 2713.010 2463.260 ;
        RECT 2713.150 2463.200 2713.470 2463.260 ;
        RECT 2712.690 2463.060 2713.470 2463.200 ;
        RECT 2712.690 2463.000 2713.010 2463.060 ;
        RECT 2713.150 2463.000 2713.470 2463.060 ;
        RECT 2712.690 2428.860 2713.010 2428.920 ;
        RECT 2713.150 2428.860 2713.470 2428.920 ;
        RECT 2712.690 2428.720 2713.470 2428.860 ;
        RECT 2712.690 2428.660 2713.010 2428.720 ;
        RECT 2713.150 2428.660 2713.470 2428.720 ;
        RECT 2712.230 2380.580 2712.550 2380.640 ;
        RECT 2713.150 2380.580 2713.470 2380.640 ;
        RECT 2712.230 2380.440 2713.470 2380.580 ;
        RECT 2712.230 2380.380 2712.550 2380.440 ;
        RECT 2713.150 2380.380 2713.470 2380.440 ;
        RECT 2712.690 2366.640 2713.010 2366.700 ;
        RECT 2713.150 2366.640 2713.470 2366.700 ;
        RECT 2712.690 2366.500 2713.470 2366.640 ;
        RECT 2712.690 2366.440 2713.010 2366.500 ;
        RECT 2713.150 2366.440 2713.470 2366.500 ;
        RECT 2713.150 2332.300 2713.470 2332.360 ;
        RECT 2712.780 2332.160 2713.470 2332.300 ;
        RECT 2712.780 2332.020 2712.920 2332.160 ;
        RECT 2713.150 2332.100 2713.470 2332.160 ;
        RECT 2712.690 2331.760 2713.010 2332.020 ;
        RECT 2711.770 2235.540 2712.090 2235.800 ;
        RECT 2711.860 2235.400 2712.000 2235.540 ;
        RECT 2712.230 2235.400 2712.550 2235.460 ;
        RECT 2711.860 2235.260 2712.550 2235.400 ;
        RECT 2712.230 2235.200 2712.550 2235.260 ;
        RECT 2710.850 2221.800 2711.170 2221.860 ;
        RECT 2712.230 2221.800 2712.550 2221.860 ;
        RECT 2710.850 2221.660 2712.550 2221.800 ;
        RECT 2710.850 2221.600 2711.170 2221.660 ;
        RECT 2712.230 2221.600 2712.550 2221.660 ;
        RECT 2711.770 2138.980 2712.090 2139.240 ;
        RECT 2711.860 2138.840 2712.000 2138.980 ;
        RECT 2712.230 2138.840 2712.550 2138.900 ;
        RECT 2711.860 2138.700 2712.550 2138.840 ;
        RECT 2712.230 2138.640 2712.550 2138.700 ;
        RECT 2710.850 2125.240 2711.170 2125.300 ;
        RECT 2712.230 2125.240 2712.550 2125.300 ;
        RECT 2710.850 2125.100 2712.550 2125.240 ;
        RECT 2710.850 2125.040 2711.170 2125.100 ;
        RECT 2712.230 2125.040 2712.550 2125.100 ;
        RECT 2711.770 2042.420 2712.090 2042.680 ;
        RECT 2711.860 2041.940 2712.000 2042.420 ;
        RECT 2712.230 2041.940 2712.550 2042.000 ;
        RECT 2711.860 2041.800 2712.550 2041.940 ;
        RECT 2712.230 2041.740 2712.550 2041.800 ;
        RECT 2710.390 2021.540 2710.710 2021.600 ;
        RECT 2712.230 2021.540 2712.550 2021.600 ;
        RECT 2710.390 2021.400 2712.550 2021.540 ;
        RECT 2710.390 2021.340 2710.710 2021.400 ;
        RECT 2712.230 2021.340 2712.550 2021.400 ;
        RECT 2710.850 1966.460 2711.170 1966.520 ;
        RECT 2711.770 1966.460 2712.090 1966.520 ;
        RECT 2710.850 1966.320 2712.090 1966.460 ;
        RECT 2710.850 1966.260 2711.170 1966.320 ;
        RECT 2711.770 1966.260 2712.090 1966.320 ;
        RECT 2710.850 1918.520 2711.170 1918.580 ;
        RECT 2712.230 1918.520 2712.550 1918.580 ;
        RECT 2710.850 1918.380 2712.550 1918.520 ;
        RECT 2710.850 1918.320 2711.170 1918.380 ;
        RECT 2712.230 1918.320 2712.550 1918.380 ;
        RECT 2712.230 1897.440 2712.550 1897.500 ;
        RECT 2713.150 1897.440 2713.470 1897.500 ;
        RECT 2712.230 1897.300 2713.470 1897.440 ;
        RECT 2712.230 1897.240 2712.550 1897.300 ;
        RECT 2713.150 1897.240 2713.470 1897.300 ;
        RECT 2712.230 1835.220 2712.550 1835.280 ;
        RECT 2713.610 1835.220 2713.930 1835.280 ;
        RECT 2712.230 1835.080 2713.930 1835.220 ;
        RECT 2712.230 1835.020 2712.550 1835.080 ;
        RECT 2713.610 1835.020 2713.930 1835.080 ;
        RECT 2712.230 1787.280 2712.550 1787.340 ;
        RECT 2712.690 1787.280 2713.010 1787.340 ;
        RECT 2712.230 1787.140 2713.010 1787.280 ;
        RECT 2712.230 1787.080 2712.550 1787.140 ;
        RECT 2712.690 1787.080 2713.010 1787.140 ;
        RECT 2712.690 1752.740 2713.010 1753.000 ;
        RECT 2712.780 1752.600 2712.920 1752.740 ;
        RECT 2713.610 1752.600 2713.930 1752.660 ;
        RECT 2712.780 1752.460 2713.930 1752.600 ;
        RECT 2713.610 1752.400 2713.930 1752.460 ;
        RECT 2614.250 1704.320 2614.570 1704.380 ;
        RECT 2713.610 1704.320 2713.930 1704.380 ;
        RECT 2614.250 1704.180 2713.930 1704.320 ;
        RECT 2614.250 1704.120 2614.570 1704.180 ;
        RECT 2713.610 1704.120 2713.930 1704.180 ;
      LAYER via ;
        RECT 2713.640 3491.160 2713.900 3491.420 ;
        RECT 2717.780 3491.160 2718.040 3491.420 ;
        RECT 2712.720 3470.420 2712.980 3470.680 ;
        RECT 2713.640 3470.420 2713.900 3470.680 ;
        RECT 2712.260 3422.480 2712.520 3422.740 ;
        RECT 2712.720 3422.480 2712.980 3422.740 ;
        RECT 2712.720 3332.720 2712.980 3332.980 ;
        RECT 2714.100 3332.720 2714.360 3332.980 ;
        RECT 2712.720 3308.580 2712.980 3308.840 ;
        RECT 2714.100 3308.580 2714.360 3308.840 ;
        RECT 2712.720 3284.440 2712.980 3284.700 ;
        RECT 2713.180 3284.440 2713.440 3284.700 ;
        RECT 2712.720 3236.160 2712.980 3236.420 ;
        RECT 2713.180 3236.160 2713.440 3236.420 ;
        RECT 2712.720 3201.820 2712.980 3202.080 ;
        RECT 2713.180 3201.820 2713.440 3202.080 ;
        RECT 2712.260 3153.200 2712.520 3153.460 ;
        RECT 2713.180 3153.200 2713.440 3153.460 ;
        RECT 2712.260 3056.640 2712.520 3056.900 ;
        RECT 2713.180 3056.640 2713.440 3056.900 ;
        RECT 2712.260 3042.700 2712.520 3042.960 ;
        RECT 2712.720 3042.700 2712.980 3042.960 ;
        RECT 2712.260 3008.360 2712.520 3008.620 ;
        RECT 2713.640 3008.360 2713.900 3008.620 ;
        RECT 2712.720 2994.420 2712.980 2994.680 ;
        RECT 2713.640 2994.420 2713.900 2994.680 ;
        RECT 2712.720 2946.480 2712.980 2946.740 ;
        RECT 2714.100 2946.480 2714.360 2946.740 ;
        RECT 2714.100 2912.140 2714.360 2912.400 ;
        RECT 2713.640 2911.460 2713.900 2911.720 ;
        RECT 2712.260 2815.580 2712.520 2815.840 ;
        RECT 2712.260 2814.900 2712.520 2815.160 ;
        RECT 2711.800 2766.960 2712.060 2767.220 ;
        RECT 2712.260 2766.620 2712.520 2766.880 ;
        RECT 2711.800 2753.020 2712.060 2753.280 ;
        RECT 2712.260 2753.020 2712.520 2753.280 ;
        RECT 2711.800 2718.680 2712.060 2718.940 ;
        RECT 2712.260 2718.000 2712.520 2718.260 ;
        RECT 2712.260 2670.060 2712.520 2670.320 ;
        RECT 2713.180 2670.060 2713.440 2670.320 ;
        RECT 2713.180 2622.120 2713.440 2622.380 ;
        RECT 2713.640 2621.780 2713.900 2622.040 ;
        RECT 2712.720 2559.900 2712.980 2560.160 ;
        RECT 2714.100 2559.900 2714.360 2560.160 ;
        RECT 2713.180 2511.620 2713.440 2511.880 ;
        RECT 2714.100 2511.620 2714.360 2511.880 ;
        RECT 2712.720 2463.000 2712.980 2463.260 ;
        RECT 2713.180 2463.000 2713.440 2463.260 ;
        RECT 2712.720 2428.660 2712.980 2428.920 ;
        RECT 2713.180 2428.660 2713.440 2428.920 ;
        RECT 2712.260 2380.380 2712.520 2380.640 ;
        RECT 2713.180 2380.380 2713.440 2380.640 ;
        RECT 2712.720 2366.440 2712.980 2366.700 ;
        RECT 2713.180 2366.440 2713.440 2366.700 ;
        RECT 2713.180 2332.100 2713.440 2332.360 ;
        RECT 2712.720 2331.760 2712.980 2332.020 ;
        RECT 2711.800 2235.540 2712.060 2235.800 ;
        RECT 2712.260 2235.200 2712.520 2235.460 ;
        RECT 2710.880 2221.600 2711.140 2221.860 ;
        RECT 2712.260 2221.600 2712.520 2221.860 ;
        RECT 2711.800 2138.980 2712.060 2139.240 ;
        RECT 2712.260 2138.640 2712.520 2138.900 ;
        RECT 2710.880 2125.040 2711.140 2125.300 ;
        RECT 2712.260 2125.040 2712.520 2125.300 ;
        RECT 2711.800 2042.420 2712.060 2042.680 ;
        RECT 2712.260 2041.740 2712.520 2042.000 ;
        RECT 2710.420 2021.340 2710.680 2021.600 ;
        RECT 2712.260 2021.340 2712.520 2021.600 ;
        RECT 2710.880 1966.260 2711.140 1966.520 ;
        RECT 2711.800 1966.260 2712.060 1966.520 ;
        RECT 2710.880 1918.320 2711.140 1918.580 ;
        RECT 2712.260 1918.320 2712.520 1918.580 ;
        RECT 2712.260 1897.240 2712.520 1897.500 ;
        RECT 2713.180 1897.240 2713.440 1897.500 ;
        RECT 2712.260 1835.020 2712.520 1835.280 ;
        RECT 2713.640 1835.020 2713.900 1835.280 ;
        RECT 2712.260 1787.080 2712.520 1787.340 ;
        RECT 2712.720 1787.080 2712.980 1787.340 ;
        RECT 2712.720 1752.740 2712.980 1753.000 ;
        RECT 2713.640 1752.400 2713.900 1752.660 ;
        RECT 2614.280 1704.120 2614.540 1704.380 ;
        RECT 2713.640 1704.120 2713.900 1704.380 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3517.370 2717.520 3517.600 ;
        RECT 2717.380 3517.230 2717.980 3517.370 ;
        RECT 2717.840 3491.450 2717.980 3517.230 ;
        RECT 2713.640 3491.130 2713.900 3491.450 ;
        RECT 2717.780 3491.130 2718.040 3491.450 ;
        RECT 2713.700 3470.710 2713.840 3491.130 ;
        RECT 2712.720 3470.390 2712.980 3470.710 ;
        RECT 2713.640 3470.390 2713.900 3470.710 ;
        RECT 2712.780 3422.770 2712.920 3470.390 ;
        RECT 2712.260 3422.450 2712.520 3422.770 ;
        RECT 2712.720 3422.450 2712.980 3422.770 ;
        RECT 2712.320 3422.285 2712.460 3422.450 ;
        RECT 2712.250 3421.915 2712.530 3422.285 ;
        RECT 2712.710 3394.035 2712.990 3394.405 ;
        RECT 2712.780 3333.010 2712.920 3394.035 ;
        RECT 2712.720 3332.690 2712.980 3333.010 ;
        RECT 2714.100 3332.690 2714.360 3333.010 ;
        RECT 2714.160 3308.870 2714.300 3332.690 ;
        RECT 2712.720 3308.550 2712.980 3308.870 ;
        RECT 2714.100 3308.550 2714.360 3308.870 ;
        RECT 2712.780 3284.730 2712.920 3308.550 ;
        RECT 2712.720 3284.410 2712.980 3284.730 ;
        RECT 2713.180 3284.410 2713.440 3284.730 ;
        RECT 2713.240 3236.450 2713.380 3284.410 ;
        RECT 2712.720 3236.130 2712.980 3236.450 ;
        RECT 2713.180 3236.130 2713.440 3236.450 ;
        RECT 2712.780 3202.110 2712.920 3236.130 ;
        RECT 2712.720 3201.790 2712.980 3202.110 ;
        RECT 2713.180 3201.790 2713.440 3202.110 ;
        RECT 2713.240 3153.490 2713.380 3201.790 ;
        RECT 2712.260 3153.170 2712.520 3153.490 ;
        RECT 2713.180 3153.170 2713.440 3153.490 ;
        RECT 2712.320 3152.890 2712.460 3153.170 ;
        RECT 2712.320 3152.750 2712.920 3152.890 ;
        RECT 2712.780 3105.290 2712.920 3152.750 ;
        RECT 2712.780 3105.150 2713.380 3105.290 ;
        RECT 2713.240 3056.930 2713.380 3105.150 ;
        RECT 2712.260 3056.610 2712.520 3056.930 ;
        RECT 2713.180 3056.610 2713.440 3056.930 ;
        RECT 2712.320 3056.330 2712.460 3056.610 ;
        RECT 2712.320 3056.190 2712.920 3056.330 ;
        RECT 2712.780 3042.990 2712.920 3056.190 ;
        RECT 2712.260 3042.670 2712.520 3042.990 ;
        RECT 2712.720 3042.670 2712.980 3042.990 ;
        RECT 2712.320 3008.650 2712.460 3042.670 ;
        RECT 2712.260 3008.330 2712.520 3008.650 ;
        RECT 2713.640 3008.330 2713.900 3008.650 ;
        RECT 2713.700 2994.710 2713.840 3008.330 ;
        RECT 2712.720 2994.390 2712.980 2994.710 ;
        RECT 2713.640 2994.390 2713.900 2994.710 ;
        RECT 2712.780 2946.770 2712.920 2994.390 ;
        RECT 2712.720 2946.450 2712.980 2946.770 ;
        RECT 2714.100 2946.450 2714.360 2946.770 ;
        RECT 2714.160 2912.430 2714.300 2946.450 ;
        RECT 2714.100 2912.110 2714.360 2912.430 ;
        RECT 2713.640 2911.430 2713.900 2911.750 ;
        RECT 2713.700 2863.210 2713.840 2911.430 ;
        RECT 2712.780 2863.070 2713.840 2863.210 ;
        RECT 2712.780 2849.610 2712.920 2863.070 ;
        RECT 2712.320 2849.470 2712.920 2849.610 ;
        RECT 2712.320 2815.870 2712.460 2849.470 ;
        RECT 2712.260 2815.550 2712.520 2815.870 ;
        RECT 2712.260 2814.870 2712.520 2815.190 ;
        RECT 2712.320 2801.330 2712.460 2814.870 ;
        RECT 2711.860 2801.190 2712.460 2801.330 ;
        RECT 2711.860 2767.250 2712.000 2801.190 ;
        RECT 2711.800 2766.930 2712.060 2767.250 ;
        RECT 2712.260 2766.590 2712.520 2766.910 ;
        RECT 2712.320 2753.310 2712.460 2766.590 ;
        RECT 2711.800 2752.990 2712.060 2753.310 ;
        RECT 2712.260 2752.990 2712.520 2753.310 ;
        RECT 2711.860 2718.970 2712.000 2752.990 ;
        RECT 2711.800 2718.650 2712.060 2718.970 ;
        RECT 2712.260 2717.970 2712.520 2718.290 ;
        RECT 2712.320 2670.350 2712.460 2717.970 ;
        RECT 2712.260 2670.030 2712.520 2670.350 ;
        RECT 2713.180 2670.030 2713.440 2670.350 ;
        RECT 2713.240 2622.410 2713.380 2670.030 ;
        RECT 2713.180 2622.090 2713.440 2622.410 ;
        RECT 2713.640 2621.750 2713.900 2622.070 ;
        RECT 2713.700 2608.325 2713.840 2621.750 ;
        RECT 2712.710 2607.955 2712.990 2608.325 ;
        RECT 2713.630 2607.955 2713.910 2608.325 ;
        RECT 2712.780 2560.190 2712.920 2607.955 ;
        RECT 2712.720 2559.870 2712.980 2560.190 ;
        RECT 2714.100 2559.870 2714.360 2560.190 ;
        RECT 2714.160 2511.910 2714.300 2559.870 ;
        RECT 2713.180 2511.590 2713.440 2511.910 ;
        RECT 2714.100 2511.590 2714.360 2511.910 ;
        RECT 2713.240 2464.165 2713.380 2511.590 ;
        RECT 2713.170 2463.795 2713.450 2464.165 ;
        RECT 2712.710 2463.115 2712.990 2463.485 ;
        RECT 2712.720 2462.970 2712.980 2463.115 ;
        RECT 2713.180 2462.970 2713.440 2463.290 ;
        RECT 2713.240 2428.950 2713.380 2462.970 ;
        RECT 2712.720 2428.630 2712.980 2428.950 ;
        RECT 2713.180 2428.630 2713.440 2428.950 ;
        RECT 2712.780 2415.090 2712.920 2428.630 ;
        RECT 2712.780 2414.950 2713.380 2415.090 ;
        RECT 2713.240 2380.670 2713.380 2414.950 ;
        RECT 2712.260 2380.410 2712.520 2380.670 ;
        RECT 2712.260 2380.350 2712.920 2380.410 ;
        RECT 2713.180 2380.350 2713.440 2380.670 ;
        RECT 2712.320 2380.270 2712.920 2380.350 ;
        RECT 2712.780 2366.730 2712.920 2380.270 ;
        RECT 2712.720 2366.410 2712.980 2366.730 ;
        RECT 2713.180 2366.410 2713.440 2366.730 ;
        RECT 2713.240 2332.390 2713.380 2366.410 ;
        RECT 2713.180 2332.070 2713.440 2332.390 ;
        RECT 2712.720 2331.730 2712.980 2332.050 ;
        RECT 2712.780 2318.530 2712.920 2331.730 ;
        RECT 2712.780 2318.390 2713.380 2318.530 ;
        RECT 2713.240 2270.365 2713.380 2318.390 ;
        RECT 2711.790 2269.995 2712.070 2270.365 ;
        RECT 2713.170 2269.995 2713.450 2270.365 ;
        RECT 2711.860 2235.830 2712.000 2269.995 ;
        RECT 2711.800 2235.510 2712.060 2235.830 ;
        RECT 2712.260 2235.170 2712.520 2235.490 ;
        RECT 2712.320 2221.890 2712.460 2235.170 ;
        RECT 2710.880 2221.570 2711.140 2221.890 ;
        RECT 2712.260 2221.570 2712.520 2221.890 ;
        RECT 2710.940 2173.805 2711.080 2221.570 ;
        RECT 2710.870 2173.435 2711.150 2173.805 ;
        RECT 2711.790 2173.435 2712.070 2173.805 ;
        RECT 2711.860 2139.270 2712.000 2173.435 ;
        RECT 2711.800 2138.950 2712.060 2139.270 ;
        RECT 2712.260 2138.610 2712.520 2138.930 ;
        RECT 2712.320 2125.330 2712.460 2138.610 ;
        RECT 2710.880 2125.010 2711.140 2125.330 ;
        RECT 2712.260 2125.010 2712.520 2125.330 ;
        RECT 2710.940 2077.245 2711.080 2125.010 ;
        RECT 2710.870 2076.875 2711.150 2077.245 ;
        RECT 2711.790 2076.875 2712.070 2077.245 ;
        RECT 2711.860 2042.710 2712.000 2076.875 ;
        RECT 2711.800 2042.390 2712.060 2042.710 ;
        RECT 2712.260 2041.710 2712.520 2042.030 ;
        RECT 2712.320 2021.630 2712.460 2041.710 ;
        RECT 2710.420 2021.310 2710.680 2021.630 ;
        RECT 2712.260 2021.310 2712.520 2021.630 ;
        RECT 2710.480 1973.885 2710.620 2021.310 ;
        RECT 2710.410 1973.515 2710.690 1973.885 ;
        RECT 2711.330 1973.770 2711.610 1973.885 ;
        RECT 2711.330 1973.630 2712.000 1973.770 ;
        RECT 2711.330 1973.515 2711.610 1973.630 ;
        RECT 2711.860 1966.550 2712.000 1973.630 ;
        RECT 2710.880 1966.230 2711.140 1966.550 ;
        RECT 2711.800 1966.230 2712.060 1966.550 ;
        RECT 2710.940 1918.610 2711.080 1966.230 ;
        RECT 2710.880 1918.290 2711.140 1918.610 ;
        RECT 2712.260 1918.290 2712.520 1918.610 ;
        RECT 2712.320 1897.530 2712.460 1918.290 ;
        RECT 2712.260 1897.210 2712.520 1897.530 ;
        RECT 2713.180 1897.210 2713.440 1897.530 ;
        RECT 2713.240 1859.530 2713.380 1897.210 ;
        RECT 2713.240 1859.390 2713.840 1859.530 ;
        RECT 2713.700 1835.310 2713.840 1859.390 ;
        RECT 2712.260 1834.990 2712.520 1835.310 ;
        RECT 2713.640 1834.990 2713.900 1835.310 ;
        RECT 2712.320 1787.370 2712.460 1834.990 ;
        RECT 2712.260 1787.050 2712.520 1787.370 ;
        RECT 2712.720 1787.050 2712.980 1787.370 ;
        RECT 2712.780 1753.030 2712.920 1787.050 ;
        RECT 2712.720 1752.710 2712.980 1753.030 ;
        RECT 2713.640 1752.370 2713.900 1752.690 ;
        RECT 2713.700 1704.410 2713.840 1752.370 ;
        RECT 2614.280 1704.090 2614.540 1704.410 ;
        RECT 2713.640 1704.090 2713.900 1704.410 ;
        RECT 2614.340 1699.845 2614.480 1704.090 ;
        RECT 2614.270 1699.475 2614.550 1699.845 ;
      LAYER via2 ;
        RECT 2712.250 3421.960 2712.530 3422.240 ;
        RECT 2712.710 3394.080 2712.990 3394.360 ;
        RECT 2712.710 2608.000 2712.990 2608.280 ;
        RECT 2713.630 2608.000 2713.910 2608.280 ;
        RECT 2713.170 2463.840 2713.450 2464.120 ;
        RECT 2712.710 2463.160 2712.990 2463.440 ;
        RECT 2711.790 2270.040 2712.070 2270.320 ;
        RECT 2713.170 2270.040 2713.450 2270.320 ;
        RECT 2710.870 2173.480 2711.150 2173.760 ;
        RECT 2711.790 2173.480 2712.070 2173.760 ;
        RECT 2710.870 2076.920 2711.150 2077.200 ;
        RECT 2711.790 2076.920 2712.070 2077.200 ;
        RECT 2710.410 1973.560 2710.690 1973.840 ;
        RECT 2711.330 1973.560 2711.610 1973.840 ;
        RECT 2614.270 1699.520 2614.550 1699.800 ;
      LAYER met3 ;
        RECT 2712.225 3422.260 2712.555 3422.265 ;
        RECT 2712.225 3422.250 2712.810 3422.260 ;
        RECT 2712.225 3421.950 2713.010 3422.250 ;
        RECT 2712.225 3421.940 2712.810 3421.950 ;
        RECT 2712.225 3421.935 2712.555 3421.940 ;
        RECT 2712.685 3394.380 2713.015 3394.385 ;
        RECT 2712.430 3394.370 2713.015 3394.380 ;
        RECT 2712.230 3394.070 2713.015 3394.370 ;
        RECT 2712.430 3394.060 2713.015 3394.070 ;
        RECT 2712.685 3394.055 2713.015 3394.060 ;
        RECT 2712.685 2608.290 2713.015 2608.305 ;
        RECT 2713.605 2608.290 2713.935 2608.305 ;
        RECT 2712.685 2607.990 2713.935 2608.290 ;
        RECT 2712.685 2607.975 2713.015 2607.990 ;
        RECT 2713.605 2607.975 2713.935 2607.990 ;
        RECT 2713.145 2464.130 2713.475 2464.145 ;
        RECT 2712.470 2463.830 2713.475 2464.130 ;
        RECT 2712.470 2463.465 2712.770 2463.830 ;
        RECT 2713.145 2463.815 2713.475 2463.830 ;
        RECT 2712.470 2463.150 2713.015 2463.465 ;
        RECT 2712.685 2463.135 2713.015 2463.150 ;
        RECT 2711.765 2270.330 2712.095 2270.345 ;
        RECT 2713.145 2270.330 2713.475 2270.345 ;
        RECT 2711.765 2270.030 2713.475 2270.330 ;
        RECT 2711.765 2270.015 2712.095 2270.030 ;
        RECT 2713.145 2270.015 2713.475 2270.030 ;
        RECT 2710.845 2173.770 2711.175 2173.785 ;
        RECT 2711.765 2173.770 2712.095 2173.785 ;
        RECT 2710.845 2173.470 2712.095 2173.770 ;
        RECT 2710.845 2173.455 2711.175 2173.470 ;
        RECT 2711.765 2173.455 2712.095 2173.470 ;
        RECT 2710.845 2077.210 2711.175 2077.225 ;
        RECT 2711.765 2077.210 2712.095 2077.225 ;
        RECT 2710.845 2076.910 2712.095 2077.210 ;
        RECT 2710.845 2076.895 2711.175 2076.910 ;
        RECT 2711.765 2076.895 2712.095 2076.910 ;
        RECT 2710.385 1973.850 2710.715 1973.865 ;
        RECT 2711.305 1973.850 2711.635 1973.865 ;
        RECT 2710.385 1973.550 2711.635 1973.850 ;
        RECT 2710.385 1973.535 2710.715 1973.550 ;
        RECT 2711.305 1973.535 2711.635 1973.550 ;
        RECT 2614.245 1699.810 2614.575 1699.825 ;
        RECT 2599.460 1699.760 2614.575 1699.810 ;
        RECT 2596.000 1699.510 2614.575 1699.760 ;
        RECT 2596.000 1699.160 2600.000 1699.510 ;
        RECT 2614.245 1699.495 2614.575 1699.510 ;
      LAYER via3 ;
        RECT 2712.460 3421.940 2712.780 3422.260 ;
        RECT 2712.460 3394.060 2712.780 3394.380 ;
      LAYER met4 ;
        RECT 2712.455 3421.935 2712.785 3422.265 ;
        RECT 2712.470 3394.385 2712.770 3421.935 ;
        RECT 2712.455 3394.055 2712.785 3394.385 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2391.610 3477.420 2391.930 3477.480 ;
        RECT 2392.070 3477.420 2392.390 3477.480 ;
        RECT 2391.610 3477.280 2392.390 3477.420 ;
        RECT 2391.610 3477.220 2391.930 3477.280 ;
        RECT 2392.070 3477.220 2392.390 3477.280 ;
        RECT 2391.610 3429.480 2391.930 3429.540 ;
        RECT 2392.530 3429.480 2392.850 3429.540 ;
        RECT 2391.610 3429.340 2392.850 3429.480 ;
        RECT 2391.610 3429.280 2391.930 3429.340 ;
        RECT 2392.530 3429.280 2392.850 3429.340 ;
        RECT 2391.150 3380.860 2391.470 3380.920 ;
        RECT 2392.070 3380.860 2392.390 3380.920 ;
        RECT 2391.150 3380.720 2392.390 3380.860 ;
        RECT 2391.150 3380.660 2391.470 3380.720 ;
        RECT 2392.070 3380.660 2392.390 3380.720 ;
        RECT 2391.150 3332.920 2391.470 3332.980 ;
        RECT 2392.530 3332.920 2392.850 3332.980 ;
        RECT 2391.150 3332.780 2392.850 3332.920 ;
        RECT 2391.150 3332.720 2391.470 3332.780 ;
        RECT 2392.530 3332.720 2392.850 3332.780 ;
        RECT 2392.990 3298.240 2393.310 3298.300 ;
        RECT 2393.910 3298.240 2394.230 3298.300 ;
        RECT 2392.990 3298.100 2394.230 3298.240 ;
        RECT 2392.990 3298.040 2393.310 3298.100 ;
        RECT 2393.910 3298.040 2394.230 3298.100 ;
        RECT 2392.530 3284.300 2392.850 3284.360 ;
        RECT 2393.910 3284.300 2394.230 3284.360 ;
        RECT 2392.530 3284.160 2394.230 3284.300 ;
        RECT 2392.530 3284.100 2392.850 3284.160 ;
        RECT 2393.910 3284.100 2394.230 3284.160 ;
        RECT 2392.530 3236.360 2392.850 3236.420 ;
        RECT 2393.450 3236.360 2393.770 3236.420 ;
        RECT 2392.530 3236.220 2393.770 3236.360 ;
        RECT 2392.530 3236.160 2392.850 3236.220 ;
        RECT 2393.450 3236.160 2393.770 3236.220 ;
        RECT 2393.450 3202.020 2393.770 3202.080 ;
        RECT 2392.620 3201.880 2393.770 3202.020 ;
        RECT 2392.620 3201.400 2392.760 3201.880 ;
        RECT 2393.450 3201.820 2393.770 3201.880 ;
        RECT 2392.530 3201.140 2392.850 3201.400 ;
        RECT 2392.530 3187.740 2392.850 3187.800 ;
        RECT 2392.990 3187.740 2393.310 3187.800 ;
        RECT 2392.530 3187.600 2393.310 3187.740 ;
        RECT 2392.530 3187.540 2392.850 3187.600 ;
        RECT 2392.990 3187.540 2393.310 3187.600 ;
        RECT 2392.990 3139.800 2393.310 3139.860 ;
        RECT 2393.910 3139.800 2394.230 3139.860 ;
        RECT 2392.990 3139.660 2394.230 3139.800 ;
        RECT 2392.990 3139.600 2393.310 3139.660 ;
        RECT 2393.910 3139.600 2394.230 3139.660 ;
        RECT 2392.530 3091.520 2392.850 3091.580 ;
        RECT 2393.910 3091.520 2394.230 3091.580 ;
        RECT 2392.530 3091.380 2394.230 3091.520 ;
        RECT 2392.530 3091.320 2392.850 3091.380 ;
        RECT 2393.910 3091.320 2394.230 3091.380 ;
        RECT 2392.530 3060.240 2392.850 3060.300 ;
        RECT 2598.150 3060.240 2598.470 3060.300 ;
        RECT 2392.530 3060.100 2598.470 3060.240 ;
        RECT 2392.530 3060.040 2392.850 3060.100 ;
        RECT 2598.150 3060.040 2598.470 3060.100 ;
      LAYER via ;
        RECT 2391.640 3477.220 2391.900 3477.480 ;
        RECT 2392.100 3477.220 2392.360 3477.480 ;
        RECT 2391.640 3429.280 2391.900 3429.540 ;
        RECT 2392.560 3429.280 2392.820 3429.540 ;
        RECT 2391.180 3380.660 2391.440 3380.920 ;
        RECT 2392.100 3380.660 2392.360 3380.920 ;
        RECT 2391.180 3332.720 2391.440 3332.980 ;
        RECT 2392.560 3332.720 2392.820 3332.980 ;
        RECT 2393.020 3298.040 2393.280 3298.300 ;
        RECT 2393.940 3298.040 2394.200 3298.300 ;
        RECT 2392.560 3284.100 2392.820 3284.360 ;
        RECT 2393.940 3284.100 2394.200 3284.360 ;
        RECT 2392.560 3236.160 2392.820 3236.420 ;
        RECT 2393.480 3236.160 2393.740 3236.420 ;
        RECT 2393.480 3201.820 2393.740 3202.080 ;
        RECT 2392.560 3201.140 2392.820 3201.400 ;
        RECT 2392.560 3187.540 2392.820 3187.800 ;
        RECT 2393.020 3187.540 2393.280 3187.800 ;
        RECT 2393.020 3139.600 2393.280 3139.860 ;
        RECT 2393.940 3139.600 2394.200 3139.860 ;
        RECT 2392.560 3091.320 2392.820 3091.580 ;
        RECT 2393.940 3091.320 2394.200 3091.580 ;
        RECT 2392.560 3060.040 2392.820 3060.300 ;
        RECT 2598.180 3060.040 2598.440 3060.300 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3517.370 2392.760 3517.600 ;
        RECT 2392.160 3517.230 2392.760 3517.370 ;
        RECT 2392.160 3477.510 2392.300 3517.230 ;
        RECT 2391.640 3477.190 2391.900 3477.510 ;
        RECT 2392.100 3477.190 2392.360 3477.510 ;
        RECT 2391.700 3429.570 2391.840 3477.190 ;
        RECT 2391.640 3429.250 2391.900 3429.570 ;
        RECT 2392.560 3429.250 2392.820 3429.570 ;
        RECT 2392.620 3395.765 2392.760 3429.250 ;
        RECT 2392.550 3395.395 2392.830 3395.765 ;
        RECT 2392.090 3381.115 2392.370 3381.485 ;
        RECT 2392.160 3380.950 2392.300 3381.115 ;
        RECT 2391.180 3380.630 2391.440 3380.950 ;
        RECT 2392.100 3380.630 2392.360 3380.950 ;
        RECT 2391.240 3333.010 2391.380 3380.630 ;
        RECT 2391.180 3332.690 2391.440 3333.010 ;
        RECT 2392.560 3332.690 2392.820 3333.010 ;
        RECT 2392.620 3298.410 2392.760 3332.690 ;
        RECT 2392.620 3298.330 2393.220 3298.410 ;
        RECT 2392.620 3298.270 2393.280 3298.330 ;
        RECT 2393.020 3298.010 2393.280 3298.270 ;
        RECT 2393.940 3298.010 2394.200 3298.330 ;
        RECT 2394.000 3284.390 2394.140 3298.010 ;
        RECT 2392.560 3284.070 2392.820 3284.390 ;
        RECT 2393.940 3284.070 2394.200 3284.390 ;
        RECT 2392.620 3236.450 2392.760 3284.070 ;
        RECT 2392.560 3236.130 2392.820 3236.450 ;
        RECT 2393.480 3236.130 2393.740 3236.450 ;
        RECT 2393.540 3202.110 2393.680 3236.130 ;
        RECT 2393.480 3201.790 2393.740 3202.110 ;
        RECT 2392.560 3201.110 2392.820 3201.430 ;
        RECT 2392.620 3187.830 2392.760 3201.110 ;
        RECT 2392.560 3187.510 2392.820 3187.830 ;
        RECT 2393.020 3187.510 2393.280 3187.830 ;
        RECT 2393.080 3139.890 2393.220 3187.510 ;
        RECT 2393.020 3139.570 2393.280 3139.890 ;
        RECT 2393.940 3139.570 2394.200 3139.890 ;
        RECT 2394.000 3091.610 2394.140 3139.570 ;
        RECT 2392.560 3091.290 2392.820 3091.610 ;
        RECT 2393.940 3091.290 2394.200 3091.610 ;
        RECT 2392.620 3060.330 2392.760 3091.290 ;
        RECT 2392.560 3060.010 2392.820 3060.330 ;
        RECT 2598.180 3060.010 2598.440 3060.330 ;
        RECT 2598.240 1732.485 2598.380 3060.010 ;
        RECT 2598.170 1732.115 2598.450 1732.485 ;
      LAYER via2 ;
        RECT 2392.550 3395.440 2392.830 3395.720 ;
        RECT 2392.090 3381.160 2392.370 3381.440 ;
        RECT 2598.170 1732.160 2598.450 1732.440 ;
      LAYER met3 ;
        RECT 2392.525 3395.740 2392.855 3395.745 ;
        RECT 2392.270 3395.730 2392.855 3395.740 ;
        RECT 2392.070 3395.430 2392.855 3395.730 ;
        RECT 2392.270 3395.420 2392.855 3395.430 ;
        RECT 2392.525 3395.415 2392.855 3395.420 ;
        RECT 2392.065 3381.460 2392.395 3381.465 ;
        RECT 2392.065 3381.450 2392.650 3381.460 ;
        RECT 2392.065 3381.150 2392.850 3381.450 ;
        RECT 2392.065 3381.140 2392.650 3381.150 ;
        RECT 2392.065 3381.135 2392.395 3381.140 ;
        RECT 2598.145 1732.450 2598.475 1732.465 ;
        RECT 2598.145 1732.135 2598.690 1732.450 ;
        RECT 2598.390 1731.720 2598.690 1732.135 ;
        RECT 2596.000 1731.120 2600.000 1731.720 ;
      LAYER via3 ;
        RECT 2392.300 3395.420 2392.620 3395.740 ;
        RECT 2392.300 3381.140 2392.620 3381.460 ;
      LAYER met4 ;
        RECT 2392.295 3395.415 2392.625 3395.745 ;
        RECT 2392.310 3381.465 2392.610 3395.415 ;
        RECT 2392.295 3381.135 2392.625 3381.465 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2067.770 3477.760 2068.090 3477.820 ;
        RECT 2068.230 3477.760 2068.550 3477.820 ;
        RECT 2067.770 3477.620 2068.550 3477.760 ;
        RECT 2067.770 3477.560 2068.090 3477.620 ;
        RECT 2068.230 3477.560 2068.550 3477.620 ;
        RECT 2068.230 3443.080 2068.550 3443.140 ;
        RECT 2069.150 3443.080 2069.470 3443.140 ;
        RECT 2068.230 3442.940 2069.470 3443.080 ;
        RECT 2068.230 3442.880 2068.550 3442.940 ;
        RECT 2069.150 3442.880 2069.470 3442.940 ;
        RECT 2067.770 3429.140 2068.090 3429.200 ;
        RECT 2069.150 3429.140 2069.470 3429.200 ;
        RECT 2067.770 3429.000 2069.470 3429.140 ;
        RECT 2067.770 3428.940 2068.090 3429.000 ;
        RECT 2069.150 3428.940 2069.470 3429.000 ;
        RECT 2067.770 3381.200 2068.090 3381.260 ;
        RECT 2068.690 3381.200 2069.010 3381.260 ;
        RECT 2067.770 3381.060 2069.010 3381.200 ;
        RECT 2067.770 3381.000 2068.090 3381.060 ;
        RECT 2068.690 3381.000 2069.010 3381.060 ;
        RECT 2068.690 3367.600 2069.010 3367.660 ;
        RECT 2069.610 3367.600 2069.930 3367.660 ;
        RECT 2068.690 3367.460 2069.930 3367.600 ;
        RECT 2068.690 3367.400 2069.010 3367.460 ;
        RECT 2069.610 3367.400 2069.930 3367.460 ;
        RECT 2068.690 3270.700 2069.010 3270.760 ;
        RECT 2069.610 3270.700 2069.930 3270.760 ;
        RECT 2068.690 3270.560 2069.930 3270.700 ;
        RECT 2068.690 3270.500 2069.010 3270.560 ;
        RECT 2069.610 3270.500 2069.930 3270.560 ;
        RECT 2068.690 3174.140 2069.010 3174.200 ;
        RECT 2069.610 3174.140 2069.930 3174.200 ;
        RECT 2068.690 3174.000 2069.930 3174.140 ;
        RECT 2068.690 3173.940 2069.010 3174.000 ;
        RECT 2069.610 3173.940 2069.930 3174.000 ;
        RECT 2068.690 3077.580 2069.010 3077.640 ;
        RECT 2069.610 3077.580 2069.930 3077.640 ;
        RECT 2068.690 3077.440 2069.930 3077.580 ;
        RECT 2068.690 3077.380 2069.010 3077.440 ;
        RECT 2069.610 3077.380 2069.930 3077.440 ;
        RECT 2067.310 2994.620 2067.630 2994.680 ;
        RECT 2068.690 2994.620 2069.010 2994.680 ;
        RECT 2067.310 2994.480 2069.010 2994.620 ;
        RECT 2067.310 2994.420 2067.630 2994.480 ;
        RECT 2068.690 2994.420 2069.010 2994.480 ;
        RECT 2067.310 2946.340 2067.630 2946.400 ;
        RECT 2067.770 2946.340 2068.090 2946.400 ;
        RECT 2067.310 2946.200 2068.090 2946.340 ;
        RECT 2067.310 2946.140 2067.630 2946.200 ;
        RECT 2067.770 2946.140 2068.090 2946.200 ;
        RECT 2067.310 2911.320 2067.630 2911.380 ;
        RECT 2068.690 2911.320 2069.010 2911.380 ;
        RECT 2067.310 2911.180 2069.010 2911.320 ;
        RECT 2067.310 2911.120 2067.630 2911.180 ;
        RECT 2068.690 2911.120 2069.010 2911.180 ;
        RECT 2067.310 2898.060 2067.630 2898.120 ;
        RECT 2068.690 2898.060 2069.010 2898.120 ;
        RECT 2067.310 2897.920 2069.010 2898.060 ;
        RECT 2067.310 2897.860 2067.630 2897.920 ;
        RECT 2068.690 2897.860 2069.010 2897.920 ;
        RECT 2067.310 2849.780 2067.630 2849.840 ;
        RECT 2068.230 2849.780 2068.550 2849.840 ;
        RECT 2067.310 2849.640 2068.550 2849.780 ;
        RECT 2067.310 2849.580 2067.630 2849.640 ;
        RECT 2068.230 2849.580 2068.550 2849.640 ;
        RECT 2068.230 2815.240 2068.550 2815.500 ;
        RECT 2068.320 2814.760 2068.460 2815.240 ;
        RECT 2068.690 2814.760 2069.010 2814.820 ;
        RECT 2068.320 2814.620 2069.010 2814.760 ;
        RECT 2068.690 2814.560 2069.010 2814.620 ;
        RECT 2068.230 2767.160 2068.550 2767.220 ;
        RECT 2068.230 2767.020 2068.920 2767.160 ;
        RECT 2068.230 2766.960 2068.550 2767.020 ;
        RECT 2068.780 2766.880 2068.920 2767.020 ;
        RECT 2068.690 2766.620 2069.010 2766.880 ;
        RECT 2068.230 2753.220 2068.550 2753.280 ;
        RECT 2068.690 2753.220 2069.010 2753.280 ;
        RECT 2068.230 2753.080 2069.010 2753.220 ;
        RECT 2068.230 2753.020 2068.550 2753.080 ;
        RECT 2068.690 2753.020 2069.010 2753.080 ;
        RECT 2068.230 2718.680 2068.550 2718.940 ;
        RECT 2068.320 2718.200 2068.460 2718.680 ;
        RECT 2068.690 2718.200 2069.010 2718.260 ;
        RECT 2068.320 2718.060 2069.010 2718.200 ;
        RECT 2068.690 2718.000 2069.010 2718.060 ;
        RECT 2068.230 2670.600 2068.550 2670.660 ;
        RECT 2068.230 2670.460 2068.920 2670.600 ;
        RECT 2068.230 2670.400 2068.550 2670.460 ;
        RECT 2068.780 2670.320 2068.920 2670.460 ;
        RECT 2068.690 2670.060 2069.010 2670.320 ;
        RECT 2068.230 2656.660 2068.550 2656.720 ;
        RECT 2068.690 2656.660 2069.010 2656.720 ;
        RECT 2068.230 2656.520 2069.010 2656.660 ;
        RECT 2068.230 2656.460 2068.550 2656.520 ;
        RECT 2068.690 2656.460 2069.010 2656.520 ;
        RECT 2068.230 2622.120 2068.550 2622.380 ;
        RECT 2068.320 2621.640 2068.460 2622.120 ;
        RECT 2068.690 2621.640 2069.010 2621.700 ;
        RECT 2068.320 2621.500 2069.010 2621.640 ;
        RECT 2068.690 2621.440 2069.010 2621.500 ;
        RECT 2067.770 2560.100 2068.090 2560.160 ;
        RECT 2069.150 2560.100 2069.470 2560.160 ;
        RECT 2067.770 2559.960 2069.470 2560.100 ;
        RECT 2067.770 2559.900 2068.090 2559.960 ;
        RECT 2069.150 2559.900 2069.470 2559.960 ;
        RECT 2069.150 2525.560 2069.470 2525.820 ;
        RECT 2069.240 2525.080 2069.380 2525.560 ;
        RECT 2069.610 2525.080 2069.930 2525.140 ;
        RECT 2069.240 2524.940 2069.930 2525.080 ;
        RECT 2069.610 2524.880 2069.930 2524.940 ;
        RECT 2067.770 2463.200 2068.090 2463.260 ;
        RECT 2069.150 2463.200 2069.470 2463.260 ;
        RECT 2067.770 2463.060 2069.470 2463.200 ;
        RECT 2067.770 2463.000 2068.090 2463.060 ;
        RECT 2069.150 2463.000 2069.470 2463.060 ;
        RECT 2068.690 2405.060 2069.010 2405.120 ;
        RECT 2600.450 2405.060 2600.770 2405.120 ;
        RECT 2068.690 2404.920 2600.770 2405.060 ;
        RECT 2068.690 2404.860 2069.010 2404.920 ;
        RECT 2600.450 2404.860 2600.770 2404.920 ;
        RECT 2600.450 2381.260 2600.770 2381.320 ;
        RECT 2599.620 2381.120 2600.770 2381.260 ;
        RECT 2599.620 2380.640 2599.760 2381.120 ;
        RECT 2600.450 2381.060 2600.770 2381.120 ;
        RECT 2599.530 2380.380 2599.850 2380.640 ;
      LAYER via ;
        RECT 2067.800 3477.560 2068.060 3477.820 ;
        RECT 2068.260 3477.560 2068.520 3477.820 ;
        RECT 2068.260 3442.880 2068.520 3443.140 ;
        RECT 2069.180 3442.880 2069.440 3443.140 ;
        RECT 2067.800 3428.940 2068.060 3429.200 ;
        RECT 2069.180 3428.940 2069.440 3429.200 ;
        RECT 2067.800 3381.000 2068.060 3381.260 ;
        RECT 2068.720 3381.000 2068.980 3381.260 ;
        RECT 2068.720 3367.400 2068.980 3367.660 ;
        RECT 2069.640 3367.400 2069.900 3367.660 ;
        RECT 2068.720 3270.500 2068.980 3270.760 ;
        RECT 2069.640 3270.500 2069.900 3270.760 ;
        RECT 2068.720 3173.940 2068.980 3174.200 ;
        RECT 2069.640 3173.940 2069.900 3174.200 ;
        RECT 2068.720 3077.380 2068.980 3077.640 ;
        RECT 2069.640 3077.380 2069.900 3077.640 ;
        RECT 2067.340 2994.420 2067.600 2994.680 ;
        RECT 2068.720 2994.420 2068.980 2994.680 ;
        RECT 2067.340 2946.140 2067.600 2946.400 ;
        RECT 2067.800 2946.140 2068.060 2946.400 ;
        RECT 2067.340 2911.120 2067.600 2911.380 ;
        RECT 2068.720 2911.120 2068.980 2911.380 ;
        RECT 2067.340 2897.860 2067.600 2898.120 ;
        RECT 2068.720 2897.860 2068.980 2898.120 ;
        RECT 2067.340 2849.580 2067.600 2849.840 ;
        RECT 2068.260 2849.580 2068.520 2849.840 ;
        RECT 2068.260 2815.240 2068.520 2815.500 ;
        RECT 2068.720 2814.560 2068.980 2814.820 ;
        RECT 2068.260 2766.960 2068.520 2767.220 ;
        RECT 2068.720 2766.620 2068.980 2766.880 ;
        RECT 2068.260 2753.020 2068.520 2753.280 ;
        RECT 2068.720 2753.020 2068.980 2753.280 ;
        RECT 2068.260 2718.680 2068.520 2718.940 ;
        RECT 2068.720 2718.000 2068.980 2718.260 ;
        RECT 2068.260 2670.400 2068.520 2670.660 ;
        RECT 2068.720 2670.060 2068.980 2670.320 ;
        RECT 2068.260 2656.460 2068.520 2656.720 ;
        RECT 2068.720 2656.460 2068.980 2656.720 ;
        RECT 2068.260 2622.120 2068.520 2622.380 ;
        RECT 2068.720 2621.440 2068.980 2621.700 ;
        RECT 2067.800 2559.900 2068.060 2560.160 ;
        RECT 2069.180 2559.900 2069.440 2560.160 ;
        RECT 2069.180 2525.560 2069.440 2525.820 ;
        RECT 2069.640 2524.880 2069.900 2525.140 ;
        RECT 2067.800 2463.000 2068.060 2463.260 ;
        RECT 2069.180 2463.000 2069.440 2463.260 ;
        RECT 2068.720 2404.860 2068.980 2405.120 ;
        RECT 2600.480 2404.860 2600.740 2405.120 ;
        RECT 2600.480 2381.060 2600.740 2381.320 ;
        RECT 2599.560 2380.380 2599.820 2380.640 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3517.370 2068.460 3517.600 ;
        RECT 2067.860 3517.230 2068.460 3517.370 ;
        RECT 2067.860 3477.850 2068.000 3517.230 ;
        RECT 2067.800 3477.530 2068.060 3477.850 ;
        RECT 2068.260 3477.530 2068.520 3477.850 ;
        RECT 2068.320 3443.170 2068.460 3477.530 ;
        RECT 2068.260 3442.850 2068.520 3443.170 ;
        RECT 2069.180 3442.850 2069.440 3443.170 ;
        RECT 2069.240 3429.230 2069.380 3442.850 ;
        RECT 2067.800 3428.910 2068.060 3429.230 ;
        RECT 2069.180 3428.910 2069.440 3429.230 ;
        RECT 2067.860 3381.290 2068.000 3428.910 ;
        RECT 2067.800 3380.970 2068.060 3381.290 ;
        RECT 2068.720 3380.970 2068.980 3381.290 ;
        RECT 2068.780 3367.690 2068.920 3380.970 ;
        RECT 2068.720 3367.370 2068.980 3367.690 ;
        RECT 2069.640 3367.370 2069.900 3367.690 ;
        RECT 2069.700 3318.810 2069.840 3367.370 ;
        RECT 2068.780 3318.670 2069.840 3318.810 ;
        RECT 2068.780 3270.790 2068.920 3318.670 ;
        RECT 2068.720 3270.470 2068.980 3270.790 ;
        RECT 2069.640 3270.470 2069.900 3270.790 ;
        RECT 2069.700 3222.250 2069.840 3270.470 ;
        RECT 2068.780 3222.110 2069.840 3222.250 ;
        RECT 2068.780 3174.230 2068.920 3222.110 ;
        RECT 2068.720 3173.910 2068.980 3174.230 ;
        RECT 2069.640 3173.910 2069.900 3174.230 ;
        RECT 2069.700 3125.690 2069.840 3173.910 ;
        RECT 2068.780 3125.550 2069.840 3125.690 ;
        RECT 2068.780 3077.670 2068.920 3125.550 ;
        RECT 2068.720 3077.410 2068.980 3077.670 ;
        RECT 2069.640 3077.410 2069.900 3077.670 ;
        RECT 2068.720 3077.350 2069.900 3077.410 ;
        RECT 2068.780 3077.270 2069.840 3077.350 ;
        RECT 2068.780 2994.710 2068.920 3077.270 ;
        RECT 2067.340 2994.390 2067.600 2994.710 ;
        RECT 2068.720 2994.390 2068.980 2994.710 ;
        RECT 2067.400 2946.850 2067.540 2994.390 ;
        RECT 2067.400 2946.710 2068.000 2946.850 ;
        RECT 2067.860 2946.430 2068.000 2946.710 ;
        RECT 2067.340 2946.110 2067.600 2946.430 ;
        RECT 2067.800 2946.110 2068.060 2946.430 ;
        RECT 2067.400 2911.410 2067.540 2946.110 ;
        RECT 2067.340 2911.090 2067.600 2911.410 ;
        RECT 2068.720 2911.090 2068.980 2911.410 ;
        RECT 2068.780 2898.150 2068.920 2911.090 ;
        RECT 2067.340 2897.830 2067.600 2898.150 ;
        RECT 2068.720 2897.830 2068.980 2898.150 ;
        RECT 2067.400 2849.870 2067.540 2897.830 ;
        RECT 2067.340 2849.550 2067.600 2849.870 ;
        RECT 2068.260 2849.550 2068.520 2849.870 ;
        RECT 2068.320 2815.530 2068.460 2849.550 ;
        RECT 2068.260 2815.210 2068.520 2815.530 ;
        RECT 2068.720 2814.530 2068.980 2814.850 ;
        RECT 2068.780 2801.330 2068.920 2814.530 ;
        RECT 2068.320 2801.190 2068.920 2801.330 ;
        RECT 2068.320 2767.250 2068.460 2801.190 ;
        RECT 2068.260 2766.930 2068.520 2767.250 ;
        RECT 2068.720 2766.590 2068.980 2766.910 ;
        RECT 2068.780 2753.310 2068.920 2766.590 ;
        RECT 2068.260 2752.990 2068.520 2753.310 ;
        RECT 2068.720 2752.990 2068.980 2753.310 ;
        RECT 2068.320 2718.970 2068.460 2752.990 ;
        RECT 2068.260 2718.650 2068.520 2718.970 ;
        RECT 2068.720 2717.970 2068.980 2718.290 ;
        RECT 2068.780 2704.770 2068.920 2717.970 ;
        RECT 2068.320 2704.630 2068.920 2704.770 ;
        RECT 2068.320 2670.690 2068.460 2704.630 ;
        RECT 2068.260 2670.370 2068.520 2670.690 ;
        RECT 2068.720 2670.030 2068.980 2670.350 ;
        RECT 2068.780 2656.750 2068.920 2670.030 ;
        RECT 2068.260 2656.430 2068.520 2656.750 ;
        RECT 2068.720 2656.430 2068.980 2656.750 ;
        RECT 2068.320 2622.410 2068.460 2656.430 ;
        RECT 2068.260 2622.090 2068.520 2622.410 ;
        RECT 2068.720 2621.410 2068.980 2621.730 ;
        RECT 2068.780 2608.325 2068.920 2621.410 ;
        RECT 2067.790 2607.955 2068.070 2608.325 ;
        RECT 2068.710 2607.955 2068.990 2608.325 ;
        RECT 2067.860 2560.190 2068.000 2607.955 ;
        RECT 2067.800 2559.870 2068.060 2560.190 ;
        RECT 2069.180 2559.870 2069.440 2560.190 ;
        RECT 2069.240 2525.850 2069.380 2559.870 ;
        RECT 2069.180 2525.530 2069.440 2525.850 ;
        RECT 2069.640 2524.850 2069.900 2525.170 ;
        RECT 2069.700 2476.970 2069.840 2524.850 ;
        RECT 2069.240 2476.830 2069.840 2476.970 ;
        RECT 2069.240 2463.290 2069.380 2476.830 ;
        RECT 2067.800 2462.970 2068.060 2463.290 ;
        RECT 2069.180 2462.970 2069.440 2463.290 ;
        RECT 2067.860 2415.205 2068.000 2462.970 ;
        RECT 2067.790 2414.835 2068.070 2415.205 ;
        RECT 2068.710 2414.835 2068.990 2415.205 ;
        RECT 2068.780 2405.150 2068.920 2414.835 ;
        RECT 2068.720 2404.830 2068.980 2405.150 ;
        RECT 2600.480 2404.830 2600.740 2405.150 ;
        RECT 2600.540 2381.350 2600.680 2404.830 ;
        RECT 2600.480 2381.030 2600.740 2381.350 ;
        RECT 2599.560 2380.350 2599.820 2380.670 ;
        RECT 2599.620 1765.805 2599.760 2380.350 ;
        RECT 2599.550 1765.435 2599.830 1765.805 ;
      LAYER via2 ;
        RECT 2067.790 2608.000 2068.070 2608.280 ;
        RECT 2068.710 2608.000 2068.990 2608.280 ;
        RECT 2067.790 2414.880 2068.070 2415.160 ;
        RECT 2068.710 2414.880 2068.990 2415.160 ;
        RECT 2599.550 1765.480 2599.830 1765.760 ;
      LAYER met3 ;
        RECT 2067.765 2608.290 2068.095 2608.305 ;
        RECT 2068.685 2608.290 2069.015 2608.305 ;
        RECT 2067.765 2607.990 2069.015 2608.290 ;
        RECT 2067.765 2607.975 2068.095 2607.990 ;
        RECT 2068.685 2607.975 2069.015 2607.990 ;
        RECT 2067.765 2415.170 2068.095 2415.185 ;
        RECT 2068.685 2415.170 2069.015 2415.185 ;
        RECT 2067.765 2414.870 2069.015 2415.170 ;
        RECT 2067.765 2414.855 2068.095 2414.870 ;
        RECT 2068.685 2414.855 2069.015 2414.870 ;
        RECT 2599.525 1765.770 2599.855 1765.785 ;
        RECT 2599.310 1765.455 2599.855 1765.770 ;
        RECT 2599.310 1763.000 2599.610 1765.455 ;
        RECT 2596.000 1762.400 2600.000 1763.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1743.930 3503.940 1744.250 3504.000 ;
        RECT 2601.370 3503.940 2601.690 3504.000 ;
        RECT 1743.930 3503.800 2601.690 3503.940 ;
        RECT 1743.930 3503.740 1744.250 3503.800 ;
        RECT 2601.370 3503.740 2601.690 3503.800 ;
      LAYER via ;
        RECT 1743.960 3503.740 1744.220 3504.000 ;
        RECT 2601.400 3503.740 2601.660 3504.000 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3504.030 1744.160 3517.600 ;
        RECT 1743.960 3503.710 1744.220 3504.030 ;
        RECT 2601.400 3503.710 2601.660 3504.030 ;
        RECT 2601.460 1795.045 2601.600 3503.710 ;
        RECT 2601.390 1794.675 2601.670 1795.045 ;
      LAYER via2 ;
        RECT 2601.390 1794.720 2601.670 1795.000 ;
      LAYER met3 ;
        RECT 2601.365 1795.010 2601.695 1795.025 ;
        RECT 2599.460 1794.960 2601.695 1795.010 ;
        RECT 2596.000 1794.710 2601.695 1794.960 ;
        RECT 2596.000 1794.360 2600.000 1794.710 ;
        RECT 2601.365 1794.695 2601.695 1794.710 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3503.260 1419.490 3503.320 ;
        RECT 2601.830 3503.260 2602.150 3503.320 ;
        RECT 1419.170 3503.120 2602.150 3503.260 ;
        RECT 1419.170 3503.060 1419.490 3503.120 ;
        RECT 2601.830 3503.060 2602.150 3503.120 ;
      LAYER via ;
        RECT 1419.200 3503.060 1419.460 3503.320 ;
        RECT 2601.860 3503.060 2602.120 3503.320 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3503.350 1419.400 3517.600 ;
        RECT 1419.200 3503.030 1419.460 3503.350 ;
        RECT 2601.860 3503.030 2602.120 3503.350 ;
        RECT 2601.920 1826.325 2602.060 3503.030 ;
        RECT 2601.850 1825.955 2602.130 1826.325 ;
      LAYER via2 ;
        RECT 2601.850 1826.000 2602.130 1826.280 ;
      LAYER met3 ;
        RECT 2601.825 1826.290 2602.155 1826.305 ;
        RECT 2599.460 1826.240 2602.155 1826.290 ;
        RECT 2596.000 1825.990 2602.155 1826.240 ;
        RECT 2596.000 1825.640 2600.000 1825.990 ;
        RECT 2601.825 1825.975 2602.155 1825.990 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2612.870 386.140 2613.190 386.200 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 2612.870 386.000 2901.150 386.140 ;
        RECT 2612.870 385.940 2613.190 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
      LAYER via ;
        RECT 2612.900 385.940 2613.160 386.200 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
      LAYER met2 ;
        RECT 2612.890 1257.475 2613.170 1257.845 ;
        RECT 2612.960 386.230 2613.100 1257.475 ;
        RECT 2612.900 385.910 2613.160 386.230 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 2612.890 1257.520 2613.170 1257.800 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 2612.865 1257.810 2613.195 1257.825 ;
        RECT 2599.460 1257.760 2613.195 1257.810 ;
        RECT 2596.000 1257.510 2613.195 1257.760 ;
        RECT 2596.000 1257.160 2600.000 1257.510 ;
        RECT 2612.865 1257.495 2613.195 1257.510 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3502.580 1095.190 3502.640 ;
        RECT 2596.770 3502.580 2597.090 3502.640 ;
        RECT 1094.870 3502.440 2597.090 3502.580 ;
        RECT 1094.870 3502.380 1095.190 3502.440 ;
        RECT 2596.770 3502.380 2597.090 3502.440 ;
        RECT 2596.770 2404.720 2597.090 2404.780 ;
        RECT 2600.910 2404.720 2601.230 2404.780 ;
        RECT 2596.770 2404.580 2601.230 2404.720 ;
        RECT 2596.770 2404.520 2597.090 2404.580 ;
        RECT 2600.910 2404.520 2601.230 2404.580 ;
        RECT 2600.910 2380.040 2601.230 2380.300 ;
        RECT 2596.770 2379.900 2597.090 2379.960 ;
        RECT 2601.000 2379.900 2601.140 2380.040 ;
        RECT 2596.770 2379.760 2601.140 2379.900 ;
        RECT 2596.770 2379.700 2597.090 2379.760 ;
        RECT 2596.770 2332.640 2597.090 2332.700 ;
        RECT 2602.290 2332.640 2602.610 2332.700 ;
        RECT 2596.770 2332.500 2602.610 2332.640 ;
        RECT 2596.770 2332.440 2597.090 2332.500 ;
        RECT 2602.290 2332.440 2602.610 2332.500 ;
        RECT 2596.770 2331.960 2597.090 2332.020 ;
        RECT 2602.290 2331.960 2602.610 2332.020 ;
        RECT 2596.770 2331.820 2602.610 2331.960 ;
        RECT 2596.770 2331.760 2597.090 2331.820 ;
        RECT 2602.290 2331.760 2602.610 2331.820 ;
        RECT 2596.770 2285.040 2597.090 2285.100 ;
        RECT 2602.290 2285.040 2602.610 2285.100 ;
        RECT 2596.770 2284.900 2602.610 2285.040 ;
        RECT 2596.770 2284.840 2597.090 2284.900 ;
        RECT 2602.290 2284.840 2602.610 2284.900 ;
      LAYER via ;
        RECT 1094.900 3502.380 1095.160 3502.640 ;
        RECT 2596.800 3502.380 2597.060 3502.640 ;
        RECT 2596.800 2404.520 2597.060 2404.780 ;
        RECT 2600.940 2404.520 2601.200 2404.780 ;
        RECT 2600.940 2380.040 2601.200 2380.300 ;
        RECT 2596.800 2379.700 2597.060 2379.960 ;
        RECT 2596.800 2332.440 2597.060 2332.700 ;
        RECT 2602.320 2332.440 2602.580 2332.700 ;
        RECT 2596.800 2331.760 2597.060 2332.020 ;
        RECT 2602.320 2331.760 2602.580 2332.020 ;
        RECT 2596.800 2284.840 2597.060 2285.100 ;
        RECT 2602.320 2284.840 2602.580 2285.100 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3502.670 1095.100 3517.600 ;
        RECT 1094.900 3502.350 1095.160 3502.670 ;
        RECT 2596.800 3502.350 2597.060 3502.670 ;
        RECT 2596.860 2404.810 2597.000 3502.350 ;
        RECT 2596.800 2404.490 2597.060 2404.810 ;
        RECT 2600.940 2404.490 2601.200 2404.810 ;
        RECT 2601.000 2380.330 2601.140 2404.490 ;
        RECT 2600.940 2380.010 2601.200 2380.330 ;
        RECT 2596.800 2379.670 2597.060 2379.990 ;
        RECT 2596.860 2332.730 2597.000 2379.670 ;
        RECT 2596.800 2332.410 2597.060 2332.730 ;
        RECT 2602.320 2332.410 2602.580 2332.730 ;
        RECT 2602.380 2332.050 2602.520 2332.410 ;
        RECT 2596.800 2331.730 2597.060 2332.050 ;
        RECT 2602.320 2331.730 2602.580 2332.050 ;
        RECT 2596.860 2285.130 2597.000 2331.730 ;
        RECT 2596.800 2284.810 2597.060 2285.130 ;
        RECT 2602.320 2284.810 2602.580 2285.130 ;
        RECT 2602.380 2185.365 2602.520 2284.810 ;
        RECT 2602.310 2184.995 2602.590 2185.365 ;
        RECT 2596.790 2161.195 2597.070 2161.565 ;
        RECT 2596.860 1860.325 2597.000 2161.195 ;
        RECT 2596.790 1859.955 2597.070 1860.325 ;
      LAYER via2 ;
        RECT 2602.310 2185.040 2602.590 2185.320 ;
        RECT 2596.790 2161.240 2597.070 2161.520 ;
        RECT 2596.790 1860.000 2597.070 1860.280 ;
      LAYER met3 ;
        RECT 2600.190 2185.330 2600.570 2185.340 ;
        RECT 2602.285 2185.330 2602.615 2185.345 ;
        RECT 2600.190 2185.030 2602.615 2185.330 ;
        RECT 2600.190 2185.020 2600.570 2185.030 ;
        RECT 2602.285 2185.015 2602.615 2185.030 ;
        RECT 2596.765 2161.530 2597.095 2161.545 ;
        RECT 2600.190 2161.530 2600.570 2161.540 ;
        RECT 2596.765 2161.230 2600.570 2161.530 ;
        RECT 2596.765 2161.215 2597.095 2161.230 ;
        RECT 2600.190 2161.220 2600.570 2161.230 ;
        RECT 2596.765 1860.290 2597.095 1860.305 ;
        RECT 2596.550 1859.975 2597.095 1860.290 ;
        RECT 2596.550 1857.520 2596.850 1859.975 ;
        RECT 2596.000 1856.920 2600.000 1857.520 ;
      LAYER via3 ;
        RECT 2600.220 2185.020 2600.540 2185.340 ;
        RECT 2600.220 2161.220 2600.540 2161.540 ;
      LAYER met4 ;
        RECT 2600.215 2185.015 2600.545 2185.345 ;
        RECT 2600.230 2161.545 2600.530 2185.015 ;
        RECT 2600.215 2161.215 2600.545 2161.545 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3501.900 770.890 3501.960 ;
        RECT 2602.290 3501.900 2602.610 3501.960 ;
        RECT 770.570 3501.760 2602.610 3501.900 ;
        RECT 770.570 3501.700 770.890 3501.760 ;
        RECT 2602.290 3501.700 2602.610 3501.760 ;
        RECT 2602.290 2356.440 2602.610 2356.500 ;
        RECT 2604.130 2356.440 2604.450 2356.500 ;
        RECT 2602.290 2356.300 2604.450 2356.440 ;
        RECT 2602.290 2356.240 2602.610 2356.300 ;
        RECT 2604.130 2356.240 2604.450 2356.300 ;
        RECT 2602.290 2184.740 2602.610 2184.800 ;
        RECT 2604.130 2184.740 2604.450 2184.800 ;
        RECT 2602.290 2184.600 2604.450 2184.740 ;
        RECT 2602.290 2184.540 2602.610 2184.600 ;
        RECT 2604.130 2184.540 2604.450 2184.600 ;
      LAYER via ;
        RECT 770.600 3501.700 770.860 3501.960 ;
        RECT 2602.320 3501.700 2602.580 3501.960 ;
        RECT 2602.320 2356.240 2602.580 2356.500 ;
        RECT 2604.160 2356.240 2604.420 2356.500 ;
        RECT 2602.320 2184.540 2602.580 2184.800 ;
        RECT 2604.160 2184.540 2604.420 2184.800 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3501.990 770.800 3517.600 ;
        RECT 770.600 3501.670 770.860 3501.990 ;
        RECT 2602.320 3501.670 2602.580 3501.990 ;
        RECT 2602.380 2356.530 2602.520 3501.670 ;
        RECT 2602.320 2356.210 2602.580 2356.530 ;
        RECT 2604.160 2356.210 2604.420 2356.530 ;
        RECT 2604.220 2184.830 2604.360 2356.210 ;
        RECT 2602.320 2184.510 2602.580 2184.830 ;
        RECT 2604.160 2184.510 2604.420 2184.830 ;
        RECT 2602.380 1889.565 2602.520 2184.510 ;
        RECT 2602.310 1889.195 2602.590 1889.565 ;
      LAYER via2 ;
        RECT 2602.310 1889.240 2602.590 1889.520 ;
      LAYER met3 ;
        RECT 2602.285 1889.530 2602.615 1889.545 ;
        RECT 2599.460 1889.480 2602.615 1889.530 ;
        RECT 2596.000 1889.230 2602.615 1889.480 ;
        RECT 2596.000 1888.880 2600.000 1889.230 ;
        RECT 2602.285 1889.215 2602.615 1889.230 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3503.885 446.040 3517.600 ;
        RECT 445.830 3503.515 446.110 3503.885 ;
      LAYER via2 ;
        RECT 445.830 3503.560 446.110 3503.840 ;
      LAYER met3 ;
        RECT 445.805 3503.850 446.135 3503.865 ;
        RECT 2602.030 3503.850 2602.410 3503.860 ;
        RECT 445.805 3503.550 2602.410 3503.850 ;
        RECT 445.805 3503.535 446.135 3503.550 ;
        RECT 2602.030 3503.540 2602.410 3503.550 ;
        RECT 2602.030 1920.810 2602.410 1920.820 ;
        RECT 2599.460 1920.760 2602.410 1920.810 ;
        RECT 2596.000 1920.510 2602.410 1920.760 ;
        RECT 2596.000 1920.160 2600.000 1920.510 ;
        RECT 2602.030 1920.500 2602.410 1920.510 ;
      LAYER via3 ;
        RECT 2602.060 3503.540 2602.380 3503.860 ;
        RECT 2602.060 1920.500 2602.380 1920.820 ;
      LAYER met4 ;
        RECT 2602.055 3503.535 2602.385 3503.865 ;
        RECT 2602.070 1920.825 2602.370 3503.535 ;
        RECT 2602.055 1920.495 2602.385 1920.825 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3502.525 121.740 3517.600 ;
        RECT 121.530 3502.155 121.810 3502.525 ;
      LAYER via2 ;
        RECT 121.530 3502.200 121.810 3502.480 ;
      LAYER met3 ;
        RECT 121.505 3502.490 121.835 3502.505 ;
        RECT 2602.950 3502.490 2603.330 3502.500 ;
        RECT 121.505 3502.190 2603.330 3502.490 ;
        RECT 121.505 3502.175 121.835 3502.190 ;
        RECT 2602.950 3502.180 2603.330 3502.190 ;
        RECT 2602.950 1952.770 2603.330 1952.780 ;
        RECT 2599.460 1952.720 2603.330 1952.770 ;
        RECT 2596.000 1952.470 2603.330 1952.720 ;
        RECT 2596.000 1952.120 2600.000 1952.470 ;
        RECT 2602.950 1952.460 2603.330 1952.470 ;
      LAYER via3 ;
        RECT 2602.980 3502.180 2603.300 3502.500 ;
        RECT 2602.980 1952.460 2603.300 1952.780 ;
      LAYER met4 ;
        RECT 2602.975 3502.175 2603.305 3502.505 ;
        RECT 2602.990 1952.785 2603.290 3502.175 ;
        RECT 2602.975 1952.455 2603.305 1952.785 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 2603.870 3339.970 2604.250 3339.980 ;
        RECT -4.800 3339.670 2604.250 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 2603.870 3339.660 2604.250 3339.670 ;
        RECT 2603.870 1984.050 2604.250 1984.060 ;
        RECT 2599.460 1984.000 2604.250 1984.050 ;
        RECT 2596.000 1983.750 2604.250 1984.000 ;
        RECT 2596.000 1983.400 2600.000 1983.750 ;
        RECT 2603.870 1983.740 2604.250 1983.750 ;
      LAYER via3 ;
        RECT 2603.900 3339.660 2604.220 3339.980 ;
        RECT 2603.900 1983.740 2604.220 1984.060 ;
      LAYER met4 ;
        RECT 2603.895 3339.655 2604.225 3339.985 ;
        RECT 2603.910 1984.065 2604.210 3339.655 ;
        RECT 2603.895 1983.735 2604.225 1984.065 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3051.740 17.410 3051.800 ;
        RECT 2604.130 3051.740 2604.450 3051.800 ;
        RECT 17.090 3051.600 2604.450 3051.740 ;
        RECT 17.090 3051.540 17.410 3051.600 ;
        RECT 2604.130 3051.540 2604.450 3051.600 ;
        RECT 2604.130 2184.060 2604.450 2184.120 ;
        RECT 2606.430 2184.060 2606.750 2184.120 ;
        RECT 2604.130 2183.920 2606.750 2184.060 ;
        RECT 2604.130 2183.860 2604.450 2183.920 ;
        RECT 2606.430 2183.860 2606.750 2183.920 ;
      LAYER via ;
        RECT 17.120 3051.540 17.380 3051.800 ;
        RECT 2604.160 3051.540 2604.420 3051.800 ;
        RECT 2604.160 2183.860 2604.420 2184.120 ;
        RECT 2606.460 2183.860 2606.720 2184.120 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3051.830 17.320 3051.995 ;
        RECT 17.120 3051.510 17.380 3051.830 ;
        RECT 2604.160 3051.510 2604.420 3051.830 ;
        RECT 2604.220 2404.890 2604.360 3051.510 ;
        RECT 2604.220 2404.750 2606.660 2404.890 ;
        RECT 2606.520 2184.150 2606.660 2404.750 ;
        RECT 2604.160 2183.830 2604.420 2184.150 ;
        RECT 2606.460 2183.830 2606.720 2184.150 ;
        RECT 2604.220 2016.045 2604.360 2183.830 ;
        RECT 2604.150 2015.675 2604.430 2016.045 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 2604.150 2015.720 2604.430 2016.000 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 2604.125 2016.010 2604.455 2016.025 ;
        RECT 2599.460 2015.960 2604.455 2016.010 ;
        RECT 2596.000 2015.710 2604.455 2015.960 ;
        RECT 2596.000 2015.360 2600.000 2015.710 ;
        RECT 2604.125 2015.695 2604.455 2015.710 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 2397.580 18.790 2397.640 ;
        RECT 2613.790 2397.580 2614.110 2397.640 ;
        RECT 18.470 2397.440 2614.110 2397.580 ;
        RECT 18.470 2397.380 18.790 2397.440 ;
        RECT 2613.790 2397.380 2614.110 2397.440 ;
      LAYER via ;
        RECT 18.500 2397.380 18.760 2397.640 ;
        RECT 2613.820 2397.380 2614.080 2397.640 ;
      LAYER met2 ;
        RECT 18.490 2765.035 18.770 2765.405 ;
        RECT 18.560 2397.670 18.700 2765.035 ;
        RECT 18.500 2397.350 18.760 2397.670 ;
        RECT 2613.820 2397.350 2614.080 2397.670 ;
        RECT 2613.880 2047.325 2614.020 2397.350 ;
        RECT 2613.810 2046.955 2614.090 2047.325 ;
      LAYER via2 ;
        RECT 18.490 2765.080 18.770 2765.360 ;
        RECT 2613.810 2047.000 2614.090 2047.280 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 18.465 2765.370 18.795 2765.385 ;
        RECT -4.800 2765.070 18.795 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 18.465 2765.055 18.795 2765.070 ;
        RECT 2613.785 2047.290 2614.115 2047.305 ;
        RECT 2599.460 2047.240 2614.115 2047.290 ;
        RECT 2596.000 2046.990 2614.115 2047.240 ;
        RECT 2596.000 2046.640 2600.000 2046.990 ;
        RECT 2613.785 2046.975 2614.115 2046.990 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2477.480 17.410 2477.540 ;
        RECT 2606.430 2477.480 2606.750 2477.540 ;
        RECT 17.090 2477.340 2606.750 2477.480 ;
        RECT 17.090 2477.280 17.410 2477.340 ;
        RECT 2606.430 2477.280 2606.750 2477.340 ;
        RECT 2607.350 2380.580 2607.670 2380.640 ;
        RECT 2608.730 2380.580 2609.050 2380.640 ;
        RECT 2607.350 2380.440 2609.050 2380.580 ;
        RECT 2607.350 2380.380 2607.670 2380.440 ;
        RECT 2608.730 2380.380 2609.050 2380.440 ;
        RECT 2607.350 2209.360 2607.670 2209.620 ;
        RECT 2607.440 2208.260 2607.580 2209.360 ;
        RECT 2607.350 2208.000 2607.670 2208.260 ;
        RECT 2606.430 2111.640 2606.750 2111.700 ;
        RECT 2607.350 2111.640 2607.670 2111.700 ;
        RECT 2606.430 2111.500 2607.670 2111.640 ;
        RECT 2606.430 2111.440 2606.750 2111.500 ;
        RECT 2607.350 2111.440 2607.670 2111.500 ;
      LAYER via ;
        RECT 17.120 2477.280 17.380 2477.540 ;
        RECT 2606.460 2477.280 2606.720 2477.540 ;
        RECT 2607.380 2380.380 2607.640 2380.640 ;
        RECT 2608.760 2380.380 2609.020 2380.640 ;
        RECT 2607.380 2209.360 2607.640 2209.620 ;
        RECT 2607.380 2208.000 2607.640 2208.260 ;
        RECT 2606.460 2111.440 2606.720 2111.700 ;
        RECT 2607.380 2111.440 2607.640 2111.700 ;
      LAYER met2 ;
        RECT 17.110 2477.395 17.390 2477.765 ;
        RECT 17.120 2477.250 17.380 2477.395 ;
        RECT 2606.460 2477.250 2606.720 2477.570 ;
        RECT 2606.520 2405.570 2606.660 2477.250 ;
        RECT 2606.520 2405.430 2608.040 2405.570 ;
        RECT 2607.900 2398.090 2608.040 2405.430 ;
        RECT 2607.900 2397.950 2608.960 2398.090 ;
        RECT 2608.820 2380.670 2608.960 2397.950 ;
        RECT 2607.380 2380.350 2607.640 2380.670 ;
        RECT 2608.760 2380.350 2609.020 2380.670 ;
        RECT 2607.440 2256.085 2607.580 2380.350 ;
        RECT 2607.370 2255.715 2607.650 2256.085 ;
        RECT 2607.370 2209.475 2607.650 2209.845 ;
        RECT 2607.380 2209.330 2607.640 2209.475 ;
        RECT 2607.380 2207.970 2607.640 2208.290 ;
        RECT 2607.440 2111.730 2607.580 2207.970 ;
        RECT 2606.460 2111.410 2606.720 2111.730 ;
        RECT 2607.380 2111.410 2607.640 2111.730 ;
        RECT 2606.520 2079.285 2606.660 2111.410 ;
        RECT 2606.450 2078.915 2606.730 2079.285 ;
      LAYER via2 ;
        RECT 17.110 2477.440 17.390 2477.720 ;
        RECT 2607.370 2255.760 2607.650 2256.040 ;
        RECT 2607.370 2209.520 2607.650 2209.800 ;
        RECT 2606.450 2078.960 2606.730 2079.240 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 17.085 2477.730 17.415 2477.745 ;
        RECT -4.800 2477.430 17.415 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 17.085 2477.415 17.415 2477.430 ;
        RECT 2607.345 2256.060 2607.675 2256.065 ;
        RECT 2607.345 2256.050 2607.930 2256.060 ;
        RECT 2607.345 2255.750 2608.130 2256.050 ;
        RECT 2607.345 2255.740 2607.930 2255.750 ;
        RECT 2607.345 2255.735 2607.675 2255.740 ;
        RECT 2607.345 2209.820 2607.675 2209.825 ;
        RECT 2607.345 2209.810 2607.930 2209.820 ;
        RECT 2607.120 2209.510 2607.930 2209.810 ;
        RECT 2607.345 2209.500 2607.930 2209.510 ;
        RECT 2607.345 2209.495 2607.675 2209.500 ;
        RECT 2606.425 2079.250 2606.755 2079.265 ;
        RECT 2599.460 2079.200 2606.755 2079.250 ;
        RECT 2596.000 2078.950 2606.755 2079.200 ;
        RECT 2596.000 2078.600 2600.000 2078.950 ;
        RECT 2606.425 2078.935 2606.755 2078.950 ;
      LAYER via3 ;
        RECT 2607.580 2255.740 2607.900 2256.060 ;
        RECT 2607.580 2209.500 2607.900 2209.820 ;
      LAYER met4 ;
        RECT 2607.575 2255.735 2607.905 2256.065 ;
        RECT 2607.590 2209.825 2607.890 2255.735 ;
        RECT 2607.575 2209.495 2607.905 2209.825 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1396.170 2392.480 1396.490 2392.540 ;
        RECT 2615.630 2392.480 2615.950 2392.540 ;
        RECT 1396.170 2392.340 2615.950 2392.480 ;
        RECT 1396.170 2392.280 1396.490 2392.340 ;
        RECT 2615.630 2392.280 2615.950 2392.340 ;
        RECT 17.550 2194.260 17.870 2194.320 ;
        RECT 1396.170 2194.260 1396.490 2194.320 ;
        RECT 17.550 2194.120 1396.490 2194.260 ;
        RECT 17.550 2194.060 17.870 2194.120 ;
        RECT 1396.170 2194.060 1396.490 2194.120 ;
      LAYER via ;
        RECT 1396.200 2392.280 1396.460 2392.540 ;
        RECT 2615.660 2392.280 2615.920 2392.540 ;
        RECT 17.580 2194.060 17.840 2194.320 ;
        RECT 1396.200 2194.060 1396.460 2194.320 ;
      LAYER met2 ;
        RECT 1396.200 2392.250 1396.460 2392.570 ;
        RECT 2615.660 2392.250 2615.920 2392.570 ;
        RECT 1396.260 2194.350 1396.400 2392.250 ;
        RECT 17.580 2194.030 17.840 2194.350 ;
        RECT 1396.200 2194.030 1396.460 2194.350 ;
        RECT 17.640 2190.125 17.780 2194.030 ;
        RECT 17.570 2189.755 17.850 2190.125 ;
        RECT 2615.720 2110.565 2615.860 2392.250 ;
        RECT 2615.650 2110.195 2615.930 2110.565 ;
      LAYER via2 ;
        RECT 17.570 2189.800 17.850 2190.080 ;
        RECT 2615.650 2110.240 2615.930 2110.520 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 17.545 2190.090 17.875 2190.105 ;
        RECT -4.800 2189.790 17.875 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 17.545 2189.775 17.875 2189.790 ;
        RECT 2615.625 2110.530 2615.955 2110.545 ;
        RECT 2599.460 2110.480 2615.955 2110.530 ;
        RECT 2596.000 2110.230 2615.955 2110.480 ;
        RECT 2596.000 2109.880 2600.000 2110.230 ;
        RECT 2615.625 2110.215 2615.955 2110.230 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1399.850 2395.540 1400.170 2395.600 ;
        RECT 2616.550 2395.540 2616.870 2395.600 ;
        RECT 1399.850 2395.400 2616.870 2395.540 ;
        RECT 1399.850 2395.340 1400.170 2395.400 ;
        RECT 2616.550 2395.340 2616.870 2395.400 ;
        RECT 2608.270 2141.900 2608.590 2141.960 ;
        RECT 2616.550 2141.900 2616.870 2141.960 ;
        RECT 2608.270 2141.760 2616.870 2141.900 ;
        RECT 2608.270 2141.700 2608.590 2141.760 ;
        RECT 2616.550 2141.700 2616.870 2141.760 ;
        RECT 17.550 1904.240 17.870 1904.300 ;
        RECT 1399.850 1904.240 1400.170 1904.300 ;
        RECT 17.550 1904.100 1400.170 1904.240 ;
        RECT 17.550 1904.040 17.870 1904.100 ;
        RECT 1399.850 1904.040 1400.170 1904.100 ;
      LAYER via ;
        RECT 1399.880 2395.340 1400.140 2395.600 ;
        RECT 2616.580 2395.340 2616.840 2395.600 ;
        RECT 2608.300 2141.700 2608.560 2141.960 ;
        RECT 2616.580 2141.700 2616.840 2141.960 ;
        RECT 17.580 1904.040 17.840 1904.300 ;
        RECT 1399.880 1904.040 1400.140 1904.300 ;
      LAYER met2 ;
        RECT 1399.880 2395.310 1400.140 2395.630 ;
        RECT 2616.580 2395.310 2616.840 2395.630 ;
        RECT 1399.940 1904.330 1400.080 2395.310 ;
        RECT 2616.640 2141.990 2616.780 2395.310 ;
        RECT 2608.300 2141.845 2608.560 2141.990 ;
        RECT 2608.290 2141.475 2608.570 2141.845 ;
        RECT 2616.580 2141.670 2616.840 2141.990 ;
        RECT 17.580 1904.010 17.840 1904.330 ;
        RECT 1399.880 1904.010 1400.140 1904.330 ;
        RECT 17.640 1903.165 17.780 1904.010 ;
        RECT 17.570 1902.795 17.850 1903.165 ;
      LAYER via2 ;
        RECT 2608.290 2141.520 2608.570 2141.800 ;
        RECT 17.570 1902.840 17.850 1903.120 ;
      LAYER met3 ;
        RECT 2608.265 2141.810 2608.595 2141.825 ;
        RECT 2599.460 2141.760 2608.595 2141.810 ;
        RECT 2596.000 2141.510 2608.595 2141.760 ;
        RECT 2596.000 2141.160 2600.000 2141.510 ;
        RECT 2608.265 2141.495 2608.595 2141.510 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 17.545 1903.130 17.875 1903.145 ;
        RECT -4.800 1902.830 17.875 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 17.545 1902.815 17.875 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2613.330 620.740 2613.650 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2613.330 620.600 2901.150 620.740 ;
        RECT 2613.330 620.540 2613.650 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2613.360 620.540 2613.620 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2613.350 1288.755 2613.630 1289.125 ;
        RECT 2613.420 620.830 2613.560 1288.755 ;
        RECT 2613.360 620.510 2613.620 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2613.350 1288.800 2613.630 1289.080 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 2613.325 1289.090 2613.655 1289.105 ;
        RECT 2599.460 1289.040 2613.655 1289.090 ;
        RECT 2596.000 1288.790 2613.655 1289.040 ;
        RECT 2596.000 1288.440 2600.000 1288.790 ;
        RECT 2613.325 1288.775 2613.655 1288.790 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2607.350 2397.240 2607.670 2397.300 ;
        RECT 2597.320 2397.100 2607.670 2397.240 ;
        RECT 1398.470 2396.900 1398.790 2396.960 ;
        RECT 2597.320 2396.900 2597.460 2397.100 ;
        RECT 2607.350 2397.040 2607.670 2397.100 ;
        RECT 1398.470 2396.760 2597.460 2396.900 ;
        RECT 1398.470 2396.700 1398.790 2396.760 ;
        RECT 2607.810 2332.300 2608.130 2332.360 ;
        RECT 2608.730 2332.300 2609.050 2332.360 ;
        RECT 2607.810 2332.160 2609.050 2332.300 ;
        RECT 2607.810 2332.100 2608.130 2332.160 ;
        RECT 2608.730 2332.100 2609.050 2332.160 ;
        RECT 17.550 1621.360 17.870 1621.420 ;
        RECT 1398.470 1621.360 1398.790 1621.420 ;
        RECT 17.550 1621.220 1398.790 1621.360 ;
        RECT 17.550 1621.160 17.870 1621.220 ;
        RECT 1398.470 1621.160 1398.790 1621.220 ;
      LAYER via ;
        RECT 1398.500 2396.700 1398.760 2396.960 ;
        RECT 2607.380 2397.040 2607.640 2397.300 ;
        RECT 2607.840 2332.100 2608.100 2332.360 ;
        RECT 2608.760 2332.100 2609.020 2332.360 ;
        RECT 17.580 1621.160 17.840 1621.420 ;
        RECT 1398.500 1621.160 1398.760 1621.420 ;
      LAYER met2 ;
        RECT 2607.380 2397.010 2607.640 2397.330 ;
        RECT 1398.500 2396.670 1398.760 2396.990 ;
        RECT 1398.560 1621.450 1398.700 2396.670 ;
        RECT 2607.440 2381.090 2607.580 2397.010 ;
        RECT 2607.440 2380.950 2608.040 2381.090 ;
        RECT 2607.900 2332.390 2608.040 2380.950 ;
        RECT 2607.840 2332.070 2608.100 2332.390 ;
        RECT 2608.760 2332.070 2609.020 2332.390 ;
        RECT 2608.820 2331.450 2608.960 2332.070 ;
        RECT 2607.900 2331.310 2608.960 2331.450 ;
        RECT 2607.900 2209.165 2608.040 2331.310 ;
        RECT 2607.830 2208.795 2608.110 2209.165 ;
        RECT 17.580 1621.130 17.840 1621.450 ;
        RECT 1398.500 1621.130 1398.760 1621.450 ;
        RECT 17.640 1615.525 17.780 1621.130 ;
        RECT 17.570 1615.155 17.850 1615.525 ;
      LAYER via2 ;
        RECT 2607.830 2208.840 2608.110 2209.120 ;
        RECT 17.570 1615.200 17.850 1615.480 ;
      LAYER met3 ;
        RECT 2607.805 2209.140 2608.135 2209.145 ;
        RECT 2607.550 2209.130 2608.135 2209.140 ;
        RECT 2607.350 2208.830 2608.135 2209.130 ;
        RECT 2607.550 2208.820 2608.135 2208.830 ;
        RECT 2607.805 2208.815 2608.135 2208.820 ;
        RECT 2607.550 2176.490 2607.930 2176.500 ;
        RECT 2599.310 2176.190 2607.930 2176.490 ;
        RECT 2599.310 2173.720 2599.610 2176.190 ;
        RECT 2607.550 2176.180 2607.930 2176.190 ;
        RECT 2596.000 2173.120 2600.000 2173.720 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 17.545 1615.490 17.875 1615.505 ;
        RECT -4.800 1615.190 17.875 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 17.545 1615.175 17.875 1615.190 ;
      LAYER via3 ;
        RECT 2607.580 2208.820 2607.900 2209.140 ;
        RECT 2607.580 2176.180 2607.900 2176.500 ;
      LAYER met4 ;
        RECT 2607.575 2208.815 2607.905 2209.145 ;
        RECT 2607.590 2176.505 2607.890 2208.815 ;
        RECT 2607.575 2176.175 2607.905 2176.505 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1397.090 2395.880 1397.410 2395.940 ;
        RECT 2611.950 2395.880 2612.270 2395.940 ;
        RECT 1397.090 2395.740 2612.270 2395.880 ;
        RECT 1397.090 2395.680 1397.410 2395.740 ;
        RECT 2611.950 2395.680 2612.270 2395.740 ;
        RECT 17.550 1400.700 17.870 1400.760 ;
        RECT 1397.090 1400.700 1397.410 1400.760 ;
        RECT 17.550 1400.560 1397.410 1400.700 ;
        RECT 17.550 1400.500 17.870 1400.560 ;
        RECT 1397.090 1400.500 1397.410 1400.560 ;
      LAYER via ;
        RECT 1397.120 2395.680 1397.380 2395.940 ;
        RECT 2611.980 2395.680 2612.240 2395.940 ;
        RECT 17.580 1400.500 17.840 1400.760 ;
        RECT 1397.120 1400.500 1397.380 1400.760 ;
      LAYER met2 ;
        RECT 1397.120 2395.650 1397.380 2395.970 ;
        RECT 2611.980 2395.650 2612.240 2395.970 ;
        RECT 1397.180 1400.790 1397.320 2395.650 ;
        RECT 2612.040 2205.085 2612.180 2395.650 ;
        RECT 2611.970 2204.715 2612.250 2205.085 ;
        RECT 17.580 1400.645 17.840 1400.790 ;
        RECT 17.570 1400.275 17.850 1400.645 ;
        RECT 1397.120 1400.470 1397.380 1400.790 ;
      LAYER via2 ;
        RECT 2611.970 2204.760 2612.250 2205.040 ;
        RECT 17.570 1400.320 17.850 1400.600 ;
      LAYER met3 ;
        RECT 2611.945 2205.050 2612.275 2205.065 ;
        RECT 2599.460 2205.000 2612.275 2205.050 ;
        RECT 2596.000 2204.750 2612.275 2205.000 ;
        RECT 2596.000 2204.400 2600.000 2204.750 ;
        RECT 2611.945 2204.735 2612.275 2204.750 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.545 1400.610 17.875 1400.625 ;
        RECT -4.800 1400.310 17.875 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.545 1400.295 17.875 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 1186.840 17.870 1186.900 ;
        RECT 2612.410 1186.840 2612.730 1186.900 ;
        RECT 17.550 1186.700 2612.730 1186.840 ;
        RECT 17.550 1186.640 17.870 1186.700 ;
        RECT 2612.410 1186.640 2612.730 1186.700 ;
      LAYER via ;
        RECT 17.580 1186.640 17.840 1186.900 ;
        RECT 2612.440 1186.640 2612.700 1186.900 ;
      LAYER met2 ;
        RECT 2612.430 2236.675 2612.710 2237.045 ;
        RECT 2612.500 1186.930 2612.640 2236.675 ;
        RECT 17.580 1186.610 17.840 1186.930 ;
        RECT 2612.440 1186.610 2612.700 1186.930 ;
        RECT 17.640 1185.085 17.780 1186.610 ;
        RECT 17.570 1184.715 17.850 1185.085 ;
      LAYER via2 ;
        RECT 2612.430 2236.720 2612.710 2237.000 ;
        RECT 17.570 1184.760 17.850 1185.040 ;
      LAYER met3 ;
        RECT 2612.405 2237.010 2612.735 2237.025 ;
        RECT 2599.460 2236.960 2612.735 2237.010 ;
        RECT 2596.000 2236.710 2612.735 2236.960 ;
        RECT 2596.000 2236.360 2600.000 2236.710 ;
        RECT 2612.405 2236.695 2612.735 2236.710 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.545 1185.050 17.875 1185.065 ;
        RECT -4.800 1184.750 17.875 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.545 1184.735 17.875 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 1005.280 15.110 1005.340 ;
        RECT 2610.110 1005.280 2610.430 1005.340 ;
        RECT 14.790 1005.140 2610.430 1005.280 ;
        RECT 14.790 1005.080 15.110 1005.140 ;
        RECT 2610.110 1005.080 2610.430 1005.140 ;
      LAYER via ;
        RECT 14.820 1005.080 15.080 1005.340 ;
        RECT 2610.140 1005.080 2610.400 1005.340 ;
      LAYER met2 ;
        RECT 2610.130 2267.955 2610.410 2268.325 ;
        RECT 2610.200 1005.370 2610.340 2267.955 ;
        RECT 14.820 1005.050 15.080 1005.370 ;
        RECT 2610.140 1005.050 2610.400 1005.370 ;
        RECT 14.880 969.525 15.020 1005.050 ;
        RECT 14.810 969.155 15.090 969.525 ;
      LAYER via2 ;
        RECT 2610.130 2268.000 2610.410 2268.280 ;
        RECT 14.810 969.200 15.090 969.480 ;
      LAYER met3 ;
        RECT 2610.105 2268.290 2610.435 2268.305 ;
        RECT 2599.460 2268.240 2610.435 2268.290 ;
        RECT 2596.000 2267.990 2610.435 2268.240 ;
        RECT 2596.000 2267.640 2600.000 2267.990 ;
        RECT 2610.105 2267.975 2610.435 2267.990 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 14.785 969.490 15.115 969.505 ;
        RECT -4.800 969.190 15.115 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 14.785 969.175 15.115 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 1005.620 18.790 1005.680 ;
        RECT 2608.730 1005.620 2609.050 1005.680 ;
        RECT 18.470 1005.480 2609.050 1005.620 ;
        RECT 18.470 1005.420 18.790 1005.480 ;
        RECT 2608.730 1005.420 2609.050 1005.480 ;
      LAYER via ;
        RECT 18.500 1005.420 18.760 1005.680 ;
        RECT 2608.760 1005.420 2609.020 1005.680 ;
      LAYER met2 ;
        RECT 2608.750 2299.915 2609.030 2300.285 ;
        RECT 2608.820 1005.710 2608.960 2299.915 ;
        RECT 18.500 1005.390 18.760 1005.710 ;
        RECT 2608.760 1005.390 2609.020 1005.710 ;
        RECT 18.560 753.965 18.700 1005.390 ;
        RECT 18.490 753.595 18.770 753.965 ;
      LAYER via2 ;
        RECT 2608.750 2299.960 2609.030 2300.240 ;
        RECT 18.490 753.640 18.770 753.920 ;
      LAYER met3 ;
        RECT 2608.725 2300.250 2609.055 2300.265 ;
        RECT 2599.460 2300.200 2609.055 2300.250 ;
        RECT 2596.000 2299.950 2609.055 2300.200 ;
        RECT 2596.000 2299.600 2600.000 2299.950 ;
        RECT 2608.725 2299.935 2609.055 2299.950 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 18.465 753.930 18.795 753.945 ;
        RECT -4.800 753.630 18.795 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 18.465 753.615 18.795 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 544.155 17.850 544.525 ;
        RECT 17.640 538.405 17.780 544.155 ;
        RECT 17.570 538.035 17.850 538.405 ;
      LAYER via2 ;
        RECT 17.570 544.200 17.850 544.480 ;
        RECT 17.570 538.080 17.850 538.360 ;
      LAYER met3 ;
        RECT 2613.070 2331.530 2613.450 2331.540 ;
        RECT 2599.460 2331.480 2613.450 2331.530 ;
        RECT 2596.000 2331.230 2613.450 2331.480 ;
        RECT 2596.000 2330.880 2600.000 2331.230 ;
        RECT 2613.070 2331.220 2613.450 2331.230 ;
        RECT 17.545 544.490 17.875 544.505 ;
        RECT 2613.070 544.490 2613.450 544.500 ;
        RECT 17.545 544.190 2613.450 544.490 ;
        RECT 17.545 544.175 17.875 544.190 ;
        RECT 2613.070 544.180 2613.450 544.190 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 17.545 538.370 17.875 538.385 ;
        RECT -4.800 538.070 17.875 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 17.545 538.055 17.875 538.070 ;
      LAYER via3 ;
        RECT 2613.100 2331.220 2613.420 2331.540 ;
        RECT 2613.100 544.180 2613.420 544.500 ;
      LAYER met4 ;
        RECT 2613.095 2331.215 2613.425 2331.545 ;
        RECT 2613.110 544.505 2613.410 2331.215 ;
        RECT 2613.095 544.175 2613.425 544.505 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2601.110 2363.490 2601.490 2363.500 ;
        RECT 2599.460 2363.440 2601.490 2363.490 ;
        RECT 2596.000 2363.190 2601.490 2363.440 ;
        RECT 2596.000 2362.840 2600.000 2363.190 ;
        RECT 2601.110 2363.180 2601.490 2363.190 ;
        RECT 2601.110 324.170 2601.490 324.180 ;
        RECT 3.070 323.870 2601.490 324.170 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 3.070 322.810 3.370 323.870 ;
        RECT 2601.110 323.860 2601.490 323.870 ;
        RECT -4.800 322.510 3.370 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
      LAYER via3 ;
        RECT 2601.140 2363.180 2601.460 2363.500 ;
        RECT 2601.140 323.860 2601.460 324.180 ;
      LAYER met4 ;
        RECT 2601.135 2363.175 2601.465 2363.505 ;
        RECT 2601.150 324.185 2601.450 2363.175 ;
        RECT 2601.135 323.855 2601.465 324.185 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2394.520 17.410 2394.580 ;
        RECT 2608.270 2394.520 2608.590 2394.580 ;
        RECT 17.090 2394.380 2608.590 2394.520 ;
        RECT 17.090 2394.320 17.410 2394.380 ;
        RECT 2608.270 2394.320 2608.590 2394.380 ;
      LAYER via ;
        RECT 17.120 2394.320 17.380 2394.580 ;
        RECT 2608.300 2394.320 2608.560 2394.580 ;
      LAYER met2 ;
        RECT 17.120 2394.290 17.380 2394.610 ;
        RECT 2608.290 2394.435 2608.570 2394.805 ;
        RECT 2608.300 2394.290 2608.560 2394.435 ;
        RECT 17.180 107.285 17.320 2394.290 ;
        RECT 17.110 106.915 17.390 107.285 ;
      LAYER via2 ;
        RECT 2608.290 2394.480 2608.570 2394.760 ;
        RECT 17.110 106.960 17.390 107.240 ;
      LAYER met3 ;
        RECT 2608.265 2394.770 2608.595 2394.785 ;
        RECT 2599.460 2394.720 2608.595 2394.770 ;
        RECT 2596.000 2394.470 2608.595 2394.720 ;
        RECT 2596.000 2394.120 2600.000 2394.470 ;
        RECT 2608.265 2394.455 2608.595 2394.470 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 17.085 107.250 17.415 107.265 ;
        RECT -4.800 106.950 17.415 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 17.085 106.935 17.415 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2613.790 1318.080 2614.110 1318.140 ;
        RECT 2619.310 1318.080 2619.630 1318.140 ;
        RECT 2613.790 1317.940 2619.630 1318.080 ;
        RECT 2613.790 1317.880 2614.110 1317.940 ;
        RECT 2619.310 1317.880 2619.630 1317.940 ;
        RECT 2619.310 855.340 2619.630 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2619.310 855.200 2901.150 855.340 ;
        RECT 2619.310 855.140 2619.630 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2613.820 1317.880 2614.080 1318.140 ;
        RECT 2619.340 1317.880 2619.600 1318.140 ;
        RECT 2619.340 855.140 2619.600 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2613.810 1320.715 2614.090 1321.085 ;
        RECT 2613.880 1318.170 2614.020 1320.715 ;
        RECT 2613.820 1317.850 2614.080 1318.170 ;
        RECT 2619.340 1317.850 2619.600 1318.170 ;
        RECT 2619.400 855.430 2619.540 1317.850 ;
        RECT 2619.340 855.110 2619.600 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2613.810 1320.760 2614.090 1321.040 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2613.785 1321.050 2614.115 1321.065 ;
        RECT 2599.460 1321.000 2614.115 1321.050 ;
        RECT 2596.000 1320.750 2614.115 1321.000 ;
        RECT 2596.000 1320.400 2600.000 1320.750 ;
        RECT 2613.785 1320.735 2614.115 1320.750 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2614.250 1345.620 2614.570 1345.680 ;
        RECT 2620.690 1345.620 2621.010 1345.680 ;
        RECT 2614.250 1345.480 2621.010 1345.620 ;
        RECT 2614.250 1345.420 2614.570 1345.480 ;
        RECT 2620.690 1345.420 2621.010 1345.480 ;
        RECT 2620.690 1089.940 2621.010 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2620.690 1089.800 2901.150 1089.940 ;
        RECT 2620.690 1089.740 2621.010 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2614.280 1345.420 2614.540 1345.680 ;
        RECT 2620.720 1345.420 2620.980 1345.680 ;
        RECT 2620.720 1089.740 2620.980 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2614.270 1351.995 2614.550 1352.365 ;
        RECT 2614.340 1345.710 2614.480 1351.995 ;
        RECT 2614.280 1345.390 2614.540 1345.710 ;
        RECT 2620.720 1345.390 2620.980 1345.710 ;
        RECT 2620.780 1090.030 2620.920 1345.390 ;
        RECT 2620.720 1089.710 2620.980 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2614.270 1352.040 2614.550 1352.320 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2614.245 1352.330 2614.575 1352.345 ;
        RECT 2599.460 1352.280 2614.575 1352.330 ;
        RECT 2596.000 1352.030 2614.575 1352.280 ;
        RECT 2596.000 1351.680 2600.000 1352.030 ;
        RECT 2614.245 1352.015 2614.575 1352.030 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2612.870 1328.280 2613.190 1328.340 ;
        RECT 2900.830 1328.280 2901.150 1328.340 ;
        RECT 2612.870 1328.140 2901.150 1328.280 ;
        RECT 2612.870 1328.080 2613.190 1328.140 ;
        RECT 2900.830 1328.080 2901.150 1328.140 ;
      LAYER via ;
        RECT 2612.900 1328.080 2613.160 1328.340 ;
        RECT 2900.860 1328.080 2901.120 1328.340 ;
      LAYER met2 ;
        RECT 2612.890 1383.955 2613.170 1384.325 ;
        RECT 2612.960 1328.370 2613.100 1383.955 ;
        RECT 2612.900 1328.050 2613.160 1328.370 ;
        RECT 2900.860 1328.050 2901.120 1328.370 ;
        RECT 2900.920 1319.725 2901.060 1328.050 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2612.890 1384.000 2613.170 1384.280 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2612.865 1384.290 2613.195 1384.305 ;
        RECT 2599.460 1384.240 2613.195 1384.290 ;
        RECT 2596.000 1383.990 2613.195 1384.240 ;
        RECT 2596.000 1383.640 2600.000 1383.990 ;
        RECT 2612.865 1383.975 2613.195 1383.990 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2613.330 1473.460 2613.650 1473.520 ;
        RECT 2903.590 1473.460 2903.910 1473.520 ;
        RECT 2613.330 1473.320 2903.910 1473.460 ;
        RECT 2613.330 1473.260 2613.650 1473.320 ;
        RECT 2903.590 1473.260 2903.910 1473.320 ;
      LAYER via ;
        RECT 2613.360 1473.260 2613.620 1473.520 ;
        RECT 2903.620 1473.260 2903.880 1473.520 ;
      LAYER met2 ;
        RECT 2903.610 1553.955 2903.890 1554.325 ;
        RECT 2903.680 1473.550 2903.820 1553.955 ;
        RECT 2613.360 1473.230 2613.620 1473.550 ;
        RECT 2903.620 1473.230 2903.880 1473.550 ;
        RECT 2613.420 1415.605 2613.560 1473.230 ;
        RECT 2613.350 1415.235 2613.630 1415.605 ;
      LAYER via2 ;
        RECT 2903.610 1554.000 2903.890 1554.280 ;
        RECT 2613.350 1415.280 2613.630 1415.560 ;
      LAYER met3 ;
        RECT 2903.585 1554.290 2903.915 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2903.585 1553.990 2924.800 1554.290 ;
        RECT 2903.585 1553.975 2903.915 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 2613.325 1415.570 2613.655 1415.585 ;
        RECT 2599.460 1415.520 2613.655 1415.570 ;
        RECT 2596.000 1415.270 2613.655 1415.520 ;
        RECT 2596.000 1414.920 2600.000 1415.270 ;
        RECT 2613.325 1415.255 2613.655 1415.270 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2614.250 1448.980 2614.570 1449.040 ;
        RECT 2902.210 1448.980 2902.530 1449.040 ;
        RECT 2614.250 1448.840 2902.530 1448.980 ;
        RECT 2614.250 1448.780 2614.570 1448.840 ;
        RECT 2902.210 1448.780 2902.530 1448.840 ;
      LAYER via ;
        RECT 2614.280 1448.780 2614.540 1449.040 ;
        RECT 2902.240 1448.780 2902.500 1449.040 ;
      LAYER met2 ;
        RECT 2902.230 1789.235 2902.510 1789.605 ;
        RECT 2902.300 1449.070 2902.440 1789.235 ;
        RECT 2614.280 1448.750 2614.540 1449.070 ;
        RECT 2902.240 1448.750 2902.500 1449.070 ;
        RECT 2614.340 1447.565 2614.480 1448.750 ;
        RECT 2614.270 1447.195 2614.550 1447.565 ;
      LAYER via2 ;
        RECT 2902.230 1789.280 2902.510 1789.560 ;
        RECT 2614.270 1447.240 2614.550 1447.520 ;
      LAYER met3 ;
        RECT 2902.205 1789.570 2902.535 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2902.205 1789.270 2924.800 1789.570 ;
        RECT 2902.205 1789.255 2902.535 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2614.245 1447.530 2614.575 1447.545 ;
        RECT 2599.460 1447.480 2614.575 1447.530 ;
        RECT 2596.000 1447.230 2614.575 1447.480 ;
        RECT 2596.000 1446.880 2600.000 1447.230 ;
        RECT 2614.245 1447.215 2614.575 1447.230 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2613.790 1483.320 2614.110 1483.380 ;
        RECT 2901.290 1483.320 2901.610 1483.380 ;
        RECT 2613.790 1483.180 2901.610 1483.320 ;
        RECT 2613.790 1483.120 2614.110 1483.180 ;
        RECT 2901.290 1483.120 2901.610 1483.180 ;
      LAYER via ;
        RECT 2613.820 1483.120 2614.080 1483.380 ;
        RECT 2901.320 1483.120 2901.580 1483.380 ;
      LAYER met2 ;
        RECT 2901.310 2023.835 2901.590 2024.205 ;
        RECT 2901.380 1483.410 2901.520 2023.835 ;
        RECT 2613.820 1483.090 2614.080 1483.410 ;
        RECT 2901.320 1483.090 2901.580 1483.410 ;
        RECT 2613.880 1478.845 2614.020 1483.090 ;
        RECT 2613.810 1478.475 2614.090 1478.845 ;
      LAYER via2 ;
        RECT 2901.310 2023.880 2901.590 2024.160 ;
        RECT 2613.810 1478.520 2614.090 1478.800 ;
      LAYER met3 ;
        RECT 2901.285 2024.170 2901.615 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2901.285 2023.870 2924.800 2024.170 ;
        RECT 2901.285 2023.855 2901.615 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 2613.785 1478.810 2614.115 1478.825 ;
        RECT 2599.460 1478.760 2614.115 1478.810 ;
        RECT 2596.000 1478.510 2614.115 1478.760 ;
        RECT 2596.000 1478.160 2600.000 1478.510 ;
        RECT 2613.785 1478.495 2614.115 1478.510 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2818.490 2256.480 2818.810 2256.540 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 2818.490 2256.340 2901.150 2256.480 ;
        RECT 2818.490 2256.280 2818.810 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
        RECT 2614.250 1510.860 2614.570 1510.920 ;
        RECT 2818.490 1510.860 2818.810 1510.920 ;
        RECT 2614.250 1510.720 2818.810 1510.860 ;
        RECT 2614.250 1510.660 2614.570 1510.720 ;
        RECT 2818.490 1510.660 2818.810 1510.720 ;
      LAYER via ;
        RECT 2818.520 2256.280 2818.780 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
        RECT 2614.280 1510.660 2614.540 1510.920 ;
        RECT 2818.520 1510.660 2818.780 1510.920 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 2818.520 2256.250 2818.780 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 2818.580 1510.950 2818.720 2256.250 ;
        RECT 2614.280 1510.630 2614.540 1510.950 ;
        RECT 2818.520 1510.630 2818.780 1510.950 ;
        RECT 2614.340 1510.125 2614.480 1510.630 ;
        RECT 2614.270 1509.755 2614.550 1510.125 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
        RECT 2614.270 1509.800 2614.550 1510.080 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 2614.245 1510.090 2614.575 1510.105 ;
        RECT 2599.460 1510.040 2614.575 1510.090 ;
        RECT 2596.000 1509.790 2614.575 1510.040 ;
        RECT 2596.000 1509.440 2600.000 1509.790 ;
        RECT 2614.245 1509.775 2614.575 1509.790 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 634.410 2325.500 634.730 2325.560 ;
        RECT 1393.410 2325.500 1393.730 2325.560 ;
        RECT 634.410 2325.360 1393.730 2325.500 ;
        RECT 634.410 2325.300 634.730 2325.360 ;
        RECT 1393.410 2325.300 1393.730 2325.360 ;
      LAYER via ;
        RECT 634.440 2325.300 634.700 2325.560 ;
        RECT 1393.440 2325.300 1393.700 2325.560 ;
      LAYER met2 ;
        RECT 1393.430 2330.515 1393.710 2330.885 ;
        RECT 1393.500 2325.590 1393.640 2330.515 ;
        RECT 634.440 2325.270 634.700 2325.590 ;
        RECT 1393.440 2325.270 1393.700 2325.590 ;
        RECT 634.500 17.410 634.640 2325.270 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2330.560 1393.710 2330.840 ;
      LAYER met3 ;
        RECT 1393.405 2330.850 1393.735 2330.865 ;
        RECT 1393.405 2330.800 1400.700 2330.850 ;
        RECT 1393.405 2330.550 1404.000 2330.800 ;
        RECT 1393.405 2330.535 1393.735 2330.550 ;
        RECT 1400.000 2330.200 1404.000 2330.550 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 655.110 2360.180 655.430 2360.240 ;
        RECT 1393.410 2360.180 1393.730 2360.240 ;
        RECT 655.110 2360.040 1393.730 2360.180 ;
        RECT 655.110 2359.980 655.430 2360.040 ;
        RECT 1393.410 2359.980 1393.730 2360.040 ;
        RECT 650.970 17.920 651.290 17.980 ;
        RECT 655.110 17.920 655.430 17.980 ;
        RECT 650.970 17.780 655.430 17.920 ;
        RECT 650.970 17.720 651.290 17.780 ;
        RECT 655.110 17.720 655.430 17.780 ;
      LAYER via ;
        RECT 655.140 2359.980 655.400 2360.240 ;
        RECT 1393.440 2359.980 1393.700 2360.240 ;
        RECT 651.000 17.720 651.260 17.980 ;
        RECT 655.140 17.720 655.400 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2362.475 1393.710 2362.845 ;
        RECT 1393.500 2360.270 1393.640 2362.475 ;
        RECT 655.140 2359.950 655.400 2360.270 ;
        RECT 1393.440 2359.950 1393.700 2360.270 ;
        RECT 655.200 18.010 655.340 2359.950 ;
        RECT 651.000 17.690 651.260 18.010 ;
        RECT 655.140 17.690 655.400 18.010 ;
        RECT 651.060 2.400 651.200 17.690 ;
        RECT 650.850 -4.800 651.410 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2362.520 1393.710 2362.800 ;
      LAYER met3 ;
        RECT 1393.405 2362.810 1393.735 2362.825 ;
        RECT 1393.405 2362.760 1400.700 2362.810 ;
        RECT 1393.405 2362.510 1404.000 2362.760 ;
        RECT 1393.405 2362.495 1393.735 2362.510 ;
        RECT 1400.000 2362.160 1404.000 2362.510 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.310 2339.440 641.630 2339.500 ;
        RECT 1393.410 2339.440 1393.730 2339.500 ;
        RECT 641.310 2339.300 1393.730 2339.440 ;
        RECT 641.310 2339.240 641.630 2339.300 ;
        RECT 1393.410 2339.240 1393.730 2339.300 ;
        RECT 639.010 17.920 639.330 17.980 ;
        RECT 641.310 17.920 641.630 17.980 ;
        RECT 639.010 17.780 641.630 17.920 ;
        RECT 639.010 17.720 639.330 17.780 ;
        RECT 641.310 17.720 641.630 17.780 ;
      LAYER via ;
        RECT 641.340 2339.240 641.600 2339.500 ;
        RECT 1393.440 2339.240 1393.700 2339.500 ;
        RECT 639.040 17.720 639.300 17.980 ;
        RECT 641.340 17.720 641.600 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2341.395 1393.710 2341.765 ;
        RECT 1393.500 2339.530 1393.640 2341.395 ;
        RECT 641.340 2339.210 641.600 2339.530 ;
        RECT 1393.440 2339.210 1393.700 2339.530 ;
        RECT 641.400 18.010 641.540 2339.210 ;
        RECT 639.040 17.690 639.300 18.010 ;
        RECT 641.340 17.690 641.600 18.010 ;
        RECT 639.100 2.400 639.240 17.690 ;
        RECT 638.890 -4.800 639.450 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2341.440 1393.710 2341.720 ;
      LAYER met3 ;
        RECT 1393.405 2341.730 1393.735 2341.745 ;
        RECT 1393.405 2341.680 1400.700 2341.730 ;
        RECT 1393.405 2341.430 1404.000 2341.680 ;
        RECT 1393.405 2341.415 1393.735 2341.430 ;
        RECT 1400.000 2341.080 1404.000 2341.430 ;
    END
  END la_data_out[0]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 2366.980 662.330 2367.040 ;
        RECT 1393.410 2366.980 1393.730 2367.040 ;
        RECT 662.010 2366.840 1393.730 2366.980 ;
        RECT 662.010 2366.780 662.330 2366.840 ;
        RECT 1393.410 2366.780 1393.730 2366.840 ;
        RECT 656.950 17.920 657.270 17.980 ;
        RECT 662.010 17.920 662.330 17.980 ;
        RECT 656.950 17.780 662.330 17.920 ;
        RECT 656.950 17.720 657.270 17.780 ;
        RECT 662.010 17.720 662.330 17.780 ;
      LAYER via ;
        RECT 662.040 2366.780 662.300 2367.040 ;
        RECT 1393.440 2366.780 1393.700 2367.040 ;
        RECT 656.980 17.720 657.240 17.980 ;
        RECT 662.040 17.720 662.300 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2373.355 1393.710 2373.725 ;
        RECT 1393.500 2367.070 1393.640 2373.355 ;
        RECT 662.040 2366.750 662.300 2367.070 ;
        RECT 1393.440 2366.750 1393.700 2367.070 ;
        RECT 662.100 18.010 662.240 2366.750 ;
        RECT 656.980 17.690 657.240 18.010 ;
        RECT 662.040 17.690 662.300 18.010 ;
        RECT 657.040 2.400 657.180 17.690 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2373.400 1393.710 2373.680 ;
      LAYER met3 ;
        RECT 1393.405 2373.690 1393.735 2373.705 ;
        RECT 1393.405 2373.640 1400.700 2373.690 ;
        RECT 1393.405 2373.390 1404.000 2373.640 ;
        RECT 1393.405 2373.375 1393.735 2373.390 ;
        RECT 1400.000 2373.040 1404.000 2373.390 ;
    END
  END la_data_out[1]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 675.810 2394.860 676.130 2394.920 ;
        RECT 1386.970 2394.860 1387.290 2394.920 ;
        RECT 675.810 2394.720 1387.290 2394.860 ;
        RECT 675.810 2394.660 676.130 2394.720 ;
        RECT 1386.970 2394.660 1387.290 2394.720 ;
      LAYER via ;
        RECT 675.840 2394.660 676.100 2394.920 ;
        RECT 1387.000 2394.660 1387.260 2394.920 ;
      LAYER met2 ;
        RECT 675.840 2394.630 676.100 2394.950 ;
        RECT 1387.000 2394.805 1387.260 2394.950 ;
        RECT 675.900 3.130 676.040 2394.630 ;
        RECT 1386.990 2394.435 1387.270 2394.805 ;
        RECT 674.520 2.990 676.040 3.130 ;
        RECT 674.520 2.400 674.660 2.990 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 1386.990 2394.480 1387.270 2394.760 ;
      LAYER met3 ;
        RECT 1386.965 2394.770 1387.295 2394.785 ;
        RECT 1386.965 2394.720 1400.700 2394.770 ;
        RECT 1386.965 2394.470 1404.000 2394.720 ;
        RECT 1386.965 2394.455 1387.295 2394.470 ;
        RECT 1400.000 2394.120 1404.000 2394.470 ;
    END
  END la_data_out[2]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 2346.240 648.530 2346.300 ;
        RECT 1389.270 2346.240 1389.590 2346.300 ;
        RECT 648.210 2346.100 1389.590 2346.240 ;
        RECT 648.210 2346.040 648.530 2346.100 ;
        RECT 1389.270 2346.040 1389.590 2346.100 ;
        RECT 644.990 17.920 645.310 17.980 ;
        RECT 648.210 17.920 648.530 17.980 ;
        RECT 644.990 17.780 648.530 17.920 ;
        RECT 644.990 17.720 645.310 17.780 ;
        RECT 648.210 17.720 648.530 17.780 ;
      LAYER via ;
        RECT 648.240 2346.040 648.500 2346.300 ;
        RECT 1389.300 2346.040 1389.560 2346.300 ;
        RECT 645.020 17.720 645.280 17.980 ;
        RECT 648.240 17.720 648.500 17.980 ;
      LAYER met2 ;
        RECT 1389.290 2351.595 1389.570 2351.965 ;
        RECT 1389.360 2346.330 1389.500 2351.595 ;
        RECT 648.240 2346.010 648.500 2346.330 ;
        RECT 1389.300 2346.010 1389.560 2346.330 ;
        RECT 648.300 18.010 648.440 2346.010 ;
        RECT 645.020 17.690 645.280 18.010 ;
        RECT 648.240 17.690 648.500 18.010 ;
        RECT 645.080 2.400 645.220 17.690 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 1389.290 2351.640 1389.570 2351.920 ;
      LAYER met3 ;
        RECT 1389.265 2351.930 1389.595 2351.945 ;
        RECT 1389.265 2351.880 1400.700 2351.930 ;
        RECT 1389.265 2351.630 1404.000 2351.880 ;
        RECT 1389.265 2351.615 1389.595 2351.630 ;
        RECT 1400.000 2351.280 1404.000 2351.630 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 2380.580 669.230 2380.640 ;
        RECT 1386.970 2380.580 1387.290 2380.640 ;
        RECT 668.910 2380.440 1387.290 2380.580 ;
        RECT 668.910 2380.380 669.230 2380.440 ;
        RECT 1386.970 2380.380 1387.290 2380.440 ;
        RECT 662.930 17.920 663.250 17.980 ;
        RECT 668.910 17.920 669.230 17.980 ;
        RECT 662.930 17.780 669.230 17.920 ;
        RECT 662.930 17.720 663.250 17.780 ;
        RECT 668.910 17.720 669.230 17.780 ;
      LAYER via ;
        RECT 668.940 2380.380 669.200 2380.640 ;
        RECT 1387.000 2380.380 1387.260 2380.640 ;
        RECT 662.960 17.720 663.220 17.980 ;
        RECT 668.940 17.720 669.200 17.980 ;
      LAYER met2 ;
        RECT 1386.990 2383.555 1387.270 2383.925 ;
        RECT 1387.060 2380.670 1387.200 2383.555 ;
        RECT 668.940 2380.350 669.200 2380.670 ;
        RECT 1387.000 2380.350 1387.260 2380.670 ;
        RECT 669.000 18.010 669.140 2380.350 ;
        RECT 662.960 17.690 663.220 18.010 ;
        RECT 668.940 17.690 669.200 18.010 ;
        RECT 663.020 2.400 663.160 17.690 ;
        RECT 662.810 -4.800 663.370 2.400 ;
      LAYER via2 ;
        RECT 1386.990 2383.600 1387.270 2383.880 ;
      LAYER met3 ;
        RECT 1386.965 2383.890 1387.295 2383.905 ;
        RECT 1386.965 2383.840 1400.700 2383.890 ;
        RECT 1386.965 2383.590 1404.000 2383.840 ;
        RECT 1386.965 2383.575 1387.295 2383.590 ;
        RECT 1400.000 2383.240 1404.000 2383.590 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1518.070 2591.040 1518.390 2591.100 ;
        RECT 2118.370 2591.040 2118.690 2591.100 ;
        RECT 1518.070 2590.900 2118.690 2591.040 ;
        RECT 1518.070 2590.840 1518.390 2590.900 ;
        RECT 2118.370 2590.840 2118.690 2590.900 ;
        RECT 1403.990 2588.320 1404.310 2588.380 ;
        RECT 1518.070 2588.320 1518.390 2588.380 ;
        RECT 1403.990 2588.180 1518.390 2588.320 ;
        RECT 1403.990 2588.120 1404.310 2588.180 ;
        RECT 1518.070 2588.120 1518.390 2588.180 ;
        RECT 1403.990 1203.500 1404.310 1203.560 ;
        RECT 1866.290 1203.500 1866.610 1203.560 ;
        RECT 1403.990 1203.360 1866.610 1203.500 ;
        RECT 1403.990 1203.300 1404.310 1203.360 ;
        RECT 1866.290 1203.300 1866.610 1203.360 ;
        RECT 6.510 1200.780 6.830 1200.840 ;
        RECT 1403.990 1200.780 1404.310 1200.840 ;
        RECT 6.510 1200.640 1404.310 1200.780 ;
        RECT 6.510 1200.580 6.830 1200.640 ;
        RECT 1403.990 1200.580 1404.310 1200.640 ;
        RECT 2.830 17.580 3.150 17.640 ;
        RECT 6.510 17.580 6.830 17.640 ;
        RECT 2.830 17.440 6.830 17.580 ;
        RECT 2.830 17.380 3.150 17.440 ;
        RECT 6.510 17.380 6.830 17.440 ;
      LAYER via ;
        RECT 1518.100 2590.840 1518.360 2591.100 ;
        RECT 2118.400 2590.840 2118.660 2591.100 ;
        RECT 1404.020 2588.120 1404.280 2588.380 ;
        RECT 1518.100 2588.120 1518.360 2588.380 ;
        RECT 1404.020 1203.300 1404.280 1203.560 ;
        RECT 1866.320 1203.300 1866.580 1203.560 ;
        RECT 6.540 1200.580 6.800 1200.840 ;
        RECT 1404.020 1200.580 1404.280 1200.840 ;
        RECT 2.860 17.380 3.120 17.640 ;
        RECT 6.540 17.380 6.800 17.640 ;
      LAYER met2 ;
        RECT 1518.090 2592.315 1518.370 2592.685 ;
        RECT 1518.160 2591.130 1518.300 2592.315 ;
        RECT 1518.100 2590.810 1518.360 2591.130 ;
        RECT 2118.390 2590.955 2118.670 2591.325 ;
        RECT 2118.400 2590.810 2118.660 2590.955 ;
        RECT 1518.160 2588.410 1518.300 2590.810 ;
        RECT 1404.020 2588.090 1404.280 2588.410 ;
        RECT 1518.100 2588.090 1518.360 2588.410 ;
        RECT 1404.080 1204.125 1404.220 2588.090 ;
        RECT 1404.010 1203.755 1404.290 1204.125 ;
        RECT 1404.080 1203.590 1404.220 1203.755 ;
        RECT 1404.020 1203.270 1404.280 1203.590 ;
        RECT 1866.320 1203.270 1866.580 1203.590 ;
        RECT 1404.080 1200.870 1404.220 1203.270 ;
        RECT 6.540 1200.550 6.800 1200.870 ;
        RECT 1404.020 1200.550 1404.280 1200.870 ;
        RECT 6.600 17.670 6.740 1200.550 ;
        RECT 1866.380 1015.765 1866.520 1203.270 ;
        RECT 1866.310 1015.395 1866.590 1015.765 ;
        RECT 2.860 17.350 3.120 17.670 ;
        RECT 6.540 17.350 6.800 17.670 ;
        RECT 2.920 2.400 3.060 17.350 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 1518.090 2592.360 1518.370 2592.640 ;
        RECT 2118.390 2591.000 2118.670 2591.280 ;
        RECT 1404.010 1203.800 1404.290 1204.080 ;
        RECT 1866.310 1015.440 1866.590 1015.720 ;
      LAYER met3 ;
        RECT 1518.065 2592.660 1518.395 2592.665 ;
        RECT 1518.065 2592.650 1518.650 2592.660 ;
        RECT 1518.065 2592.350 1518.850 2592.650 ;
        RECT 1518.065 2592.340 1518.650 2592.350 ;
        RECT 1518.065 2592.335 1518.395 2592.340 ;
        RECT 2118.365 2591.290 2118.695 2591.305 ;
        RECT 2119.030 2591.290 2119.410 2591.300 ;
        RECT 2118.365 2590.990 2119.410 2591.290 ;
        RECT 2118.365 2590.975 2118.695 2590.990 ;
        RECT 2119.030 2590.980 2119.410 2590.990 ;
        RECT 1400.000 1204.800 1404.000 1205.400 ;
        RECT 1403.310 1204.090 1403.610 1204.800 ;
        RECT 1403.985 1204.090 1404.315 1204.105 ;
        RECT 1403.310 1203.790 1404.315 1204.090 ;
        RECT 1403.985 1203.775 1404.315 1203.790 ;
        RECT 1866.285 1015.730 1866.615 1015.745 ;
        RECT 1866.950 1015.730 1867.330 1015.740 ;
        RECT 2464.030 1015.730 2464.410 1015.740 ;
        RECT 1866.285 1015.430 2464.410 1015.730 ;
        RECT 1866.285 1015.415 1866.615 1015.430 ;
        RECT 1866.950 1015.420 1867.330 1015.430 ;
        RECT 2464.030 1015.420 2464.410 1015.430 ;
      LAYER via3 ;
        RECT 1518.300 2592.340 1518.620 2592.660 ;
        RECT 2119.060 2590.980 2119.380 2591.300 ;
        RECT 1866.980 1015.420 1867.300 1015.740 ;
        RECT 2464.060 1015.420 2464.380 1015.740 ;
      LAYER met4 ;
        RECT 1519.015 2601.150 1519.315 2604.600 ;
        RECT 1518.310 2600.850 1519.315 2601.150 ;
        RECT 1518.310 2592.665 1518.610 2600.850 ;
        RECT 1519.015 2600.000 1519.315 2600.850 ;
        RECT 2119.015 2601.150 2119.315 2604.600 ;
        RECT 2119.015 2600.000 2119.370 2601.150 ;
        RECT 1518.295 2592.335 1518.625 2592.665 ;
        RECT 2119.070 2591.305 2119.370 2600.000 ;
        RECT 2119.055 2590.975 2119.385 2591.305 ;
        RECT 1866.975 1015.415 1867.305 1015.745 ;
        RECT 2464.055 1015.415 2464.385 1015.745 ;
        RECT 1866.990 1006.235 1867.290 1015.415 ;
        RECT 1866.990 1004.550 1867.465 1006.235 ;
        RECT 2464.070 1004.850 2464.370 1015.415 ;
        RECT 2467.165 1004.850 2467.465 1006.235 ;
        RECT 2464.070 1004.550 2467.465 1004.850 ;
        RECT 1867.165 1001.635 1867.465 1004.550 ;
        RECT 2467.165 1001.635 2467.465 1004.550 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.410 1214.720 13.730 1214.780 ;
        RECT 1393.410 1214.720 1393.730 1214.780 ;
        RECT 13.410 1214.580 1393.730 1214.720 ;
        RECT 13.410 1214.520 13.730 1214.580 ;
        RECT 1393.410 1214.520 1393.730 1214.580 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 13.410 17.580 13.730 17.640 ;
        RECT 8.350 17.440 13.730 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 13.410 17.380 13.730 17.440 ;
      LAYER via ;
        RECT 13.440 1214.520 13.700 1214.780 ;
        RECT 1393.440 1214.520 1393.700 1214.780 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 13.440 17.380 13.700 17.640 ;
      LAYER met2 ;
        RECT 1393.430 1215.315 1393.710 1215.685 ;
        RECT 1393.500 1214.810 1393.640 1215.315 ;
        RECT 13.440 1214.490 13.700 1214.810 ;
        RECT 1393.440 1214.490 1393.700 1214.810 ;
        RECT 13.500 17.670 13.640 1214.490 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 13.440 17.350 13.700 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1215.360 1393.710 1215.640 ;
      LAYER met3 ;
        RECT 1393.405 1215.650 1393.735 1215.665 ;
        RECT 1393.405 1215.600 1400.700 1215.650 ;
        RECT 1393.405 1215.350 1404.000 1215.600 ;
        RECT 1393.405 1215.335 1393.735 1215.350 ;
        RECT 1400.000 1215.000 1404.000 1215.350 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 17.580 14.650 17.640 ;
        RECT 1390.650 17.580 1390.970 17.640 ;
        RECT 14.330 17.440 1390.970 17.580 ;
        RECT 14.330 17.380 14.650 17.440 ;
        RECT 1390.650 17.380 1390.970 17.440 ;
      LAYER via ;
        RECT 14.360 17.380 14.620 17.640 ;
        RECT 1390.680 17.380 1390.940 17.640 ;
      LAYER met2 ;
        RECT 1390.670 1226.195 1390.950 1226.565 ;
        RECT 1390.740 17.670 1390.880 1226.195 ;
        RECT 14.360 17.350 14.620 17.670 ;
        RECT 1390.680 17.350 1390.940 17.670 ;
        RECT 14.420 2.400 14.560 17.350 ;
        RECT 14.210 -4.800 14.770 2.400 ;
      LAYER via2 ;
        RECT 1390.670 1226.240 1390.950 1226.520 ;
      LAYER met3 ;
        RECT 1390.645 1226.530 1390.975 1226.545 ;
        RECT 1390.645 1226.480 1400.700 1226.530 ;
        RECT 1390.645 1226.230 1404.000 1226.480 ;
        RECT 1390.645 1226.215 1390.975 1226.230 ;
        RECT 1400.000 1225.880 1404.000 1226.230 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 41.010 1263.000 41.330 1263.060 ;
        RECT 1389.270 1263.000 1389.590 1263.060 ;
        RECT 41.010 1262.860 1389.590 1263.000 ;
        RECT 41.010 1262.800 41.330 1262.860 ;
        RECT 1389.270 1262.800 1389.590 1262.860 ;
        RECT 38.250 17.920 38.570 17.980 ;
        RECT 41.010 17.920 41.330 17.980 ;
        RECT 38.250 17.780 41.330 17.920 ;
        RECT 38.250 17.720 38.570 17.780 ;
        RECT 41.010 17.720 41.330 17.780 ;
      LAYER via ;
        RECT 41.040 1262.800 41.300 1263.060 ;
        RECT 1389.300 1262.800 1389.560 1263.060 ;
        RECT 38.280 17.720 38.540 17.980 ;
        RECT 41.040 17.720 41.300 17.980 ;
      LAYER met2 ;
        RECT 1389.290 1268.355 1389.570 1268.725 ;
        RECT 1389.360 1263.090 1389.500 1268.355 ;
        RECT 41.040 1262.770 41.300 1263.090 ;
        RECT 1389.300 1262.770 1389.560 1263.090 ;
        RECT 41.100 18.010 41.240 1262.770 ;
        RECT 38.280 17.690 38.540 18.010 ;
        RECT 41.040 17.690 41.300 18.010 ;
        RECT 38.340 2.400 38.480 17.690 ;
        RECT 38.130 -4.800 38.690 2.400 ;
      LAYER via2 ;
        RECT 1389.290 1268.400 1389.570 1268.680 ;
      LAYER met3 ;
        RECT 1389.265 1268.690 1389.595 1268.705 ;
        RECT 1389.265 1268.640 1400.700 1268.690 ;
        RECT 1389.265 1268.390 1404.000 1268.640 ;
        RECT 1389.265 1268.375 1389.595 1268.390 ;
        RECT 1400.000 1268.040 1404.000 1268.390 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 1628.500 241.430 1628.560 ;
        RECT 1390.190 1628.500 1390.510 1628.560 ;
        RECT 241.110 1628.360 1390.510 1628.500 ;
        RECT 241.110 1628.300 241.430 1628.360 ;
        RECT 1390.190 1628.300 1390.510 1628.360 ;
      LAYER via ;
        RECT 241.140 1628.300 241.400 1628.560 ;
        RECT 1390.220 1628.300 1390.480 1628.560 ;
      LAYER met2 ;
        RECT 1390.210 1629.435 1390.490 1629.805 ;
        RECT 1390.280 1628.590 1390.420 1629.435 ;
        RECT 241.140 1628.270 241.400 1628.590 ;
        RECT 1390.220 1628.270 1390.480 1628.590 ;
        RECT 241.200 17.410 241.340 1628.270 ;
        RECT 240.740 17.270 241.340 17.410 ;
        RECT 240.740 2.400 240.880 17.270 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 1390.210 1629.480 1390.490 1629.760 ;
      LAYER met3 ;
        RECT 1390.185 1629.770 1390.515 1629.785 ;
        RECT 1390.185 1629.720 1400.700 1629.770 ;
        RECT 1390.185 1629.470 1404.000 1629.720 ;
        RECT 1390.185 1629.455 1390.515 1629.470 ;
        RECT 1400.000 1629.120 1404.000 1629.470 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 261.810 1656.380 262.130 1656.440 ;
        RECT 1393.410 1656.380 1393.730 1656.440 ;
        RECT 261.810 1656.240 1393.730 1656.380 ;
        RECT 261.810 1656.180 262.130 1656.240 ;
        RECT 1393.410 1656.180 1393.730 1656.240 ;
        RECT 258.130 17.920 258.450 17.980 ;
        RECT 261.810 17.920 262.130 17.980 ;
        RECT 258.130 17.780 262.130 17.920 ;
        RECT 258.130 17.720 258.450 17.780 ;
        RECT 261.810 17.720 262.130 17.780 ;
      LAYER via ;
        RECT 261.840 1656.180 262.100 1656.440 ;
        RECT 1393.440 1656.180 1393.700 1656.440 ;
        RECT 258.160 17.720 258.420 17.980 ;
        RECT 261.840 17.720 262.100 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1661.395 1393.710 1661.765 ;
        RECT 1393.500 1656.470 1393.640 1661.395 ;
        RECT 261.840 1656.150 262.100 1656.470 ;
        RECT 1393.440 1656.150 1393.700 1656.470 ;
        RECT 261.900 18.010 262.040 1656.150 ;
        RECT 258.160 17.690 258.420 18.010 ;
        RECT 261.840 17.690 262.100 18.010 ;
        RECT 258.220 2.400 258.360 17.690 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1661.440 1393.710 1661.720 ;
      LAYER met3 ;
        RECT 1393.405 1661.730 1393.735 1661.745 ;
        RECT 1393.405 1661.680 1400.700 1661.730 ;
        RECT 1393.405 1661.430 1404.000 1661.680 ;
        RECT 1393.405 1661.415 1393.735 1661.430 ;
        RECT 1400.000 1661.080 1404.000 1661.430 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 1690.720 282.370 1690.780 ;
        RECT 1393.410 1690.720 1393.730 1690.780 ;
        RECT 282.050 1690.580 1393.730 1690.720 ;
        RECT 282.050 1690.520 282.370 1690.580 ;
        RECT 1393.410 1690.520 1393.730 1690.580 ;
        RECT 276.070 17.920 276.390 17.980 ;
        RECT 282.050 17.920 282.370 17.980 ;
        RECT 276.070 17.780 282.370 17.920 ;
        RECT 276.070 17.720 276.390 17.780 ;
        RECT 282.050 17.720 282.370 17.780 ;
      LAYER via ;
        RECT 282.080 1690.520 282.340 1690.780 ;
        RECT 1393.440 1690.520 1393.700 1690.780 ;
        RECT 276.100 17.720 276.360 17.980 ;
        RECT 282.080 17.720 282.340 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1693.355 1393.710 1693.725 ;
        RECT 1393.500 1690.810 1393.640 1693.355 ;
        RECT 282.080 1690.490 282.340 1690.810 ;
        RECT 1393.440 1690.490 1393.700 1690.810 ;
        RECT 282.140 18.010 282.280 1690.490 ;
        RECT 276.100 17.690 276.360 18.010 ;
        RECT 282.080 17.690 282.340 18.010 ;
        RECT 276.160 2.400 276.300 17.690 ;
        RECT 275.950 -4.800 276.510 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1693.400 1393.710 1693.680 ;
      LAYER met3 ;
        RECT 1393.405 1693.690 1393.735 1693.705 ;
        RECT 1393.405 1693.640 1400.700 1693.690 ;
        RECT 1393.405 1693.390 1404.000 1693.640 ;
        RECT 1393.405 1693.375 1393.735 1693.390 ;
        RECT 1400.000 1693.040 1404.000 1693.390 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 296.310 1725.400 296.630 1725.460 ;
        RECT 1393.410 1725.400 1393.730 1725.460 ;
        RECT 296.310 1725.260 1393.730 1725.400 ;
        RECT 296.310 1725.200 296.630 1725.260 ;
        RECT 1393.410 1725.200 1393.730 1725.260 ;
        RECT 294.010 17.920 294.330 17.980 ;
        RECT 296.310 17.920 296.630 17.980 ;
        RECT 294.010 17.780 296.630 17.920 ;
        RECT 294.010 17.720 294.330 17.780 ;
        RECT 296.310 17.720 296.630 17.780 ;
      LAYER via ;
        RECT 296.340 1725.200 296.600 1725.460 ;
        RECT 1393.440 1725.200 1393.700 1725.460 ;
        RECT 294.040 17.720 294.300 17.980 ;
        RECT 296.340 17.720 296.600 17.980 ;
      LAYER met2 ;
        RECT 296.340 1725.170 296.600 1725.490 ;
        RECT 1393.430 1725.315 1393.710 1725.685 ;
        RECT 1393.440 1725.170 1393.700 1725.315 ;
        RECT 296.400 18.010 296.540 1725.170 ;
        RECT 294.040 17.690 294.300 18.010 ;
        RECT 296.340 17.690 296.600 18.010 ;
        RECT 294.100 2.400 294.240 17.690 ;
        RECT 293.890 -4.800 294.450 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1725.360 1393.710 1725.640 ;
      LAYER met3 ;
        RECT 1393.405 1725.650 1393.735 1725.665 ;
        RECT 1393.405 1725.600 1400.700 1725.650 ;
        RECT 1393.405 1725.350 1404.000 1725.600 ;
        RECT 1393.405 1725.335 1393.735 1725.350 ;
        RECT 1400.000 1725.000 1404.000 1725.350 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.010 1752.940 317.330 1753.000 ;
        RECT 1393.410 1752.940 1393.730 1753.000 ;
        RECT 317.010 1752.800 1393.730 1752.940 ;
        RECT 317.010 1752.740 317.330 1752.800 ;
        RECT 1393.410 1752.740 1393.730 1752.800 ;
        RECT 311.950 15.880 312.270 15.940 ;
        RECT 317.010 15.880 317.330 15.940 ;
        RECT 311.950 15.740 317.330 15.880 ;
        RECT 311.950 15.680 312.270 15.740 ;
        RECT 317.010 15.680 317.330 15.740 ;
      LAYER via ;
        RECT 317.040 1752.740 317.300 1753.000 ;
        RECT 1393.440 1752.740 1393.700 1753.000 ;
        RECT 311.980 15.680 312.240 15.940 ;
        RECT 317.040 15.680 317.300 15.940 ;
      LAYER met2 ;
        RECT 1393.430 1757.275 1393.710 1757.645 ;
        RECT 1393.500 1753.030 1393.640 1757.275 ;
        RECT 317.040 1752.710 317.300 1753.030 ;
        RECT 1393.440 1752.710 1393.700 1753.030 ;
        RECT 317.100 15.970 317.240 1752.710 ;
        RECT 311.980 15.650 312.240 15.970 ;
        RECT 317.040 15.650 317.300 15.970 ;
        RECT 312.040 2.400 312.180 15.650 ;
        RECT 311.830 -4.800 312.390 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1757.320 1393.710 1757.600 ;
      LAYER met3 ;
        RECT 1393.405 1757.610 1393.735 1757.625 ;
        RECT 1393.405 1757.560 1400.700 1757.610 ;
        RECT 1393.405 1757.310 1404.000 1757.560 ;
        RECT 1393.405 1757.295 1393.735 1757.310 ;
        RECT 1400.000 1756.960 1404.000 1757.310 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 330.810 1787.280 331.130 1787.340 ;
        RECT 1393.410 1787.280 1393.730 1787.340 ;
        RECT 330.810 1787.140 1393.730 1787.280 ;
        RECT 330.810 1787.080 331.130 1787.140 ;
        RECT 1393.410 1787.080 1393.730 1787.140 ;
      LAYER via ;
        RECT 330.840 1787.080 331.100 1787.340 ;
        RECT 1393.440 1787.080 1393.700 1787.340 ;
      LAYER met2 ;
        RECT 1393.430 1789.235 1393.710 1789.605 ;
        RECT 1393.500 1787.370 1393.640 1789.235 ;
        RECT 330.840 1787.050 331.100 1787.370 ;
        RECT 1393.440 1787.050 1393.700 1787.370 ;
        RECT 330.900 17.410 331.040 1787.050 ;
        RECT 329.980 17.270 331.040 17.410 ;
        RECT 329.980 2.400 330.120 17.270 ;
        RECT 329.770 -4.800 330.330 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1789.280 1393.710 1789.560 ;
      LAYER met3 ;
        RECT 1393.405 1789.570 1393.735 1789.585 ;
        RECT 1393.405 1789.520 1400.700 1789.570 ;
        RECT 1393.405 1789.270 1404.000 1789.520 ;
        RECT 1393.405 1789.255 1393.735 1789.270 ;
        RECT 1400.000 1788.920 1404.000 1789.270 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 351.510 1814.820 351.830 1814.880 ;
        RECT 1389.270 1814.820 1389.590 1814.880 ;
        RECT 351.510 1814.680 1389.590 1814.820 ;
        RECT 351.510 1814.620 351.830 1814.680 ;
        RECT 1389.270 1814.620 1389.590 1814.680 ;
        RECT 347.370 17.920 347.690 17.980 ;
        RECT 351.510 17.920 351.830 17.980 ;
        RECT 347.370 17.780 351.830 17.920 ;
        RECT 347.370 17.720 347.690 17.780 ;
        RECT 351.510 17.720 351.830 17.780 ;
      LAYER via ;
        RECT 351.540 1814.620 351.800 1814.880 ;
        RECT 1389.300 1814.620 1389.560 1814.880 ;
        RECT 347.400 17.720 347.660 17.980 ;
        RECT 351.540 17.720 351.800 17.980 ;
      LAYER met2 ;
        RECT 1389.290 1820.515 1389.570 1820.885 ;
        RECT 1389.360 1814.910 1389.500 1820.515 ;
        RECT 351.540 1814.590 351.800 1814.910 ;
        RECT 1389.300 1814.590 1389.560 1814.910 ;
        RECT 351.600 18.010 351.740 1814.590 ;
        RECT 347.400 17.690 347.660 18.010 ;
        RECT 351.540 17.690 351.800 18.010 ;
        RECT 347.460 2.400 347.600 17.690 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 1389.290 1820.560 1389.570 1820.840 ;
      LAYER met3 ;
        RECT 1389.265 1820.850 1389.595 1820.865 ;
        RECT 1389.265 1820.800 1400.700 1820.850 ;
        RECT 1389.265 1820.550 1404.000 1820.800 ;
        RECT 1389.265 1820.535 1389.595 1820.550 ;
        RECT 1400.000 1820.200 1404.000 1820.550 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 1849.500 365.630 1849.560 ;
        RECT 1391.570 1849.500 1391.890 1849.560 ;
        RECT 365.310 1849.360 1391.890 1849.500 ;
        RECT 365.310 1849.300 365.630 1849.360 ;
        RECT 1391.570 1849.300 1391.890 1849.360 ;
      LAYER via ;
        RECT 365.340 1849.300 365.600 1849.560 ;
        RECT 1391.600 1849.300 1391.860 1849.560 ;
      LAYER met2 ;
        RECT 1391.590 1852.475 1391.870 1852.845 ;
        RECT 1391.660 1849.590 1391.800 1852.475 ;
        RECT 365.340 1849.270 365.600 1849.590 ;
        RECT 1391.600 1849.270 1391.860 1849.590 ;
        RECT 365.400 2.400 365.540 1849.270 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 1391.590 1852.520 1391.870 1852.800 ;
      LAYER met3 ;
        RECT 1391.565 1852.810 1391.895 1852.825 ;
        RECT 1391.565 1852.760 1400.700 1852.810 ;
        RECT 1391.565 1852.510 1404.000 1852.760 ;
        RECT 1391.565 1852.495 1391.895 1852.510 ;
        RECT 1400.000 1852.160 1404.000 1852.510 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 386.010 1883.840 386.330 1883.900 ;
        RECT 1393.410 1883.840 1393.730 1883.900 ;
        RECT 386.010 1883.700 1393.730 1883.840 ;
        RECT 386.010 1883.640 386.330 1883.700 ;
        RECT 1393.410 1883.640 1393.730 1883.700 ;
        RECT 383.250 17.920 383.570 17.980 ;
        RECT 386.010 17.920 386.330 17.980 ;
        RECT 383.250 17.780 386.330 17.920 ;
        RECT 383.250 17.720 383.570 17.780 ;
        RECT 386.010 17.720 386.330 17.780 ;
      LAYER via ;
        RECT 386.040 1883.640 386.300 1883.900 ;
        RECT 1393.440 1883.640 1393.700 1883.900 ;
        RECT 383.280 17.720 383.540 17.980 ;
        RECT 386.040 17.720 386.300 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1884.435 1393.710 1884.805 ;
        RECT 1393.500 1883.930 1393.640 1884.435 ;
        RECT 386.040 1883.610 386.300 1883.930 ;
        RECT 1393.440 1883.610 1393.700 1883.930 ;
        RECT 386.100 18.010 386.240 1883.610 ;
        RECT 383.280 17.690 383.540 18.010 ;
        RECT 386.040 17.690 386.300 18.010 ;
        RECT 383.340 2.400 383.480 17.690 ;
        RECT 383.130 -4.800 383.690 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1884.480 1393.710 1884.760 ;
      LAYER met3 ;
        RECT 1393.405 1884.770 1393.735 1884.785 ;
        RECT 1393.405 1884.720 1400.700 1884.770 ;
        RECT 1393.405 1884.470 1404.000 1884.720 ;
        RECT 1393.405 1884.455 1393.735 1884.470 ;
        RECT 1400.000 1884.120 1404.000 1884.470 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 406.710 1911.380 407.030 1911.440 ;
        RECT 1393.410 1911.380 1393.730 1911.440 ;
        RECT 406.710 1911.240 1393.730 1911.380 ;
        RECT 406.710 1911.180 407.030 1911.240 ;
        RECT 1393.410 1911.180 1393.730 1911.240 ;
        RECT 401.190 17.920 401.510 17.980 ;
        RECT 406.710 17.920 407.030 17.980 ;
        RECT 401.190 17.780 407.030 17.920 ;
        RECT 401.190 17.720 401.510 17.780 ;
        RECT 406.710 17.720 407.030 17.780 ;
      LAYER via ;
        RECT 406.740 1911.180 407.000 1911.440 ;
        RECT 1393.440 1911.180 1393.700 1911.440 ;
        RECT 401.220 17.720 401.480 17.980 ;
        RECT 406.740 17.720 407.000 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1916.395 1393.710 1916.765 ;
        RECT 1393.500 1911.470 1393.640 1916.395 ;
        RECT 406.740 1911.150 407.000 1911.470 ;
        RECT 1393.440 1911.150 1393.700 1911.470 ;
        RECT 406.800 18.010 406.940 1911.150 ;
        RECT 401.220 17.690 401.480 18.010 ;
        RECT 406.740 17.690 407.000 18.010 ;
        RECT 401.280 2.400 401.420 17.690 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1916.440 1393.710 1916.720 ;
      LAYER met3 ;
        RECT 1393.405 1916.730 1393.735 1916.745 ;
        RECT 1393.405 1916.680 1400.700 1916.730 ;
        RECT 1393.405 1916.430 1404.000 1916.680 ;
        RECT 1393.405 1916.415 1393.735 1916.430 ;
        RECT 1400.000 1916.080 1404.000 1916.430 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 1311.280 68.470 1311.340 ;
        RECT 1393.410 1311.280 1393.730 1311.340 ;
        RECT 68.150 1311.140 1393.730 1311.280 ;
        RECT 68.150 1311.080 68.470 1311.140 ;
        RECT 1393.410 1311.080 1393.730 1311.140 ;
        RECT 62.170 17.920 62.490 17.980 ;
        RECT 68.150 17.920 68.470 17.980 ;
        RECT 62.170 17.780 68.470 17.920 ;
        RECT 62.170 17.720 62.490 17.780 ;
        RECT 68.150 17.720 68.470 17.780 ;
      LAYER via ;
        RECT 68.180 1311.080 68.440 1311.340 ;
        RECT 1393.440 1311.080 1393.700 1311.340 ;
        RECT 62.200 17.720 62.460 17.980 ;
        RECT 68.180 17.720 68.440 17.980 ;
      LAYER met2 ;
        RECT 68.180 1311.050 68.440 1311.370 ;
        RECT 1393.430 1311.195 1393.710 1311.565 ;
        RECT 1393.440 1311.050 1393.700 1311.195 ;
        RECT 68.240 18.010 68.380 1311.050 ;
        RECT 62.200 17.690 62.460 18.010 ;
        RECT 68.180 17.690 68.440 18.010 ;
        RECT 62.260 2.400 62.400 17.690 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1311.240 1393.710 1311.520 ;
      LAYER met3 ;
        RECT 1393.405 1311.530 1393.735 1311.545 ;
        RECT 1393.405 1311.480 1400.700 1311.530 ;
        RECT 1393.405 1311.230 1404.000 1311.480 ;
        RECT 1393.405 1311.215 1393.735 1311.230 ;
        RECT 1400.000 1310.880 1404.000 1311.230 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 420.510 1946.060 420.830 1946.120 ;
        RECT 1393.410 1946.060 1393.730 1946.120 ;
        RECT 420.510 1945.920 1393.730 1946.060 ;
        RECT 420.510 1945.860 420.830 1945.920 ;
        RECT 1393.410 1945.860 1393.730 1945.920 ;
      LAYER via ;
        RECT 420.540 1945.860 420.800 1946.120 ;
        RECT 1393.440 1945.860 1393.700 1946.120 ;
      LAYER met2 ;
        RECT 1393.430 1948.355 1393.710 1948.725 ;
        RECT 1393.500 1946.150 1393.640 1948.355 ;
        RECT 420.540 1945.830 420.800 1946.150 ;
        RECT 1393.440 1945.830 1393.700 1946.150 ;
        RECT 420.600 17.410 420.740 1945.830 ;
        RECT 419.220 17.270 420.740 17.410 ;
        RECT 419.220 2.400 419.360 17.270 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1948.400 1393.710 1948.680 ;
      LAYER met3 ;
        RECT 1393.405 1948.690 1393.735 1948.705 ;
        RECT 1393.405 1948.640 1400.700 1948.690 ;
        RECT 1393.405 1948.390 1404.000 1948.640 ;
        RECT 1393.405 1948.375 1393.735 1948.390 ;
        RECT 1400.000 1948.040 1404.000 1948.390 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 441.210 1980.400 441.530 1980.460 ;
        RECT 1393.410 1980.400 1393.730 1980.460 ;
        RECT 441.210 1980.260 1393.730 1980.400 ;
        RECT 441.210 1980.200 441.530 1980.260 ;
        RECT 1393.410 1980.200 1393.730 1980.260 ;
        RECT 436.610 17.920 436.930 17.980 ;
        RECT 441.210 17.920 441.530 17.980 ;
        RECT 436.610 17.780 441.530 17.920 ;
        RECT 436.610 17.720 436.930 17.780 ;
        RECT 441.210 17.720 441.530 17.780 ;
      LAYER via ;
        RECT 441.240 1980.200 441.500 1980.460 ;
        RECT 1393.440 1980.200 1393.700 1980.460 ;
        RECT 436.640 17.720 436.900 17.980 ;
        RECT 441.240 17.720 441.500 17.980 ;
      LAYER met2 ;
        RECT 441.240 1980.170 441.500 1980.490 ;
        RECT 1393.430 1980.315 1393.710 1980.685 ;
        RECT 1393.440 1980.170 1393.700 1980.315 ;
        RECT 441.300 18.010 441.440 1980.170 ;
        RECT 436.640 17.690 436.900 18.010 ;
        RECT 441.240 17.690 441.500 18.010 ;
        RECT 436.700 2.400 436.840 17.690 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1980.360 1393.710 1980.640 ;
      LAYER met3 ;
        RECT 1393.405 1980.650 1393.735 1980.665 ;
        RECT 1393.405 1980.600 1400.700 1980.650 ;
        RECT 1393.405 1980.350 1404.000 1980.600 ;
        RECT 1393.405 1980.335 1393.735 1980.350 ;
        RECT 1400.000 1980.000 1404.000 1980.350 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 455.010 2008.280 455.330 2008.340 ;
        RECT 1392.030 2008.280 1392.350 2008.340 ;
        RECT 455.010 2008.140 1392.350 2008.280 ;
        RECT 455.010 2008.080 455.330 2008.140 ;
        RECT 1392.030 2008.080 1392.350 2008.140 ;
      LAYER via ;
        RECT 455.040 2008.080 455.300 2008.340 ;
        RECT 1392.060 2008.080 1392.320 2008.340 ;
      LAYER met2 ;
        RECT 1392.050 2012.275 1392.330 2012.645 ;
        RECT 1392.120 2008.370 1392.260 2012.275 ;
        RECT 455.040 2008.050 455.300 2008.370 ;
        RECT 1392.060 2008.050 1392.320 2008.370 ;
        RECT 455.100 17.410 455.240 2008.050 ;
        RECT 454.640 17.270 455.240 17.410 ;
        RECT 454.640 2.400 454.780 17.270 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 1392.050 2012.320 1392.330 2012.600 ;
      LAYER met3 ;
        RECT 1392.025 2012.610 1392.355 2012.625 ;
        RECT 1392.025 2012.560 1400.700 2012.610 ;
        RECT 1392.025 2012.310 1404.000 2012.560 ;
        RECT 1392.025 2012.295 1392.355 2012.310 ;
        RECT 1400.000 2011.960 1404.000 2012.310 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 475.710 2042.620 476.030 2042.680 ;
        RECT 1393.410 2042.620 1393.730 2042.680 ;
        RECT 475.710 2042.480 1393.730 2042.620 ;
        RECT 475.710 2042.420 476.030 2042.480 ;
        RECT 1393.410 2042.420 1393.730 2042.480 ;
        RECT 472.490 17.920 472.810 17.980 ;
        RECT 475.710 17.920 476.030 17.980 ;
        RECT 472.490 17.780 476.030 17.920 ;
        RECT 472.490 17.720 472.810 17.780 ;
        RECT 475.710 17.720 476.030 17.780 ;
      LAYER via ;
        RECT 475.740 2042.420 476.000 2042.680 ;
        RECT 1393.440 2042.420 1393.700 2042.680 ;
        RECT 472.520 17.720 472.780 17.980 ;
        RECT 475.740 17.720 476.000 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2043.555 1393.710 2043.925 ;
        RECT 1393.500 2042.710 1393.640 2043.555 ;
        RECT 475.740 2042.390 476.000 2042.710 ;
        RECT 1393.440 2042.390 1393.700 2042.710 ;
        RECT 475.800 18.010 475.940 2042.390 ;
        RECT 472.520 17.690 472.780 18.010 ;
        RECT 475.740 17.690 476.000 18.010 ;
        RECT 472.580 2.400 472.720 17.690 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2043.600 1393.710 2043.880 ;
      LAYER met3 ;
        RECT 1393.405 2043.890 1393.735 2043.905 ;
        RECT 1393.405 2043.840 1400.700 2043.890 ;
        RECT 1393.405 2043.590 1404.000 2043.840 ;
        RECT 1393.405 2043.575 1393.735 2043.590 ;
        RECT 1400.000 2043.240 1404.000 2043.590 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 495.950 2070.160 496.270 2070.220 ;
        RECT 1389.270 2070.160 1389.590 2070.220 ;
        RECT 495.950 2070.020 1389.590 2070.160 ;
        RECT 495.950 2069.960 496.270 2070.020 ;
        RECT 1389.270 2069.960 1389.590 2070.020 ;
        RECT 490.430 17.920 490.750 17.980 ;
        RECT 495.950 17.920 496.270 17.980 ;
        RECT 490.430 17.780 496.270 17.920 ;
        RECT 490.430 17.720 490.750 17.780 ;
        RECT 495.950 17.720 496.270 17.780 ;
      LAYER via ;
        RECT 495.980 2069.960 496.240 2070.220 ;
        RECT 1389.300 2069.960 1389.560 2070.220 ;
        RECT 490.460 17.720 490.720 17.980 ;
        RECT 495.980 17.720 496.240 17.980 ;
      LAYER met2 ;
        RECT 1389.290 2075.515 1389.570 2075.885 ;
        RECT 1389.360 2070.250 1389.500 2075.515 ;
        RECT 495.980 2069.930 496.240 2070.250 ;
        RECT 1389.300 2069.930 1389.560 2070.250 ;
        RECT 496.040 18.010 496.180 2069.930 ;
        RECT 490.460 17.690 490.720 18.010 ;
        RECT 495.980 17.690 496.240 18.010 ;
        RECT 490.520 2.400 490.660 17.690 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 1389.290 2075.560 1389.570 2075.840 ;
      LAYER met3 ;
        RECT 1389.265 2075.850 1389.595 2075.865 ;
        RECT 1389.265 2075.800 1400.700 2075.850 ;
        RECT 1389.265 2075.550 1404.000 2075.800 ;
        RECT 1389.265 2075.535 1389.595 2075.550 ;
        RECT 1400.000 2075.200 1404.000 2075.550 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 510.210 2104.840 510.530 2104.900 ;
        RECT 1393.410 2104.840 1393.730 2104.900 ;
        RECT 510.210 2104.700 1393.730 2104.840 ;
        RECT 510.210 2104.640 510.530 2104.700 ;
        RECT 1393.410 2104.640 1393.730 2104.700 ;
        RECT 507.910 16.560 508.230 16.620 ;
        RECT 510.210 16.560 510.530 16.620 ;
        RECT 507.910 16.420 510.530 16.560 ;
        RECT 507.910 16.360 508.230 16.420 ;
        RECT 510.210 16.360 510.530 16.420 ;
      LAYER via ;
        RECT 510.240 2104.640 510.500 2104.900 ;
        RECT 1393.440 2104.640 1393.700 2104.900 ;
        RECT 507.940 16.360 508.200 16.620 ;
        RECT 510.240 16.360 510.500 16.620 ;
      LAYER met2 ;
        RECT 1393.430 2107.475 1393.710 2107.845 ;
        RECT 1393.500 2104.930 1393.640 2107.475 ;
        RECT 510.240 2104.610 510.500 2104.930 ;
        RECT 1393.440 2104.610 1393.700 2104.930 ;
        RECT 510.300 16.650 510.440 2104.610 ;
        RECT 507.940 16.330 508.200 16.650 ;
        RECT 510.240 16.330 510.500 16.650 ;
        RECT 508.000 2.400 508.140 16.330 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2107.520 1393.710 2107.800 ;
      LAYER met3 ;
        RECT 1393.405 2107.810 1393.735 2107.825 ;
        RECT 1393.405 2107.760 1400.700 2107.810 ;
        RECT 1393.405 2107.510 1404.000 2107.760 ;
        RECT 1393.405 2107.495 1393.735 2107.510 ;
        RECT 1400.000 2107.160 1404.000 2107.510 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 530.910 2139.180 531.230 2139.240 ;
        RECT 1393.410 2139.180 1393.730 2139.240 ;
        RECT 530.910 2139.040 1393.730 2139.180 ;
        RECT 530.910 2138.980 531.230 2139.040 ;
        RECT 1393.410 2138.980 1393.730 2139.040 ;
        RECT 525.850 17.920 526.170 17.980 ;
        RECT 530.910 17.920 531.230 17.980 ;
        RECT 525.850 17.780 531.230 17.920 ;
        RECT 525.850 17.720 526.170 17.780 ;
        RECT 530.910 17.720 531.230 17.780 ;
      LAYER via ;
        RECT 530.940 2138.980 531.200 2139.240 ;
        RECT 1393.440 2138.980 1393.700 2139.240 ;
        RECT 525.880 17.720 526.140 17.980 ;
        RECT 530.940 17.720 531.200 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2139.435 1393.710 2139.805 ;
        RECT 1393.500 2139.270 1393.640 2139.435 ;
        RECT 530.940 2138.950 531.200 2139.270 ;
        RECT 1393.440 2138.950 1393.700 2139.270 ;
        RECT 531.000 18.010 531.140 2138.950 ;
        RECT 525.880 17.690 526.140 18.010 ;
        RECT 530.940 17.690 531.200 18.010 ;
        RECT 525.940 2.400 526.080 17.690 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2139.480 1393.710 2139.760 ;
      LAYER met3 ;
        RECT 1393.405 2139.770 1393.735 2139.785 ;
        RECT 1393.405 2139.720 1400.700 2139.770 ;
        RECT 1393.405 2139.470 1404.000 2139.720 ;
        RECT 1393.405 2139.455 1393.735 2139.470 ;
        RECT 1400.000 2139.120 1404.000 2139.470 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 544.710 2166.720 545.030 2166.780 ;
        RECT 1393.410 2166.720 1393.730 2166.780 ;
        RECT 544.710 2166.580 1393.730 2166.720 ;
        RECT 544.710 2166.520 545.030 2166.580 ;
        RECT 1393.410 2166.520 1393.730 2166.580 ;
      LAYER via ;
        RECT 544.740 2166.520 545.000 2166.780 ;
        RECT 1393.440 2166.520 1393.700 2166.780 ;
      LAYER met2 ;
        RECT 1393.430 2171.395 1393.710 2171.765 ;
        RECT 1393.500 2166.810 1393.640 2171.395 ;
        RECT 544.740 2166.490 545.000 2166.810 ;
        RECT 1393.440 2166.490 1393.700 2166.810 ;
        RECT 544.800 17.410 544.940 2166.490 ;
        RECT 543.880 17.270 544.940 17.410 ;
        RECT 543.880 2.400 544.020 17.270 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2171.440 1393.710 2171.720 ;
      LAYER met3 ;
        RECT 1393.405 2171.730 1393.735 2171.745 ;
        RECT 1393.405 2171.680 1400.700 2171.730 ;
        RECT 1393.405 2171.430 1404.000 2171.680 ;
        RECT 1393.405 2171.415 1393.735 2171.430 ;
        RECT 1400.000 2171.080 1404.000 2171.430 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 2201.400 565.730 2201.460 ;
        RECT 1393.410 2201.400 1393.730 2201.460 ;
        RECT 565.410 2201.260 1393.730 2201.400 ;
        RECT 565.410 2201.200 565.730 2201.260 ;
        RECT 1393.410 2201.200 1393.730 2201.260 ;
        RECT 561.730 17.920 562.050 17.980 ;
        RECT 565.410 17.920 565.730 17.980 ;
        RECT 561.730 17.780 565.730 17.920 ;
        RECT 561.730 17.720 562.050 17.780 ;
        RECT 565.410 17.720 565.730 17.780 ;
      LAYER via ;
        RECT 565.440 2201.200 565.700 2201.460 ;
        RECT 1393.440 2201.200 1393.700 2201.460 ;
        RECT 561.760 17.720 562.020 17.980 ;
        RECT 565.440 17.720 565.700 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2203.355 1393.710 2203.725 ;
        RECT 1393.500 2201.490 1393.640 2203.355 ;
        RECT 565.440 2201.170 565.700 2201.490 ;
        RECT 1393.440 2201.170 1393.700 2201.490 ;
        RECT 565.500 18.010 565.640 2201.170 ;
        RECT 561.760 17.690 562.020 18.010 ;
        RECT 565.440 17.690 565.700 18.010 ;
        RECT 561.820 2.400 561.960 17.690 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2203.400 1393.710 2203.680 ;
      LAYER met3 ;
        RECT 1393.405 2203.690 1393.735 2203.705 ;
        RECT 1393.405 2203.640 1400.700 2203.690 ;
        RECT 1393.405 2203.390 1404.000 2203.640 ;
        RECT 1393.405 2203.375 1393.735 2203.390 ;
        RECT 1400.000 2203.040 1404.000 2203.390 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 2228.940 585.970 2229.000 ;
        RECT 1393.410 2228.940 1393.730 2229.000 ;
        RECT 585.650 2228.800 1393.730 2228.940 ;
        RECT 585.650 2228.740 585.970 2228.800 ;
        RECT 1393.410 2228.740 1393.730 2228.800 ;
        RECT 579.670 17.920 579.990 17.980 ;
        RECT 585.650 17.920 585.970 17.980 ;
        RECT 579.670 17.780 585.970 17.920 ;
        RECT 579.670 17.720 579.990 17.780 ;
        RECT 585.650 17.720 585.970 17.780 ;
      LAYER via ;
        RECT 585.680 2228.740 585.940 2229.000 ;
        RECT 1393.440 2228.740 1393.700 2229.000 ;
        RECT 579.700 17.720 579.960 17.980 ;
        RECT 585.680 17.720 585.940 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2235.315 1393.710 2235.685 ;
        RECT 1393.500 2229.030 1393.640 2235.315 ;
        RECT 585.680 2228.710 585.940 2229.030 ;
        RECT 1393.440 2228.710 1393.700 2229.030 ;
        RECT 585.740 18.010 585.880 2228.710 ;
        RECT 579.700 17.690 579.960 18.010 ;
        RECT 585.680 17.690 585.940 18.010 ;
        RECT 579.760 2.400 579.900 17.690 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2235.360 1393.710 2235.640 ;
      LAYER met3 ;
        RECT 1393.405 2235.650 1393.735 2235.665 ;
        RECT 1393.405 2235.600 1400.700 2235.650 ;
        RECT 1393.405 2235.350 1404.000 2235.600 ;
        RECT 1393.405 2235.335 1393.735 2235.350 ;
        RECT 1400.000 2235.000 1404.000 2235.350 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 89.310 1352.760 89.630 1352.820 ;
        RECT 1393.410 1352.760 1393.730 1352.820 ;
        RECT 89.310 1352.620 1393.730 1352.760 ;
        RECT 89.310 1352.560 89.630 1352.620 ;
        RECT 1393.410 1352.560 1393.730 1352.620 ;
        RECT 86.090 17.920 86.410 17.980 ;
        RECT 89.310 17.920 89.630 17.980 ;
        RECT 86.090 17.780 89.630 17.920 ;
        RECT 86.090 17.720 86.410 17.780 ;
        RECT 89.310 17.720 89.630 17.780 ;
      LAYER via ;
        RECT 89.340 1352.560 89.600 1352.820 ;
        RECT 1393.440 1352.560 1393.700 1352.820 ;
        RECT 86.120 17.720 86.380 17.980 ;
        RECT 89.340 17.720 89.600 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1353.355 1393.710 1353.725 ;
        RECT 1393.500 1352.850 1393.640 1353.355 ;
        RECT 89.340 1352.530 89.600 1352.850 ;
        RECT 1393.440 1352.530 1393.700 1352.850 ;
        RECT 89.400 18.010 89.540 1352.530 ;
        RECT 86.120 17.690 86.380 18.010 ;
        RECT 89.340 17.690 89.600 18.010 ;
        RECT 86.180 2.400 86.320 17.690 ;
        RECT 85.970 -4.800 86.530 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1353.400 1393.710 1353.680 ;
      LAYER met3 ;
        RECT 1393.405 1353.690 1393.735 1353.705 ;
        RECT 1393.405 1353.640 1400.700 1353.690 ;
        RECT 1393.405 1353.390 1404.000 1353.640 ;
        RECT 1393.405 1353.375 1393.735 1353.390 ;
        RECT 1400.000 1353.040 1404.000 1353.390 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 2263.280 600.230 2263.340 ;
        RECT 1393.410 2263.280 1393.730 2263.340 ;
        RECT 599.910 2263.140 1393.730 2263.280 ;
        RECT 599.910 2263.080 600.230 2263.140 ;
        RECT 1393.410 2263.080 1393.730 2263.140 ;
        RECT 597.150 17.920 597.470 17.980 ;
        RECT 599.910 17.920 600.230 17.980 ;
        RECT 597.150 17.780 600.230 17.920 ;
        RECT 597.150 17.720 597.470 17.780 ;
        RECT 599.910 17.720 600.230 17.780 ;
      LAYER via ;
        RECT 599.940 2263.080 600.200 2263.340 ;
        RECT 1393.440 2263.080 1393.700 2263.340 ;
        RECT 597.180 17.720 597.440 17.980 ;
        RECT 599.940 17.720 600.200 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2266.595 1393.710 2266.965 ;
        RECT 1393.500 2263.370 1393.640 2266.595 ;
        RECT 599.940 2263.050 600.200 2263.370 ;
        RECT 1393.440 2263.050 1393.700 2263.370 ;
        RECT 600.000 18.010 600.140 2263.050 ;
        RECT 597.180 17.690 597.440 18.010 ;
        RECT 599.940 17.690 600.200 18.010 ;
        RECT 597.240 2.400 597.380 17.690 ;
        RECT 597.030 -4.800 597.590 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2266.640 1393.710 2266.920 ;
      LAYER met3 ;
        RECT 1393.405 2266.930 1393.735 2266.945 ;
        RECT 1393.405 2266.880 1400.700 2266.930 ;
        RECT 1393.405 2266.630 1404.000 2266.880 ;
        RECT 1393.405 2266.615 1393.735 2266.630 ;
        RECT 1400.000 2266.280 1404.000 2266.630 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 2297.960 620.930 2298.020 ;
        RECT 1393.410 2297.960 1393.730 2298.020 ;
        RECT 620.610 2297.820 1393.730 2297.960 ;
        RECT 620.610 2297.760 620.930 2297.820 ;
        RECT 1393.410 2297.760 1393.730 2297.820 ;
        RECT 615.090 17.920 615.410 17.980 ;
        RECT 620.610 17.920 620.930 17.980 ;
        RECT 615.090 17.780 620.930 17.920 ;
        RECT 615.090 17.720 615.410 17.780 ;
        RECT 620.610 17.720 620.930 17.780 ;
      LAYER via ;
        RECT 620.640 2297.760 620.900 2298.020 ;
        RECT 1393.440 2297.760 1393.700 2298.020 ;
        RECT 615.120 17.720 615.380 17.980 ;
        RECT 620.640 17.720 620.900 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2298.555 1393.710 2298.925 ;
        RECT 1393.500 2298.050 1393.640 2298.555 ;
        RECT 620.640 2297.730 620.900 2298.050 ;
        RECT 1393.440 2297.730 1393.700 2298.050 ;
        RECT 620.700 18.010 620.840 2297.730 ;
        RECT 615.120 17.690 615.380 18.010 ;
        RECT 620.640 17.690 620.900 18.010 ;
        RECT 615.180 2.400 615.320 17.690 ;
        RECT 614.970 -4.800 615.530 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2298.600 1393.710 2298.880 ;
      LAYER met3 ;
        RECT 1393.405 2298.890 1393.735 2298.905 ;
        RECT 1393.405 2298.840 1400.700 2298.890 ;
        RECT 1393.405 2298.590 1404.000 2298.840 ;
        RECT 1393.405 2298.575 1393.735 2298.590 ;
        RECT 1400.000 2298.240 1404.000 2298.590 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 1393.900 110.330 1393.960 ;
        RECT 1393.410 1393.900 1393.730 1393.960 ;
        RECT 110.010 1393.760 1393.730 1393.900 ;
        RECT 110.010 1393.700 110.330 1393.760 ;
        RECT 1393.410 1393.700 1393.730 1393.760 ;
      LAYER via ;
        RECT 110.040 1393.700 110.300 1393.960 ;
        RECT 1393.440 1393.700 1393.700 1393.960 ;
      LAYER met2 ;
        RECT 1393.430 1396.195 1393.710 1396.565 ;
        RECT 1393.500 1393.990 1393.640 1396.195 ;
        RECT 110.040 1393.670 110.300 1393.990 ;
        RECT 1393.440 1393.670 1393.700 1393.990 ;
        RECT 110.100 17.410 110.240 1393.670 ;
        RECT 109.640 17.270 110.240 17.410 ;
        RECT 109.640 2.400 109.780 17.270 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1396.240 1393.710 1396.520 ;
      LAYER met3 ;
        RECT 1393.405 1396.530 1393.735 1396.545 ;
        RECT 1393.405 1396.480 1400.700 1396.530 ;
        RECT 1393.405 1396.230 1404.000 1396.480 ;
        RECT 1393.405 1396.215 1393.735 1396.230 ;
        RECT 1400.000 1395.880 1404.000 1396.230 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 137.610 1435.380 137.930 1435.440 ;
        RECT 1393.410 1435.380 1393.730 1435.440 ;
        RECT 137.610 1435.240 1393.730 1435.380 ;
        RECT 137.610 1435.180 137.930 1435.240 ;
        RECT 1393.410 1435.180 1393.730 1435.240 ;
        RECT 133.470 17.920 133.790 17.980 ;
        RECT 137.610 17.920 137.930 17.980 ;
        RECT 133.470 17.780 137.930 17.920 ;
        RECT 133.470 17.720 133.790 17.780 ;
        RECT 137.610 17.720 137.930 17.780 ;
      LAYER via ;
        RECT 137.640 1435.180 137.900 1435.440 ;
        RECT 1393.440 1435.180 1393.700 1435.440 ;
        RECT 133.500 17.720 133.760 17.980 ;
        RECT 137.640 17.720 137.900 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1438.355 1393.710 1438.725 ;
        RECT 1393.500 1435.470 1393.640 1438.355 ;
        RECT 137.640 1435.150 137.900 1435.470 ;
        RECT 1393.440 1435.150 1393.700 1435.470 ;
        RECT 137.700 18.010 137.840 1435.150 ;
        RECT 133.500 17.690 133.760 18.010 ;
        RECT 137.640 17.690 137.900 18.010 ;
        RECT 133.560 2.400 133.700 17.690 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1438.400 1393.710 1438.680 ;
      LAYER met3 ;
        RECT 1393.405 1438.690 1393.735 1438.705 ;
        RECT 1393.405 1438.640 1400.700 1438.690 ;
        RECT 1393.405 1438.390 1404.000 1438.640 ;
        RECT 1393.405 1438.375 1393.735 1438.390 ;
        RECT 1400.000 1438.040 1404.000 1438.390 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 1470.060 151.730 1470.120 ;
        RECT 1393.410 1470.060 1393.730 1470.120 ;
        RECT 151.410 1469.920 1393.730 1470.060 ;
        RECT 151.410 1469.860 151.730 1469.920 ;
        RECT 1393.410 1469.860 1393.730 1469.920 ;
      LAYER via ;
        RECT 151.440 1469.860 151.700 1470.120 ;
        RECT 1393.440 1469.860 1393.700 1470.120 ;
      LAYER met2 ;
        RECT 1393.430 1470.315 1393.710 1470.685 ;
        RECT 1393.500 1470.150 1393.640 1470.315 ;
        RECT 151.440 1469.830 151.700 1470.150 ;
        RECT 1393.440 1469.830 1393.700 1470.150 ;
        RECT 151.500 2.400 151.640 1469.830 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1470.360 1393.710 1470.640 ;
      LAYER met3 ;
        RECT 1393.405 1470.650 1393.735 1470.665 ;
        RECT 1393.405 1470.600 1400.700 1470.650 ;
        RECT 1393.405 1470.350 1404.000 1470.600 ;
        RECT 1393.405 1470.335 1393.735 1470.350 ;
        RECT 1400.000 1470.000 1404.000 1470.350 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 172.110 1497.600 172.430 1497.660 ;
        RECT 1393.410 1497.600 1393.730 1497.660 ;
        RECT 172.110 1497.460 1393.730 1497.600 ;
        RECT 172.110 1497.400 172.430 1497.460 ;
        RECT 1393.410 1497.400 1393.730 1497.460 ;
        RECT 169.350 17.920 169.670 17.980 ;
        RECT 172.110 17.920 172.430 17.980 ;
        RECT 169.350 17.780 172.430 17.920 ;
        RECT 169.350 17.720 169.670 17.780 ;
        RECT 172.110 17.720 172.430 17.780 ;
      LAYER via ;
        RECT 172.140 1497.400 172.400 1497.660 ;
        RECT 1393.440 1497.400 1393.700 1497.660 ;
        RECT 169.380 17.720 169.640 17.980 ;
        RECT 172.140 17.720 172.400 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1502.275 1393.710 1502.645 ;
        RECT 1393.500 1497.690 1393.640 1502.275 ;
        RECT 172.140 1497.370 172.400 1497.690 ;
        RECT 1393.440 1497.370 1393.700 1497.690 ;
        RECT 172.200 18.010 172.340 1497.370 ;
        RECT 169.380 17.690 169.640 18.010 ;
        RECT 172.140 17.690 172.400 18.010 ;
        RECT 169.440 2.400 169.580 17.690 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1502.320 1393.710 1502.600 ;
      LAYER met3 ;
        RECT 1393.405 1502.610 1393.735 1502.625 ;
        RECT 1393.405 1502.560 1400.700 1502.610 ;
        RECT 1393.405 1502.310 1404.000 1502.560 ;
        RECT 1393.405 1502.295 1393.735 1502.310 ;
        RECT 1400.000 1501.960 1404.000 1502.310 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.350 1531.940 192.670 1532.000 ;
        RECT 1393.410 1531.940 1393.730 1532.000 ;
        RECT 192.350 1531.800 1393.730 1531.940 ;
        RECT 192.350 1531.740 192.670 1531.800 ;
        RECT 1393.410 1531.740 1393.730 1531.800 ;
        RECT 186.830 17.920 187.150 17.980 ;
        RECT 192.350 17.920 192.670 17.980 ;
        RECT 186.830 17.780 192.670 17.920 ;
        RECT 186.830 17.720 187.150 17.780 ;
        RECT 192.350 17.720 192.670 17.780 ;
      LAYER via ;
        RECT 192.380 1531.740 192.640 1532.000 ;
        RECT 1393.440 1531.740 1393.700 1532.000 ;
        RECT 186.860 17.720 187.120 17.980 ;
        RECT 192.380 17.720 192.640 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1534.235 1393.710 1534.605 ;
        RECT 1393.500 1532.030 1393.640 1534.235 ;
        RECT 192.380 1531.710 192.640 1532.030 ;
        RECT 1393.440 1531.710 1393.700 1532.030 ;
        RECT 192.440 18.010 192.580 1531.710 ;
        RECT 186.860 17.690 187.120 18.010 ;
        RECT 192.380 17.690 192.640 18.010 ;
        RECT 186.920 2.400 187.060 17.690 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1534.280 1393.710 1534.560 ;
      LAYER met3 ;
        RECT 1393.405 1534.570 1393.735 1534.585 ;
        RECT 1393.405 1534.520 1400.700 1534.570 ;
        RECT 1393.405 1534.270 1404.000 1534.520 ;
        RECT 1393.405 1534.255 1393.735 1534.270 ;
        RECT 1400.000 1533.920 1404.000 1534.270 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 206.610 1566.620 206.930 1566.680 ;
        RECT 1393.410 1566.620 1393.730 1566.680 ;
        RECT 206.610 1566.480 1393.730 1566.620 ;
        RECT 206.610 1566.420 206.930 1566.480 ;
        RECT 1393.410 1566.420 1393.730 1566.480 ;
      LAYER via ;
        RECT 206.640 1566.420 206.900 1566.680 ;
        RECT 1393.440 1566.420 1393.700 1566.680 ;
      LAYER met2 ;
        RECT 206.640 1566.390 206.900 1566.710 ;
        RECT 1393.440 1566.565 1393.700 1566.710 ;
        RECT 206.700 17.410 206.840 1566.390 ;
        RECT 1393.430 1566.195 1393.710 1566.565 ;
        RECT 204.860 17.270 206.840 17.410 ;
        RECT 204.860 2.400 205.000 17.270 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1566.240 1393.710 1566.520 ;
      LAYER met3 ;
        RECT 1393.405 1566.530 1393.735 1566.545 ;
        RECT 1393.405 1566.480 1400.700 1566.530 ;
        RECT 1393.405 1566.230 1404.000 1566.480 ;
        RECT 1393.405 1566.215 1393.735 1566.230 ;
        RECT 1400.000 1565.880 1404.000 1566.230 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 227.310 1594.160 227.630 1594.220 ;
        RECT 1393.410 1594.160 1393.730 1594.220 ;
        RECT 227.310 1594.020 1393.730 1594.160 ;
        RECT 227.310 1593.960 227.630 1594.020 ;
        RECT 1393.410 1593.960 1393.730 1594.020 ;
        RECT 222.710 17.920 223.030 17.980 ;
        RECT 227.310 17.920 227.630 17.980 ;
        RECT 222.710 17.780 227.630 17.920 ;
        RECT 222.710 17.720 223.030 17.780 ;
        RECT 227.310 17.720 227.630 17.780 ;
      LAYER via ;
        RECT 227.340 1593.960 227.600 1594.220 ;
        RECT 1393.440 1593.960 1393.700 1594.220 ;
        RECT 222.740 17.720 223.000 17.980 ;
        RECT 227.340 17.720 227.600 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1597.475 1393.710 1597.845 ;
        RECT 1393.500 1594.250 1393.640 1597.475 ;
        RECT 227.340 1593.930 227.600 1594.250 ;
        RECT 1393.440 1593.930 1393.700 1594.250 ;
        RECT 227.400 18.010 227.540 1593.930 ;
        RECT 222.740 17.690 223.000 18.010 ;
        RECT 227.340 17.690 227.600 18.010 ;
        RECT 222.800 2.400 222.940 17.690 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1597.520 1393.710 1597.800 ;
      LAYER met3 ;
        RECT 1393.405 1597.810 1393.735 1597.825 ;
        RECT 1393.405 1597.760 1400.700 1597.810 ;
        RECT 1393.405 1597.510 1404.000 1597.760 ;
        RECT 1393.405 1597.495 1393.735 1597.510 ;
        RECT 1400.000 1597.160 1404.000 1597.510 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 17.240 20.630 17.300 ;
        RECT 1390.190 17.240 1390.510 17.300 ;
        RECT 20.310 17.100 1390.510 17.240 ;
        RECT 20.310 17.040 20.630 17.100 ;
        RECT 1390.190 17.040 1390.510 17.100 ;
      LAYER via ;
        RECT 20.340 17.040 20.600 17.300 ;
        RECT 1390.220 17.040 1390.480 17.300 ;
      LAYER met2 ;
        RECT 1390.210 1236.395 1390.490 1236.765 ;
        RECT 1390.280 17.330 1390.420 1236.395 ;
        RECT 20.340 17.010 20.600 17.330 ;
        RECT 1390.220 17.010 1390.480 17.330 ;
        RECT 20.400 2.400 20.540 17.010 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 1390.210 1236.440 1390.490 1236.720 ;
      LAYER met3 ;
        RECT 1390.185 1236.730 1390.515 1236.745 ;
        RECT 1390.185 1236.680 1400.700 1236.730 ;
        RECT 1390.185 1236.430 1404.000 1236.680 ;
        RECT 1390.185 1236.415 1390.515 1236.430 ;
        RECT 1400.000 1236.080 1404.000 1236.430 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 1276.600 48.230 1276.660 ;
        RECT 1393.410 1276.600 1393.730 1276.660 ;
        RECT 47.910 1276.460 1393.730 1276.600 ;
        RECT 47.910 1276.400 48.230 1276.460 ;
        RECT 1393.410 1276.400 1393.730 1276.460 ;
        RECT 44.230 17.920 44.550 17.980 ;
        RECT 47.910 17.920 48.230 17.980 ;
        RECT 44.230 17.780 48.230 17.920 ;
        RECT 44.230 17.720 44.550 17.780 ;
        RECT 47.910 17.720 48.230 17.780 ;
      LAYER via ;
        RECT 47.940 1276.400 48.200 1276.660 ;
        RECT 1393.440 1276.400 1393.700 1276.660 ;
        RECT 44.260 17.720 44.520 17.980 ;
        RECT 47.940 17.720 48.200 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1279.235 1393.710 1279.605 ;
        RECT 1393.500 1276.690 1393.640 1279.235 ;
        RECT 47.940 1276.370 48.200 1276.690 ;
        RECT 1393.440 1276.370 1393.700 1276.690 ;
        RECT 48.000 18.010 48.140 1276.370 ;
        RECT 44.260 17.690 44.520 18.010 ;
        RECT 47.940 17.690 48.200 18.010 ;
        RECT 44.320 2.400 44.460 17.690 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1279.280 1393.710 1279.560 ;
      LAYER met3 ;
        RECT 1393.405 1279.570 1393.735 1279.585 ;
        RECT 1393.405 1279.520 1400.700 1279.570 ;
        RECT 1393.405 1279.270 1404.000 1279.520 ;
        RECT 1393.405 1279.255 1393.735 1279.270 ;
        RECT 1400.000 1278.920 1404.000 1279.270 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 1635.640 248.330 1635.700 ;
        RECT 1393.410 1635.640 1393.730 1635.700 ;
        RECT 248.010 1635.500 1393.730 1635.640 ;
        RECT 248.010 1635.440 248.330 1635.500 ;
        RECT 1393.410 1635.440 1393.730 1635.500 ;
      LAYER via ;
        RECT 248.040 1635.440 248.300 1635.700 ;
        RECT 1393.440 1635.440 1393.700 1635.700 ;
      LAYER met2 ;
        RECT 1393.430 1640.315 1393.710 1640.685 ;
        RECT 1393.500 1635.730 1393.640 1640.315 ;
        RECT 248.040 1635.410 248.300 1635.730 ;
        RECT 1393.440 1635.410 1393.700 1635.730 ;
        RECT 248.100 17.410 248.240 1635.410 ;
        RECT 246.720 17.270 248.240 17.410 ;
        RECT 246.720 2.400 246.860 17.270 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1640.360 1393.710 1640.640 ;
      LAYER met3 ;
        RECT 1393.405 1640.650 1393.735 1640.665 ;
        RECT 1393.405 1640.600 1400.700 1640.650 ;
        RECT 1393.405 1640.350 1404.000 1640.600 ;
        RECT 1393.405 1640.335 1393.735 1640.350 ;
        RECT 1400.000 1640.000 1404.000 1640.350 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.710 1669.980 269.030 1670.040 ;
        RECT 1393.410 1669.980 1393.730 1670.040 ;
        RECT 268.710 1669.840 1393.730 1669.980 ;
        RECT 268.710 1669.780 269.030 1669.840 ;
        RECT 1393.410 1669.780 1393.730 1669.840 ;
        RECT 264.110 17.920 264.430 17.980 ;
        RECT 268.710 17.920 269.030 17.980 ;
        RECT 264.110 17.780 269.030 17.920 ;
        RECT 264.110 17.720 264.430 17.780 ;
        RECT 268.710 17.720 269.030 17.780 ;
      LAYER via ;
        RECT 268.740 1669.780 269.000 1670.040 ;
        RECT 1393.440 1669.780 1393.700 1670.040 ;
        RECT 264.140 17.720 264.400 17.980 ;
        RECT 268.740 17.720 269.000 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1672.275 1393.710 1672.645 ;
        RECT 1393.500 1670.070 1393.640 1672.275 ;
        RECT 268.740 1669.750 269.000 1670.070 ;
        RECT 1393.440 1669.750 1393.700 1670.070 ;
        RECT 268.800 18.010 268.940 1669.750 ;
        RECT 264.140 17.690 264.400 18.010 ;
        RECT 268.740 17.690 269.000 18.010 ;
        RECT 264.200 2.400 264.340 17.690 ;
        RECT 263.990 -4.800 264.550 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1672.320 1393.710 1672.600 ;
      LAYER met3 ;
        RECT 1393.405 1672.610 1393.735 1672.625 ;
        RECT 1393.405 1672.560 1400.700 1672.610 ;
        RECT 1393.405 1672.310 1404.000 1672.560 ;
        RECT 1393.405 1672.295 1393.735 1672.310 ;
        RECT 1400.000 1671.960 1404.000 1672.310 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.510 1704.660 282.830 1704.720 ;
        RECT 1393.410 1704.660 1393.730 1704.720 ;
        RECT 282.510 1704.520 1393.730 1704.660 ;
        RECT 282.510 1704.460 282.830 1704.520 ;
        RECT 1393.410 1704.460 1393.730 1704.520 ;
      LAYER via ;
        RECT 282.540 1704.460 282.800 1704.720 ;
        RECT 1393.440 1704.460 1393.700 1704.720 ;
      LAYER met2 ;
        RECT 282.540 1704.430 282.800 1704.750 ;
        RECT 1393.440 1704.605 1393.700 1704.750 ;
        RECT 282.600 17.410 282.740 1704.430 ;
        RECT 1393.430 1704.235 1393.710 1704.605 ;
        RECT 282.140 17.270 282.740 17.410 ;
        RECT 282.140 2.400 282.280 17.270 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1704.280 1393.710 1704.560 ;
      LAYER met3 ;
        RECT 1393.405 1704.570 1393.735 1704.585 ;
        RECT 1393.405 1704.520 1400.700 1704.570 ;
        RECT 1393.405 1704.270 1404.000 1704.520 ;
        RECT 1393.405 1704.255 1393.735 1704.270 ;
        RECT 1400.000 1703.920 1404.000 1704.270 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 303.210 1732.200 303.530 1732.260 ;
        RECT 1393.410 1732.200 1393.730 1732.260 ;
        RECT 303.210 1732.060 1393.730 1732.200 ;
        RECT 303.210 1732.000 303.530 1732.060 ;
        RECT 1393.410 1732.000 1393.730 1732.060 ;
        RECT 299.990 17.920 300.310 17.980 ;
        RECT 303.210 17.920 303.530 17.980 ;
        RECT 299.990 17.780 303.530 17.920 ;
        RECT 299.990 17.720 300.310 17.780 ;
        RECT 303.210 17.720 303.530 17.780 ;
      LAYER via ;
        RECT 303.240 1732.000 303.500 1732.260 ;
        RECT 1393.440 1732.000 1393.700 1732.260 ;
        RECT 300.020 17.720 300.280 17.980 ;
        RECT 303.240 17.720 303.500 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1735.515 1393.710 1735.885 ;
        RECT 1393.500 1732.290 1393.640 1735.515 ;
        RECT 303.240 1731.970 303.500 1732.290 ;
        RECT 1393.440 1731.970 1393.700 1732.290 ;
        RECT 303.300 18.010 303.440 1731.970 ;
        RECT 300.020 17.690 300.280 18.010 ;
        RECT 303.240 17.690 303.500 18.010 ;
        RECT 300.080 2.400 300.220 17.690 ;
        RECT 299.870 -4.800 300.430 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1735.560 1393.710 1735.840 ;
      LAYER met3 ;
        RECT 1393.405 1735.850 1393.735 1735.865 ;
        RECT 1393.405 1735.800 1400.700 1735.850 ;
        RECT 1393.405 1735.550 1404.000 1735.800 ;
        RECT 1393.405 1735.535 1393.735 1735.550 ;
        RECT 1400.000 1735.200 1404.000 1735.550 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.450 1766.540 323.770 1766.600 ;
        RECT 1390.190 1766.540 1390.510 1766.600 ;
        RECT 323.450 1766.400 1390.510 1766.540 ;
        RECT 323.450 1766.340 323.770 1766.400 ;
        RECT 1390.190 1766.340 1390.510 1766.400 ;
        RECT 317.930 17.920 318.250 17.980 ;
        RECT 323.450 17.920 323.770 17.980 ;
        RECT 317.930 17.780 323.770 17.920 ;
        RECT 317.930 17.720 318.250 17.780 ;
        RECT 323.450 17.720 323.770 17.780 ;
      LAYER via ;
        RECT 323.480 1766.340 323.740 1766.600 ;
        RECT 1390.220 1766.340 1390.480 1766.600 ;
        RECT 317.960 17.720 318.220 17.980 ;
        RECT 323.480 17.720 323.740 17.980 ;
      LAYER met2 ;
        RECT 1390.210 1767.475 1390.490 1767.845 ;
        RECT 1390.280 1766.630 1390.420 1767.475 ;
        RECT 323.480 1766.310 323.740 1766.630 ;
        RECT 1390.220 1766.310 1390.480 1766.630 ;
        RECT 323.540 18.010 323.680 1766.310 ;
        RECT 317.960 17.690 318.220 18.010 ;
        RECT 323.480 17.690 323.740 18.010 ;
        RECT 318.020 2.400 318.160 17.690 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 1390.210 1767.520 1390.490 1767.800 ;
      LAYER met3 ;
        RECT 1390.185 1767.810 1390.515 1767.825 ;
        RECT 1390.185 1767.760 1400.700 1767.810 ;
        RECT 1390.185 1767.510 1404.000 1767.760 ;
        RECT 1390.185 1767.495 1390.515 1767.510 ;
        RECT 1400.000 1767.160 1404.000 1767.510 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 337.710 1794.080 338.030 1794.140 ;
        RECT 1389.270 1794.080 1389.590 1794.140 ;
        RECT 337.710 1793.940 1389.590 1794.080 ;
        RECT 337.710 1793.880 338.030 1793.940 ;
        RECT 1389.270 1793.880 1389.590 1793.940 ;
      LAYER via ;
        RECT 337.740 1793.880 338.000 1794.140 ;
        RECT 1389.300 1793.880 1389.560 1794.140 ;
      LAYER met2 ;
        RECT 1389.290 1799.435 1389.570 1799.805 ;
        RECT 1389.360 1794.170 1389.500 1799.435 ;
        RECT 337.740 1793.850 338.000 1794.170 ;
        RECT 1389.300 1793.850 1389.560 1794.170 ;
        RECT 337.800 17.410 337.940 1793.850 ;
        RECT 335.960 17.270 337.940 17.410 ;
        RECT 335.960 2.400 336.100 17.270 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 1389.290 1799.480 1389.570 1799.760 ;
      LAYER met3 ;
        RECT 1389.265 1799.770 1389.595 1799.785 ;
        RECT 1389.265 1799.720 1400.700 1799.770 ;
        RECT 1389.265 1799.470 1404.000 1799.720 ;
        RECT 1389.265 1799.455 1389.595 1799.470 ;
        RECT 1400.000 1799.120 1404.000 1799.470 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 358.410 1828.760 358.730 1828.820 ;
        RECT 1393.410 1828.760 1393.730 1828.820 ;
        RECT 358.410 1828.620 1393.730 1828.760 ;
        RECT 358.410 1828.560 358.730 1828.620 ;
        RECT 1393.410 1828.560 1393.730 1828.620 ;
        RECT 353.350 17.920 353.670 17.980 ;
        RECT 358.410 17.920 358.730 17.980 ;
        RECT 353.350 17.780 358.730 17.920 ;
        RECT 353.350 17.720 353.670 17.780 ;
        RECT 358.410 17.720 358.730 17.780 ;
      LAYER via ;
        RECT 358.440 1828.560 358.700 1828.820 ;
        RECT 1393.440 1828.560 1393.700 1828.820 ;
        RECT 353.380 17.720 353.640 17.980 ;
        RECT 358.440 17.720 358.700 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1831.395 1393.710 1831.765 ;
        RECT 1393.500 1828.850 1393.640 1831.395 ;
        RECT 358.440 1828.530 358.700 1828.850 ;
        RECT 1393.440 1828.530 1393.700 1828.850 ;
        RECT 358.500 18.010 358.640 1828.530 ;
        RECT 353.380 17.690 353.640 18.010 ;
        RECT 358.440 17.690 358.700 18.010 ;
        RECT 353.440 2.400 353.580 17.690 ;
        RECT 353.230 -4.800 353.790 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1831.440 1393.710 1831.720 ;
      LAYER met3 ;
        RECT 1393.405 1831.730 1393.735 1831.745 ;
        RECT 1393.405 1831.680 1400.700 1831.730 ;
        RECT 1393.405 1831.430 1404.000 1831.680 ;
        RECT 1393.405 1831.415 1393.735 1831.430 ;
        RECT 1400.000 1831.080 1404.000 1831.430 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 1863.100 372.530 1863.160 ;
        RECT 1390.190 1863.100 1390.510 1863.160 ;
        RECT 372.210 1862.960 1390.510 1863.100 ;
        RECT 372.210 1862.900 372.530 1862.960 ;
        RECT 1390.190 1862.900 1390.510 1862.960 ;
      LAYER via ;
        RECT 372.240 1862.900 372.500 1863.160 ;
        RECT 1390.220 1862.900 1390.480 1863.160 ;
      LAYER met2 ;
        RECT 1390.210 1863.355 1390.490 1863.725 ;
        RECT 1390.280 1863.190 1390.420 1863.355 ;
        RECT 372.240 1862.870 372.500 1863.190 ;
        RECT 1390.220 1862.870 1390.480 1863.190 ;
        RECT 372.300 17.410 372.440 1862.870 ;
        RECT 371.380 17.270 372.440 17.410 ;
        RECT 371.380 2.400 371.520 17.270 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 1390.210 1863.400 1390.490 1863.680 ;
      LAYER met3 ;
        RECT 1390.185 1863.690 1390.515 1863.705 ;
        RECT 1390.185 1863.640 1400.700 1863.690 ;
        RECT 1390.185 1863.390 1404.000 1863.640 ;
        RECT 1390.185 1863.375 1390.515 1863.390 ;
        RECT 1400.000 1863.040 1404.000 1863.390 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 1890.980 393.230 1891.040 ;
        RECT 1393.410 1890.980 1393.730 1891.040 ;
        RECT 392.910 1890.840 1393.730 1890.980 ;
        RECT 392.910 1890.780 393.230 1890.840 ;
        RECT 1393.410 1890.780 1393.730 1890.840 ;
        RECT 389.230 17.920 389.550 17.980 ;
        RECT 392.910 17.920 393.230 17.980 ;
        RECT 389.230 17.780 393.230 17.920 ;
        RECT 389.230 17.720 389.550 17.780 ;
        RECT 392.910 17.720 393.230 17.780 ;
      LAYER via ;
        RECT 392.940 1890.780 393.200 1891.040 ;
        RECT 1393.440 1890.780 1393.700 1891.040 ;
        RECT 389.260 17.720 389.520 17.980 ;
        RECT 392.940 17.720 393.200 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1895.315 1393.710 1895.685 ;
        RECT 1393.500 1891.070 1393.640 1895.315 ;
        RECT 392.940 1890.750 393.200 1891.070 ;
        RECT 1393.440 1890.750 1393.700 1891.070 ;
        RECT 393.000 18.010 393.140 1890.750 ;
        RECT 389.260 17.690 389.520 18.010 ;
        RECT 392.940 17.690 393.200 18.010 ;
        RECT 389.320 2.400 389.460 17.690 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1895.360 1393.710 1895.640 ;
      LAYER met3 ;
        RECT 1393.405 1895.650 1393.735 1895.665 ;
        RECT 1393.405 1895.600 1400.700 1895.650 ;
        RECT 1393.405 1895.350 1404.000 1895.600 ;
        RECT 1393.405 1895.335 1393.735 1895.350 ;
        RECT 1400.000 1895.000 1404.000 1895.350 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.150 1925.320 413.470 1925.380 ;
        RECT 1388.350 1925.320 1388.670 1925.380 ;
        RECT 413.150 1925.180 1388.670 1925.320 ;
        RECT 413.150 1925.120 413.470 1925.180 ;
        RECT 1388.350 1925.120 1388.670 1925.180 ;
        RECT 407.170 17.920 407.490 17.980 ;
        RECT 413.150 17.920 413.470 17.980 ;
        RECT 407.170 17.780 413.470 17.920 ;
        RECT 407.170 17.720 407.490 17.780 ;
        RECT 413.150 17.720 413.470 17.780 ;
      LAYER via ;
        RECT 413.180 1925.120 413.440 1925.380 ;
        RECT 1388.380 1925.120 1388.640 1925.380 ;
        RECT 407.200 17.720 407.460 17.980 ;
        RECT 413.180 17.720 413.440 17.980 ;
      LAYER met2 ;
        RECT 1388.370 1927.275 1388.650 1927.645 ;
        RECT 1388.440 1925.410 1388.580 1927.275 ;
        RECT 413.180 1925.090 413.440 1925.410 ;
        RECT 1388.380 1925.090 1388.640 1925.410 ;
        RECT 413.240 18.010 413.380 1925.090 ;
        RECT 407.200 17.690 407.460 18.010 ;
        RECT 413.180 17.690 413.440 18.010 ;
        RECT 407.260 2.400 407.400 17.690 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 1388.370 1927.320 1388.650 1927.600 ;
      LAYER met3 ;
        RECT 1388.345 1927.610 1388.675 1927.625 ;
        RECT 1388.345 1927.560 1400.700 1927.610 ;
        RECT 1388.345 1927.310 1404.000 1927.560 ;
        RECT 1388.345 1927.295 1388.675 1927.310 ;
        RECT 1400.000 1926.960 1404.000 1927.310 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.610 1318.080 68.930 1318.140 ;
        RECT 1393.410 1318.080 1393.730 1318.140 ;
        RECT 68.610 1317.940 1393.730 1318.080 ;
        RECT 68.610 1317.880 68.930 1317.940 ;
        RECT 1393.410 1317.880 1393.730 1317.940 ;
      LAYER via ;
        RECT 68.640 1317.880 68.900 1318.140 ;
        RECT 1393.440 1317.880 1393.700 1318.140 ;
      LAYER met2 ;
        RECT 1393.430 1321.395 1393.710 1321.765 ;
        RECT 1393.500 1318.170 1393.640 1321.395 ;
        RECT 68.640 1317.850 68.900 1318.170 ;
        RECT 1393.440 1317.850 1393.700 1318.170 ;
        RECT 68.700 17.410 68.840 1317.850 ;
        RECT 68.240 17.270 68.840 17.410 ;
        RECT 68.240 2.400 68.380 17.270 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1321.440 1393.710 1321.720 ;
      LAYER met3 ;
        RECT 1393.405 1321.730 1393.735 1321.745 ;
        RECT 1393.405 1321.680 1400.700 1321.730 ;
        RECT 1393.405 1321.430 1404.000 1321.680 ;
        RECT 1393.405 1321.415 1393.735 1321.430 ;
        RECT 1400.000 1321.080 1404.000 1321.430 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 1952.860 427.730 1952.920 ;
        RECT 1391.570 1952.860 1391.890 1952.920 ;
        RECT 427.410 1952.720 1391.890 1952.860 ;
        RECT 427.410 1952.660 427.730 1952.720 ;
        RECT 1391.570 1952.660 1391.890 1952.720 ;
        RECT 424.650 17.920 424.970 17.980 ;
        RECT 427.410 17.920 427.730 17.980 ;
        RECT 424.650 17.780 427.730 17.920 ;
        RECT 424.650 17.720 424.970 17.780 ;
        RECT 427.410 17.720 427.730 17.780 ;
      LAYER via ;
        RECT 427.440 1952.660 427.700 1952.920 ;
        RECT 1391.600 1952.660 1391.860 1952.920 ;
        RECT 424.680 17.720 424.940 17.980 ;
        RECT 427.440 17.720 427.700 17.980 ;
      LAYER met2 ;
        RECT 1391.590 1958.555 1391.870 1958.925 ;
        RECT 1391.660 1952.950 1391.800 1958.555 ;
        RECT 427.440 1952.630 427.700 1952.950 ;
        RECT 1391.600 1952.630 1391.860 1952.950 ;
        RECT 427.500 18.010 427.640 1952.630 ;
        RECT 424.680 17.690 424.940 18.010 ;
        RECT 427.440 17.690 427.700 18.010 ;
        RECT 424.740 2.400 424.880 17.690 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 1391.590 1958.600 1391.870 1958.880 ;
      LAYER met3 ;
        RECT 1391.565 1958.890 1391.895 1958.905 ;
        RECT 1391.565 1958.840 1400.700 1958.890 ;
        RECT 1391.565 1958.590 1404.000 1958.840 ;
        RECT 1391.565 1958.575 1391.895 1958.590 ;
        RECT 1400.000 1958.240 1404.000 1958.590 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 1987.540 448.430 1987.600 ;
        RECT 1393.410 1987.540 1393.730 1987.600 ;
        RECT 448.110 1987.400 1393.730 1987.540 ;
        RECT 448.110 1987.340 448.430 1987.400 ;
        RECT 1393.410 1987.340 1393.730 1987.400 ;
        RECT 442.590 17.920 442.910 17.980 ;
        RECT 448.110 17.920 448.430 17.980 ;
        RECT 442.590 17.780 448.430 17.920 ;
        RECT 442.590 17.720 442.910 17.780 ;
        RECT 448.110 17.720 448.430 17.780 ;
      LAYER via ;
        RECT 448.140 1987.340 448.400 1987.600 ;
        RECT 1393.440 1987.340 1393.700 1987.600 ;
        RECT 442.620 17.720 442.880 17.980 ;
        RECT 448.140 17.720 448.400 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1990.515 1393.710 1990.885 ;
        RECT 1393.500 1987.630 1393.640 1990.515 ;
        RECT 448.140 1987.310 448.400 1987.630 ;
        RECT 1393.440 1987.310 1393.700 1987.630 ;
        RECT 448.200 18.010 448.340 1987.310 ;
        RECT 442.620 17.690 442.880 18.010 ;
        RECT 448.140 17.690 448.400 18.010 ;
        RECT 442.680 2.400 442.820 17.690 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1990.560 1393.710 1990.840 ;
      LAYER met3 ;
        RECT 1393.405 1990.850 1393.735 1990.865 ;
        RECT 1393.405 1990.800 1400.700 1990.850 ;
        RECT 1393.405 1990.550 1404.000 1990.800 ;
        RECT 1393.405 1990.535 1393.735 1990.550 ;
        RECT 1400.000 1990.200 1404.000 1990.550 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 2021.880 462.230 2021.940 ;
        RECT 1393.410 2021.880 1393.730 2021.940 ;
        RECT 461.910 2021.740 1393.730 2021.880 ;
        RECT 461.910 2021.680 462.230 2021.740 ;
        RECT 1393.410 2021.680 1393.730 2021.740 ;
      LAYER via ;
        RECT 461.940 2021.680 462.200 2021.940 ;
        RECT 1393.440 2021.680 1393.700 2021.940 ;
      LAYER met2 ;
        RECT 1393.430 2022.475 1393.710 2022.845 ;
        RECT 1393.500 2021.970 1393.640 2022.475 ;
        RECT 461.940 2021.650 462.200 2021.970 ;
        RECT 1393.440 2021.650 1393.700 2021.970 ;
        RECT 462.000 17.410 462.140 2021.650 ;
        RECT 460.620 17.270 462.140 17.410 ;
        RECT 460.620 2.400 460.760 17.270 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2022.520 1393.710 2022.800 ;
      LAYER met3 ;
        RECT 1393.405 2022.810 1393.735 2022.825 ;
        RECT 1393.405 2022.760 1400.700 2022.810 ;
        RECT 1393.405 2022.510 1404.000 2022.760 ;
        RECT 1393.405 2022.495 1393.735 2022.510 ;
        RECT 1400.000 2022.160 1404.000 2022.510 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 2049.420 482.930 2049.480 ;
        RECT 1393.410 2049.420 1393.730 2049.480 ;
        RECT 482.610 2049.280 1393.730 2049.420 ;
        RECT 482.610 2049.220 482.930 2049.280 ;
        RECT 1393.410 2049.220 1393.730 2049.280 ;
        RECT 478.470 17.920 478.790 17.980 ;
        RECT 482.610 17.920 482.930 17.980 ;
        RECT 478.470 17.780 482.930 17.920 ;
        RECT 478.470 17.720 478.790 17.780 ;
        RECT 482.610 17.720 482.930 17.780 ;
      LAYER via ;
        RECT 482.640 2049.220 482.900 2049.480 ;
        RECT 1393.440 2049.220 1393.700 2049.480 ;
        RECT 478.500 17.720 478.760 17.980 ;
        RECT 482.640 17.720 482.900 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2054.435 1393.710 2054.805 ;
        RECT 1393.500 2049.510 1393.640 2054.435 ;
        RECT 482.640 2049.190 482.900 2049.510 ;
        RECT 1393.440 2049.190 1393.700 2049.510 ;
        RECT 482.700 18.010 482.840 2049.190 ;
        RECT 478.500 17.690 478.760 18.010 ;
        RECT 482.640 17.690 482.900 18.010 ;
        RECT 478.560 2.400 478.700 17.690 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2054.480 1393.710 2054.760 ;
      LAYER met3 ;
        RECT 1393.405 2054.770 1393.735 2054.785 ;
        RECT 1393.405 2054.720 1400.700 2054.770 ;
        RECT 1393.405 2054.470 1404.000 2054.720 ;
        RECT 1393.405 2054.455 1393.735 2054.470 ;
        RECT 1400.000 2054.120 1404.000 2054.470 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 2084.100 496.730 2084.160 ;
        RECT 1393.410 2084.100 1393.730 2084.160 ;
        RECT 496.410 2083.960 1393.730 2084.100 ;
        RECT 496.410 2083.900 496.730 2083.960 ;
        RECT 1393.410 2083.900 1393.730 2083.960 ;
      LAYER via ;
        RECT 496.440 2083.900 496.700 2084.160 ;
        RECT 1393.440 2083.900 1393.700 2084.160 ;
      LAYER met2 ;
        RECT 1393.430 2086.395 1393.710 2086.765 ;
        RECT 1393.500 2084.190 1393.640 2086.395 ;
        RECT 496.440 2083.870 496.700 2084.190 ;
        RECT 1393.440 2083.870 1393.700 2084.190 ;
        RECT 496.500 2.400 496.640 2083.870 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2086.440 1393.710 2086.720 ;
      LAYER met3 ;
        RECT 1393.405 2086.730 1393.735 2086.745 ;
        RECT 1393.405 2086.680 1400.700 2086.730 ;
        RECT 1393.405 2086.430 1404.000 2086.680 ;
        RECT 1393.405 2086.415 1393.735 2086.430 ;
        RECT 1400.000 2086.080 1404.000 2086.430 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 2118.440 517.430 2118.500 ;
        RECT 1393.410 2118.440 1393.730 2118.500 ;
        RECT 517.110 2118.300 1393.730 2118.440 ;
        RECT 517.110 2118.240 517.430 2118.300 ;
        RECT 1393.410 2118.240 1393.730 2118.300 ;
        RECT 513.890 17.920 514.210 17.980 ;
        RECT 517.110 17.920 517.430 17.980 ;
        RECT 513.890 17.780 517.430 17.920 ;
        RECT 513.890 17.720 514.210 17.780 ;
        RECT 517.110 17.720 517.430 17.780 ;
      LAYER via ;
        RECT 517.140 2118.240 517.400 2118.500 ;
        RECT 1393.440 2118.240 1393.700 2118.500 ;
        RECT 513.920 17.720 514.180 17.980 ;
        RECT 517.140 17.720 517.400 17.980 ;
      LAYER met2 ;
        RECT 517.140 2118.210 517.400 2118.530 ;
        RECT 1393.430 2118.355 1393.710 2118.725 ;
        RECT 1393.440 2118.210 1393.700 2118.355 ;
        RECT 517.200 18.010 517.340 2118.210 ;
        RECT 513.920 17.690 514.180 18.010 ;
        RECT 517.140 17.690 517.400 18.010 ;
        RECT 513.980 2.400 514.120 17.690 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2118.400 1393.710 2118.680 ;
      LAYER met3 ;
        RECT 1393.405 2118.690 1393.735 2118.705 ;
        RECT 1393.405 2118.640 1400.700 2118.690 ;
        RECT 1393.405 2118.390 1404.000 2118.640 ;
        RECT 1393.405 2118.375 1393.735 2118.390 ;
        RECT 1400.000 2118.040 1404.000 2118.390 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.350 2145.980 537.670 2146.040 ;
        RECT 1388.350 2145.980 1388.670 2146.040 ;
        RECT 537.350 2145.840 1388.670 2145.980 ;
        RECT 537.350 2145.780 537.670 2145.840 ;
        RECT 1388.350 2145.780 1388.670 2145.840 ;
        RECT 531.830 17.920 532.150 17.980 ;
        RECT 537.350 17.920 537.670 17.980 ;
        RECT 531.830 17.780 537.670 17.920 ;
        RECT 531.830 17.720 532.150 17.780 ;
        RECT 537.350 17.720 537.670 17.780 ;
      LAYER via ;
        RECT 537.380 2145.780 537.640 2146.040 ;
        RECT 1388.380 2145.780 1388.640 2146.040 ;
        RECT 531.860 17.720 532.120 17.980 ;
        RECT 537.380 17.720 537.640 17.980 ;
      LAYER met2 ;
        RECT 1388.370 2150.315 1388.650 2150.685 ;
        RECT 1388.440 2146.070 1388.580 2150.315 ;
        RECT 537.380 2145.750 537.640 2146.070 ;
        RECT 1388.380 2145.750 1388.640 2146.070 ;
        RECT 537.440 18.010 537.580 2145.750 ;
        RECT 531.860 17.690 532.120 18.010 ;
        RECT 537.380 17.690 537.640 18.010 ;
        RECT 531.920 2.400 532.060 17.690 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 1388.370 2150.360 1388.650 2150.640 ;
      LAYER met3 ;
        RECT 1388.345 2150.650 1388.675 2150.665 ;
        RECT 1388.345 2150.600 1400.700 2150.650 ;
        RECT 1388.345 2150.350 1404.000 2150.600 ;
        RECT 1388.345 2150.335 1388.675 2150.350 ;
        RECT 1400.000 2150.000 1404.000 2150.350 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 2180.660 551.930 2180.720 ;
        RECT 1390.190 2180.660 1390.510 2180.720 ;
        RECT 551.610 2180.520 1390.510 2180.660 ;
        RECT 551.610 2180.460 551.930 2180.520 ;
        RECT 1390.190 2180.460 1390.510 2180.520 ;
      LAYER via ;
        RECT 551.640 2180.460 551.900 2180.720 ;
        RECT 1390.220 2180.460 1390.480 2180.720 ;
      LAYER met2 ;
        RECT 1390.210 2181.595 1390.490 2181.965 ;
        RECT 1390.280 2180.750 1390.420 2181.595 ;
        RECT 551.640 2180.430 551.900 2180.750 ;
        RECT 1390.220 2180.430 1390.480 2180.750 ;
        RECT 551.700 17.410 551.840 2180.430 ;
        RECT 549.860 17.270 551.840 17.410 ;
        RECT 549.860 2.400 550.000 17.270 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 1390.210 2181.640 1390.490 2181.920 ;
      LAYER met3 ;
        RECT 1390.185 2181.930 1390.515 2181.945 ;
        RECT 1390.185 2181.880 1400.700 2181.930 ;
        RECT 1390.185 2181.630 1404.000 2181.880 ;
        RECT 1390.185 2181.615 1390.515 2181.630 ;
        RECT 1400.000 2181.280 1404.000 2181.630 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 2208.200 572.630 2208.260 ;
        RECT 1389.270 2208.200 1389.590 2208.260 ;
        RECT 572.310 2208.060 1389.590 2208.200 ;
        RECT 572.310 2208.000 572.630 2208.060 ;
        RECT 1389.270 2208.000 1389.590 2208.060 ;
        RECT 567.710 17.920 568.030 17.980 ;
        RECT 572.310 17.920 572.630 17.980 ;
        RECT 567.710 17.780 572.630 17.920 ;
        RECT 567.710 17.720 568.030 17.780 ;
        RECT 572.310 17.720 572.630 17.780 ;
      LAYER via ;
        RECT 572.340 2208.000 572.600 2208.260 ;
        RECT 1389.300 2208.000 1389.560 2208.260 ;
        RECT 567.740 17.720 568.000 17.980 ;
        RECT 572.340 17.720 572.600 17.980 ;
      LAYER met2 ;
        RECT 1389.290 2213.555 1389.570 2213.925 ;
        RECT 1389.360 2208.290 1389.500 2213.555 ;
        RECT 572.340 2207.970 572.600 2208.290 ;
        RECT 1389.300 2207.970 1389.560 2208.290 ;
        RECT 572.400 18.010 572.540 2207.970 ;
        RECT 567.740 17.690 568.000 18.010 ;
        RECT 572.340 17.690 572.600 18.010 ;
        RECT 567.800 2.400 567.940 17.690 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1389.290 2213.600 1389.570 2213.880 ;
      LAYER met3 ;
        RECT 1389.265 2213.890 1389.595 2213.905 ;
        RECT 1389.265 2213.840 1400.700 2213.890 ;
        RECT 1389.265 2213.590 1404.000 2213.840 ;
        RECT 1389.265 2213.575 1389.595 2213.590 ;
        RECT 1400.000 2213.240 1404.000 2213.590 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 586.110 2242.880 586.430 2242.940 ;
        RECT 1393.410 2242.880 1393.730 2242.940 ;
        RECT 586.110 2242.740 1393.730 2242.880 ;
        RECT 586.110 2242.680 586.430 2242.740 ;
        RECT 1393.410 2242.680 1393.730 2242.740 ;
      LAYER via ;
        RECT 586.140 2242.680 586.400 2242.940 ;
        RECT 1393.440 2242.680 1393.700 2242.940 ;
      LAYER met2 ;
        RECT 1393.430 2245.515 1393.710 2245.885 ;
        RECT 1393.500 2242.970 1393.640 2245.515 ;
        RECT 586.140 2242.650 586.400 2242.970 ;
        RECT 1393.440 2242.650 1393.700 2242.970 ;
        RECT 586.200 17.410 586.340 2242.650 ;
        RECT 585.740 17.270 586.340 17.410 ;
        RECT 585.740 2.400 585.880 17.270 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2245.560 1393.710 2245.840 ;
      LAYER met3 ;
        RECT 1393.405 2245.850 1393.735 2245.865 ;
        RECT 1393.405 2245.800 1400.700 2245.850 ;
        RECT 1393.405 2245.550 1404.000 2245.800 ;
        RECT 1393.405 2245.535 1393.735 2245.550 ;
        RECT 1400.000 2245.200 1404.000 2245.550 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 96.210 1359.560 96.530 1359.620 ;
        RECT 1393.410 1359.560 1393.730 1359.620 ;
        RECT 96.210 1359.420 1393.730 1359.560 ;
        RECT 96.210 1359.360 96.530 1359.420 ;
        RECT 1393.410 1359.360 1393.730 1359.420 ;
        RECT 91.610 17.920 91.930 17.980 ;
        RECT 96.210 17.920 96.530 17.980 ;
        RECT 91.610 17.780 96.530 17.920 ;
        RECT 91.610 17.720 91.930 17.780 ;
        RECT 96.210 17.720 96.530 17.780 ;
      LAYER via ;
        RECT 96.240 1359.360 96.500 1359.620 ;
        RECT 1393.440 1359.360 1393.700 1359.620 ;
        RECT 91.640 17.720 91.900 17.980 ;
        RECT 96.240 17.720 96.500 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1364.235 1393.710 1364.605 ;
        RECT 1393.500 1359.650 1393.640 1364.235 ;
        RECT 96.240 1359.330 96.500 1359.650 ;
        RECT 1393.440 1359.330 1393.700 1359.650 ;
        RECT 96.300 18.010 96.440 1359.330 ;
        RECT 91.640 17.690 91.900 18.010 ;
        RECT 96.240 17.690 96.500 18.010 ;
        RECT 91.700 2.400 91.840 17.690 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1364.280 1393.710 1364.560 ;
      LAYER met3 ;
        RECT 1393.405 1364.570 1393.735 1364.585 ;
        RECT 1393.405 1364.520 1400.700 1364.570 ;
        RECT 1393.405 1364.270 1404.000 1364.520 ;
        RECT 1393.405 1364.255 1393.735 1364.270 ;
        RECT 1400.000 1363.920 1404.000 1364.270 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 2277.220 607.130 2277.280 ;
        RECT 1393.410 2277.220 1393.730 2277.280 ;
        RECT 606.810 2277.080 1393.730 2277.220 ;
        RECT 606.810 2277.020 607.130 2277.080 ;
        RECT 1393.410 2277.020 1393.730 2277.080 ;
        RECT 603.130 17.920 603.450 17.980 ;
        RECT 606.810 17.920 607.130 17.980 ;
        RECT 603.130 17.780 607.130 17.920 ;
        RECT 603.130 17.720 603.450 17.780 ;
        RECT 606.810 17.720 607.130 17.780 ;
      LAYER via ;
        RECT 606.840 2277.020 607.100 2277.280 ;
        RECT 1393.440 2277.020 1393.700 2277.280 ;
        RECT 603.160 17.720 603.420 17.980 ;
        RECT 606.840 17.720 607.100 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2277.475 1393.710 2277.845 ;
        RECT 1393.500 2277.310 1393.640 2277.475 ;
        RECT 606.840 2276.990 607.100 2277.310 ;
        RECT 1393.440 2276.990 1393.700 2277.310 ;
        RECT 606.900 18.010 607.040 2276.990 ;
        RECT 603.160 17.690 603.420 18.010 ;
        RECT 606.840 17.690 607.100 18.010 ;
        RECT 603.220 2.400 603.360 17.690 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2277.520 1393.710 2277.800 ;
      LAYER met3 ;
        RECT 1393.405 2277.810 1393.735 2277.825 ;
        RECT 1393.405 2277.760 1400.700 2277.810 ;
        RECT 1393.405 2277.510 1404.000 2277.760 ;
        RECT 1393.405 2277.495 1393.735 2277.510 ;
        RECT 1400.000 2277.160 1404.000 2277.510 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.050 2304.760 627.370 2304.820 ;
        RECT 1393.410 2304.760 1393.730 2304.820 ;
        RECT 627.050 2304.620 1393.730 2304.760 ;
        RECT 627.050 2304.560 627.370 2304.620 ;
        RECT 1393.410 2304.560 1393.730 2304.620 ;
        RECT 621.070 17.920 621.390 17.980 ;
        RECT 627.050 17.920 627.370 17.980 ;
        RECT 621.070 17.780 627.370 17.920 ;
        RECT 621.070 17.720 621.390 17.780 ;
        RECT 627.050 17.720 627.370 17.780 ;
      LAYER via ;
        RECT 627.080 2304.560 627.340 2304.820 ;
        RECT 1393.440 2304.560 1393.700 2304.820 ;
        RECT 621.100 17.720 621.360 17.980 ;
        RECT 627.080 17.720 627.340 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2309.435 1393.710 2309.805 ;
        RECT 1393.500 2304.850 1393.640 2309.435 ;
        RECT 627.080 2304.530 627.340 2304.850 ;
        RECT 1393.440 2304.530 1393.700 2304.850 ;
        RECT 627.140 18.010 627.280 2304.530 ;
        RECT 621.100 17.690 621.360 18.010 ;
        RECT 627.080 17.690 627.340 18.010 ;
        RECT 621.160 2.400 621.300 17.690 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2309.480 1393.710 2309.760 ;
      LAYER met3 ;
        RECT 1393.405 2309.770 1393.735 2309.785 ;
        RECT 1393.405 2309.720 1400.700 2309.770 ;
        RECT 1393.405 2309.470 1404.000 2309.720 ;
        RECT 1393.405 2309.455 1393.735 2309.470 ;
        RECT 1400.000 2309.120 1404.000 2309.470 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 1401.040 117.230 1401.100 ;
        RECT 1389.270 1401.040 1389.590 1401.100 ;
        RECT 116.910 1400.900 1389.590 1401.040 ;
        RECT 116.910 1400.840 117.230 1400.900 ;
        RECT 1389.270 1400.840 1389.590 1400.900 ;
      LAYER via ;
        RECT 116.940 1400.840 117.200 1401.100 ;
        RECT 1389.300 1400.840 1389.560 1401.100 ;
      LAYER met2 ;
        RECT 1389.290 1406.395 1389.570 1406.765 ;
        RECT 1389.360 1401.130 1389.500 1406.395 ;
        RECT 116.940 1400.810 117.200 1401.130 ;
        RECT 1389.300 1400.810 1389.560 1401.130 ;
        RECT 117.000 17.410 117.140 1400.810 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 1389.290 1406.440 1389.570 1406.720 ;
      LAYER met3 ;
        RECT 1389.265 1406.730 1389.595 1406.745 ;
        RECT 1389.265 1406.680 1400.700 1406.730 ;
        RECT 1389.265 1406.430 1404.000 1406.680 ;
        RECT 1389.265 1406.415 1389.595 1406.430 ;
        RECT 1400.000 1406.080 1404.000 1406.430 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 144.510 1449.320 144.830 1449.380 ;
        RECT 1393.410 1449.320 1393.730 1449.380 ;
        RECT 144.510 1449.180 1393.730 1449.320 ;
        RECT 144.510 1449.120 144.830 1449.180 ;
        RECT 1393.410 1449.120 1393.730 1449.180 ;
        RECT 139.450 17.920 139.770 17.980 ;
        RECT 144.510 17.920 144.830 17.980 ;
        RECT 139.450 17.780 144.830 17.920 ;
        RECT 139.450 17.720 139.770 17.780 ;
        RECT 144.510 17.720 144.830 17.780 ;
      LAYER via ;
        RECT 144.540 1449.120 144.800 1449.380 ;
        RECT 1393.440 1449.120 1393.700 1449.380 ;
        RECT 139.480 17.720 139.740 17.980 ;
        RECT 144.540 17.720 144.800 17.980 ;
      LAYER met2 ;
        RECT 144.540 1449.090 144.800 1449.410 ;
        RECT 1393.430 1449.235 1393.710 1449.605 ;
        RECT 1393.440 1449.090 1393.700 1449.235 ;
        RECT 144.600 18.010 144.740 1449.090 ;
        RECT 139.480 17.690 139.740 18.010 ;
        RECT 144.540 17.690 144.800 18.010 ;
        RECT 139.540 2.400 139.680 17.690 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1449.280 1393.710 1449.560 ;
      LAYER met3 ;
        RECT 1393.405 1449.570 1393.735 1449.585 ;
        RECT 1393.405 1449.520 1400.700 1449.570 ;
        RECT 1393.405 1449.270 1404.000 1449.520 ;
        RECT 1393.405 1449.255 1393.735 1449.270 ;
        RECT 1400.000 1448.920 1404.000 1449.270 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 1476.860 158.630 1476.920 ;
        RECT 1393.410 1476.860 1393.730 1476.920 ;
        RECT 158.310 1476.720 1393.730 1476.860 ;
        RECT 158.310 1476.660 158.630 1476.720 ;
        RECT 1393.410 1476.660 1393.730 1476.720 ;
      LAYER via ;
        RECT 158.340 1476.660 158.600 1476.920 ;
        RECT 1393.440 1476.660 1393.700 1476.920 ;
      LAYER met2 ;
        RECT 1393.430 1481.195 1393.710 1481.565 ;
        RECT 1393.500 1476.950 1393.640 1481.195 ;
        RECT 158.340 1476.630 158.600 1476.950 ;
        RECT 1393.440 1476.630 1393.700 1476.950 ;
        RECT 158.400 17.410 158.540 1476.630 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1481.240 1393.710 1481.520 ;
      LAYER met3 ;
        RECT 1393.405 1481.530 1393.735 1481.545 ;
        RECT 1393.405 1481.480 1400.700 1481.530 ;
        RECT 1393.405 1481.230 1404.000 1481.480 ;
        RECT 1393.405 1481.215 1393.735 1481.230 ;
        RECT 1400.000 1480.880 1404.000 1481.230 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 179.010 1511.200 179.330 1511.260 ;
        RECT 1393.410 1511.200 1393.730 1511.260 ;
        RECT 179.010 1511.060 1393.730 1511.200 ;
        RECT 179.010 1511.000 179.330 1511.060 ;
        RECT 1393.410 1511.000 1393.730 1511.060 ;
        RECT 174.870 17.920 175.190 17.980 ;
        RECT 179.010 17.920 179.330 17.980 ;
        RECT 174.870 17.780 179.330 17.920 ;
        RECT 174.870 17.720 175.190 17.780 ;
        RECT 179.010 17.720 179.330 17.780 ;
      LAYER via ;
        RECT 179.040 1511.000 179.300 1511.260 ;
        RECT 1393.440 1511.000 1393.700 1511.260 ;
        RECT 174.900 17.720 175.160 17.980 ;
        RECT 179.040 17.720 179.300 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1512.475 1393.710 1512.845 ;
        RECT 1393.500 1511.290 1393.640 1512.475 ;
        RECT 179.040 1510.970 179.300 1511.290 ;
        RECT 1393.440 1510.970 1393.700 1511.290 ;
        RECT 179.100 18.010 179.240 1510.970 ;
        RECT 174.900 17.690 175.160 18.010 ;
        RECT 179.040 17.690 179.300 18.010 ;
        RECT 174.960 2.400 175.100 17.690 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1512.520 1393.710 1512.800 ;
      LAYER met3 ;
        RECT 1393.405 1512.810 1393.735 1512.825 ;
        RECT 1393.405 1512.760 1400.700 1512.810 ;
        RECT 1393.405 1512.510 1404.000 1512.760 ;
        RECT 1393.405 1512.495 1393.735 1512.510 ;
        RECT 1400.000 1512.160 1404.000 1512.510 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 1539.080 193.130 1539.140 ;
        RECT 1389.270 1539.080 1389.590 1539.140 ;
        RECT 192.810 1538.940 1389.590 1539.080 ;
        RECT 192.810 1538.880 193.130 1538.940 ;
        RECT 1389.270 1538.880 1389.590 1538.940 ;
      LAYER via ;
        RECT 192.840 1538.880 193.100 1539.140 ;
        RECT 1389.300 1538.880 1389.560 1539.140 ;
      LAYER met2 ;
        RECT 1389.290 1544.435 1389.570 1544.805 ;
        RECT 1389.360 1539.170 1389.500 1544.435 ;
        RECT 192.840 1538.850 193.100 1539.170 ;
        RECT 1389.300 1538.850 1389.560 1539.170 ;
        RECT 192.900 2.400 193.040 1538.850 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 1389.290 1544.480 1389.570 1544.760 ;
      LAYER met3 ;
        RECT 1389.265 1544.770 1389.595 1544.785 ;
        RECT 1389.265 1544.720 1400.700 1544.770 ;
        RECT 1389.265 1544.470 1404.000 1544.720 ;
        RECT 1389.265 1544.455 1389.595 1544.470 ;
        RECT 1400.000 1544.120 1404.000 1544.470 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 1573.420 213.830 1573.480 ;
        RECT 1393.410 1573.420 1393.730 1573.480 ;
        RECT 213.510 1573.280 1393.730 1573.420 ;
        RECT 213.510 1573.220 213.830 1573.280 ;
        RECT 1393.410 1573.220 1393.730 1573.280 ;
        RECT 210.750 17.920 211.070 17.980 ;
        RECT 213.510 17.920 213.830 17.980 ;
        RECT 210.750 17.780 213.830 17.920 ;
        RECT 210.750 17.720 211.070 17.780 ;
        RECT 213.510 17.720 213.830 17.780 ;
      LAYER via ;
        RECT 213.540 1573.220 213.800 1573.480 ;
        RECT 1393.440 1573.220 1393.700 1573.480 ;
        RECT 210.780 17.720 211.040 17.980 ;
        RECT 213.540 17.720 213.800 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1576.395 1393.710 1576.765 ;
        RECT 1393.500 1573.510 1393.640 1576.395 ;
        RECT 213.540 1573.190 213.800 1573.510 ;
        RECT 1393.440 1573.190 1393.700 1573.510 ;
        RECT 213.600 18.010 213.740 1573.190 ;
        RECT 210.780 17.690 211.040 18.010 ;
        RECT 213.540 17.690 213.800 18.010 ;
        RECT 210.840 2.400 210.980 17.690 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1576.440 1393.710 1576.720 ;
      LAYER met3 ;
        RECT 1393.405 1576.730 1393.735 1576.745 ;
        RECT 1393.405 1576.680 1400.700 1576.730 ;
        RECT 1393.405 1576.430 1404.000 1576.680 ;
        RECT 1393.405 1576.415 1393.735 1576.430 ;
        RECT 1400.000 1576.080 1404.000 1576.430 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 234.210 1608.100 234.530 1608.160 ;
        RECT 1390.190 1608.100 1390.510 1608.160 ;
        RECT 234.210 1607.960 1390.510 1608.100 ;
        RECT 234.210 1607.900 234.530 1607.960 ;
        RECT 1390.190 1607.900 1390.510 1607.960 ;
        RECT 228.690 17.920 229.010 17.980 ;
        RECT 234.210 17.920 234.530 17.980 ;
        RECT 228.690 17.780 234.530 17.920 ;
        RECT 228.690 17.720 229.010 17.780 ;
        RECT 234.210 17.720 234.530 17.780 ;
      LAYER via ;
        RECT 234.240 1607.900 234.500 1608.160 ;
        RECT 1390.220 1607.900 1390.480 1608.160 ;
        RECT 228.720 17.720 228.980 17.980 ;
        RECT 234.240 17.720 234.500 17.980 ;
      LAYER met2 ;
        RECT 1390.210 1608.355 1390.490 1608.725 ;
        RECT 1390.280 1608.190 1390.420 1608.355 ;
        RECT 234.240 1607.870 234.500 1608.190 ;
        RECT 1390.220 1607.870 1390.480 1608.190 ;
        RECT 234.300 18.010 234.440 1607.870 ;
        RECT 228.720 17.690 228.980 18.010 ;
        RECT 234.240 17.690 234.500 18.010 ;
        RECT 228.780 2.400 228.920 17.690 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 1390.210 1608.400 1390.490 1608.680 ;
      LAYER met3 ;
        RECT 1390.185 1608.690 1390.515 1608.705 ;
        RECT 1390.185 1608.640 1400.700 1608.690 ;
        RECT 1390.185 1608.390 1404.000 1608.640 ;
        RECT 1390.185 1608.375 1390.515 1608.390 ;
        RECT 1400.000 1608.040 1404.000 1608.390 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 54.810 1283.740 55.130 1283.800 ;
        RECT 1389.270 1283.740 1389.590 1283.800 ;
        RECT 54.810 1283.600 1389.590 1283.740 ;
        RECT 54.810 1283.540 55.130 1283.600 ;
        RECT 1389.270 1283.540 1389.590 1283.600 ;
        RECT 50.210 17.920 50.530 17.980 ;
        RECT 54.810 17.920 55.130 17.980 ;
        RECT 50.210 17.780 55.130 17.920 ;
        RECT 50.210 17.720 50.530 17.780 ;
        RECT 54.810 17.720 55.130 17.780 ;
      LAYER via ;
        RECT 54.840 1283.540 55.100 1283.800 ;
        RECT 1389.300 1283.540 1389.560 1283.800 ;
        RECT 50.240 17.720 50.500 17.980 ;
        RECT 54.840 17.720 55.100 17.980 ;
      LAYER met2 ;
        RECT 1389.290 1289.435 1389.570 1289.805 ;
        RECT 1389.360 1283.830 1389.500 1289.435 ;
        RECT 54.840 1283.510 55.100 1283.830 ;
        RECT 1389.300 1283.510 1389.560 1283.830 ;
        RECT 54.900 18.010 55.040 1283.510 ;
        RECT 50.240 17.690 50.500 18.010 ;
        RECT 54.840 17.690 55.100 18.010 ;
        RECT 50.300 2.400 50.440 17.690 ;
        RECT 50.090 -4.800 50.650 2.400 ;
      LAYER via2 ;
        RECT 1389.290 1289.480 1389.570 1289.760 ;
      LAYER met3 ;
        RECT 1389.265 1289.770 1389.595 1289.785 ;
        RECT 1389.265 1289.720 1400.700 1289.770 ;
        RECT 1389.265 1289.470 1404.000 1289.720 ;
        RECT 1389.265 1289.455 1389.595 1289.470 ;
        RECT 1400.000 1289.120 1404.000 1289.470 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 1649.240 255.230 1649.300 ;
        RECT 1393.410 1649.240 1393.730 1649.300 ;
        RECT 254.910 1649.100 1393.730 1649.240 ;
        RECT 254.910 1649.040 255.230 1649.100 ;
        RECT 1393.410 1649.040 1393.730 1649.100 ;
        RECT 252.610 17.920 252.930 17.980 ;
        RECT 254.910 17.920 255.230 17.980 ;
        RECT 252.610 17.780 255.230 17.920 ;
        RECT 252.610 17.720 252.930 17.780 ;
        RECT 254.910 17.720 255.230 17.780 ;
      LAYER via ;
        RECT 254.940 1649.040 255.200 1649.300 ;
        RECT 1393.440 1649.040 1393.700 1649.300 ;
        RECT 252.640 17.720 252.900 17.980 ;
        RECT 254.940 17.720 255.200 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1651.195 1393.710 1651.565 ;
        RECT 1393.500 1649.330 1393.640 1651.195 ;
        RECT 254.940 1649.010 255.200 1649.330 ;
        RECT 1393.440 1649.010 1393.700 1649.330 ;
        RECT 255.000 18.010 255.140 1649.010 ;
        RECT 252.640 17.690 252.900 18.010 ;
        RECT 254.940 17.690 255.200 18.010 ;
        RECT 252.700 2.400 252.840 17.690 ;
        RECT 252.490 -4.800 253.050 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1651.240 1393.710 1651.520 ;
      LAYER met3 ;
        RECT 1393.405 1651.530 1393.735 1651.545 ;
        RECT 1393.405 1651.480 1400.700 1651.530 ;
        RECT 1393.405 1651.230 1404.000 1651.480 ;
        RECT 1393.405 1651.215 1393.735 1651.230 ;
        RECT 1400.000 1650.880 1404.000 1651.230 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 275.610 1676.780 275.930 1676.840 ;
        RECT 1389.270 1676.780 1389.590 1676.840 ;
        RECT 275.610 1676.640 1389.590 1676.780 ;
        RECT 275.610 1676.580 275.930 1676.640 ;
        RECT 1389.270 1676.580 1389.590 1676.640 ;
        RECT 270.090 17.920 270.410 17.980 ;
        RECT 275.610 17.920 275.930 17.980 ;
        RECT 270.090 17.780 275.930 17.920 ;
        RECT 270.090 17.720 270.410 17.780 ;
        RECT 275.610 17.720 275.930 17.780 ;
      LAYER via ;
        RECT 275.640 1676.580 275.900 1676.840 ;
        RECT 1389.300 1676.580 1389.560 1676.840 ;
        RECT 270.120 17.720 270.380 17.980 ;
        RECT 275.640 17.720 275.900 17.980 ;
      LAYER met2 ;
        RECT 1389.290 1682.475 1389.570 1682.845 ;
        RECT 1389.360 1676.870 1389.500 1682.475 ;
        RECT 275.640 1676.550 275.900 1676.870 ;
        RECT 1389.300 1676.550 1389.560 1676.870 ;
        RECT 275.700 18.010 275.840 1676.550 ;
        RECT 270.120 17.690 270.380 18.010 ;
        RECT 275.640 17.690 275.900 18.010 ;
        RECT 270.180 2.400 270.320 17.690 ;
        RECT 269.970 -4.800 270.530 2.400 ;
      LAYER via2 ;
        RECT 1389.290 1682.520 1389.570 1682.800 ;
      LAYER met3 ;
        RECT 1389.265 1682.810 1389.595 1682.825 ;
        RECT 1389.265 1682.760 1400.700 1682.810 ;
        RECT 1389.265 1682.510 1404.000 1682.760 ;
        RECT 1389.265 1682.495 1389.595 1682.510 ;
        RECT 1400.000 1682.160 1404.000 1682.510 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 1711.460 289.730 1711.520 ;
        RECT 1391.570 1711.460 1391.890 1711.520 ;
        RECT 289.410 1711.320 1391.890 1711.460 ;
        RECT 289.410 1711.260 289.730 1711.320 ;
        RECT 1391.570 1711.260 1391.890 1711.320 ;
      LAYER via ;
        RECT 289.440 1711.260 289.700 1711.520 ;
        RECT 1391.600 1711.260 1391.860 1711.520 ;
      LAYER met2 ;
        RECT 1391.590 1714.435 1391.870 1714.805 ;
        RECT 1391.660 1711.550 1391.800 1714.435 ;
        RECT 289.440 1711.230 289.700 1711.550 ;
        RECT 1391.600 1711.230 1391.860 1711.550 ;
        RECT 289.500 17.410 289.640 1711.230 ;
        RECT 288.120 17.270 289.640 17.410 ;
        RECT 288.120 2.400 288.260 17.270 ;
        RECT 287.910 -4.800 288.470 2.400 ;
      LAYER via2 ;
        RECT 1391.590 1714.480 1391.870 1714.760 ;
      LAYER met3 ;
        RECT 1391.565 1714.770 1391.895 1714.785 ;
        RECT 1391.565 1714.720 1400.700 1714.770 ;
        RECT 1391.565 1714.470 1404.000 1714.720 ;
        RECT 1391.565 1714.455 1391.895 1714.470 ;
        RECT 1400.000 1714.120 1404.000 1714.470 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 310.110 1745.800 310.430 1745.860 ;
        RECT 1393.410 1745.800 1393.730 1745.860 ;
        RECT 310.110 1745.660 1393.730 1745.800 ;
        RECT 310.110 1745.600 310.430 1745.660 ;
        RECT 1393.410 1745.600 1393.730 1745.660 ;
        RECT 305.970 17.920 306.290 17.980 ;
        RECT 310.110 17.920 310.430 17.980 ;
        RECT 305.970 17.780 310.430 17.920 ;
        RECT 305.970 17.720 306.290 17.780 ;
        RECT 310.110 17.720 310.430 17.780 ;
      LAYER via ;
        RECT 310.140 1745.600 310.400 1745.860 ;
        RECT 1393.440 1745.600 1393.700 1745.860 ;
        RECT 306.000 17.720 306.260 17.980 ;
        RECT 310.140 17.720 310.400 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1746.395 1393.710 1746.765 ;
        RECT 1393.500 1745.890 1393.640 1746.395 ;
        RECT 310.140 1745.570 310.400 1745.890 ;
        RECT 1393.440 1745.570 1393.700 1745.890 ;
        RECT 310.200 18.010 310.340 1745.570 ;
        RECT 306.000 17.690 306.260 18.010 ;
        RECT 310.140 17.690 310.400 18.010 ;
        RECT 306.060 2.400 306.200 17.690 ;
        RECT 305.850 -4.800 306.410 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1746.440 1393.710 1746.720 ;
      LAYER met3 ;
        RECT 1393.405 1746.730 1393.735 1746.745 ;
        RECT 1393.405 1746.680 1400.700 1746.730 ;
        RECT 1393.405 1746.430 1404.000 1746.680 ;
        RECT 1393.405 1746.415 1393.735 1746.430 ;
        RECT 1400.000 1746.080 1404.000 1746.430 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 1773.680 324.230 1773.740 ;
        RECT 1393.410 1773.680 1393.730 1773.740 ;
        RECT 323.910 1773.540 1393.730 1773.680 ;
        RECT 323.910 1773.480 324.230 1773.540 ;
        RECT 1393.410 1773.480 1393.730 1773.540 ;
      LAYER via ;
        RECT 323.940 1773.480 324.200 1773.740 ;
        RECT 1393.440 1773.480 1393.700 1773.740 ;
      LAYER met2 ;
        RECT 1393.430 1778.355 1393.710 1778.725 ;
        RECT 1393.500 1773.770 1393.640 1778.355 ;
        RECT 323.940 1773.450 324.200 1773.770 ;
        RECT 1393.440 1773.450 1393.700 1773.770 ;
        RECT 324.000 2.400 324.140 1773.450 ;
        RECT 323.790 -4.800 324.350 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1778.400 1393.710 1778.680 ;
      LAYER met3 ;
        RECT 1393.405 1778.690 1393.735 1778.705 ;
        RECT 1393.405 1778.640 1400.700 1778.690 ;
        RECT 1393.405 1778.390 1404.000 1778.640 ;
        RECT 1393.405 1778.375 1393.735 1778.390 ;
        RECT 1400.000 1778.040 1404.000 1778.390 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 344.610 1808.020 344.930 1808.080 ;
        RECT 1393.410 1808.020 1393.730 1808.080 ;
        RECT 344.610 1807.880 1393.730 1808.020 ;
        RECT 344.610 1807.820 344.930 1807.880 ;
        RECT 1393.410 1807.820 1393.730 1807.880 ;
        RECT 341.390 17.920 341.710 17.980 ;
        RECT 344.610 17.920 344.930 17.980 ;
        RECT 341.390 17.780 344.930 17.920 ;
        RECT 341.390 17.720 341.710 17.780 ;
        RECT 344.610 17.720 344.930 17.780 ;
      LAYER via ;
        RECT 344.640 1807.820 344.900 1808.080 ;
        RECT 1393.440 1807.820 1393.700 1808.080 ;
        RECT 341.420 17.720 341.680 17.980 ;
        RECT 344.640 17.720 344.900 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1810.315 1393.710 1810.685 ;
        RECT 1393.500 1808.110 1393.640 1810.315 ;
        RECT 344.640 1807.790 344.900 1808.110 ;
        RECT 1393.440 1807.790 1393.700 1808.110 ;
        RECT 344.700 18.010 344.840 1807.790 ;
        RECT 341.420 17.690 341.680 18.010 ;
        RECT 344.640 17.690 344.900 18.010 ;
        RECT 341.480 2.400 341.620 17.690 ;
        RECT 341.270 -4.800 341.830 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1810.360 1393.710 1810.640 ;
      LAYER met3 ;
        RECT 1393.405 1810.650 1393.735 1810.665 ;
        RECT 1393.405 1810.600 1400.700 1810.650 ;
        RECT 1393.405 1810.350 1404.000 1810.600 ;
        RECT 1393.405 1810.335 1393.735 1810.350 ;
        RECT 1400.000 1810.000 1404.000 1810.350 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 1842.700 365.170 1842.760 ;
        RECT 1393.410 1842.700 1393.730 1842.760 ;
        RECT 364.850 1842.560 1393.730 1842.700 ;
        RECT 364.850 1842.500 365.170 1842.560 ;
        RECT 1393.410 1842.500 1393.730 1842.560 ;
        RECT 359.330 17.920 359.650 17.980 ;
        RECT 364.850 17.920 365.170 17.980 ;
        RECT 359.330 17.780 365.170 17.920 ;
        RECT 359.330 17.720 359.650 17.780 ;
        RECT 364.850 17.720 365.170 17.780 ;
      LAYER via ;
        RECT 364.880 1842.500 365.140 1842.760 ;
        RECT 1393.440 1842.500 1393.700 1842.760 ;
        RECT 359.360 17.720 359.620 17.980 ;
        RECT 364.880 17.720 365.140 17.980 ;
      LAYER met2 ;
        RECT 364.880 1842.470 365.140 1842.790 ;
        RECT 1393.440 1842.645 1393.700 1842.790 ;
        RECT 364.940 18.010 365.080 1842.470 ;
        RECT 1393.430 1842.275 1393.710 1842.645 ;
        RECT 359.360 17.690 359.620 18.010 ;
        RECT 364.880 17.690 365.140 18.010 ;
        RECT 359.420 2.400 359.560 17.690 ;
        RECT 359.210 -4.800 359.770 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1842.320 1393.710 1842.600 ;
      LAYER met3 ;
        RECT 1393.405 1842.610 1393.735 1842.625 ;
        RECT 1393.405 1842.560 1400.700 1842.610 ;
        RECT 1393.405 1842.310 1404.000 1842.560 ;
        RECT 1393.405 1842.295 1393.735 1842.310 ;
        RECT 1400.000 1841.960 1404.000 1842.310 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 379.110 1870.240 379.430 1870.300 ;
        RECT 1392.030 1870.240 1392.350 1870.300 ;
        RECT 379.110 1870.100 1392.350 1870.240 ;
        RECT 379.110 1870.040 379.430 1870.100 ;
        RECT 1392.030 1870.040 1392.350 1870.100 ;
      LAYER via ;
        RECT 379.140 1870.040 379.400 1870.300 ;
        RECT 1392.060 1870.040 1392.320 1870.300 ;
      LAYER met2 ;
        RECT 1392.050 1874.235 1392.330 1874.605 ;
        RECT 1392.120 1870.330 1392.260 1874.235 ;
        RECT 379.140 1870.010 379.400 1870.330 ;
        RECT 1392.060 1870.010 1392.320 1870.330 ;
        RECT 379.200 17.410 379.340 1870.010 ;
        RECT 377.360 17.270 379.340 17.410 ;
        RECT 377.360 2.400 377.500 17.270 ;
        RECT 377.150 -4.800 377.710 2.400 ;
      LAYER via2 ;
        RECT 1392.050 1874.280 1392.330 1874.560 ;
      LAYER met3 ;
        RECT 1392.025 1874.570 1392.355 1874.585 ;
        RECT 1392.025 1874.520 1400.700 1874.570 ;
        RECT 1392.025 1874.270 1404.000 1874.520 ;
        RECT 1392.025 1874.255 1392.355 1874.270 ;
        RECT 1400.000 1873.920 1404.000 1874.270 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 399.810 1904.580 400.130 1904.640 ;
        RECT 1390.190 1904.580 1390.510 1904.640 ;
        RECT 399.810 1904.440 1390.510 1904.580 ;
        RECT 399.810 1904.380 400.130 1904.440 ;
        RECT 1390.190 1904.380 1390.510 1904.440 ;
        RECT 395.210 17.920 395.530 17.980 ;
        RECT 399.810 17.920 400.130 17.980 ;
        RECT 395.210 17.780 400.130 17.920 ;
        RECT 395.210 17.720 395.530 17.780 ;
        RECT 399.810 17.720 400.130 17.780 ;
      LAYER via ;
        RECT 399.840 1904.380 400.100 1904.640 ;
        RECT 1390.220 1904.380 1390.480 1904.640 ;
        RECT 395.240 17.720 395.500 17.980 ;
        RECT 399.840 17.720 400.100 17.980 ;
      LAYER met2 ;
        RECT 1390.210 1905.515 1390.490 1905.885 ;
        RECT 1390.280 1904.670 1390.420 1905.515 ;
        RECT 399.840 1904.350 400.100 1904.670 ;
        RECT 1390.220 1904.350 1390.480 1904.670 ;
        RECT 399.900 18.010 400.040 1904.350 ;
        RECT 395.240 17.690 395.500 18.010 ;
        RECT 399.840 17.690 400.100 18.010 ;
        RECT 395.300 2.400 395.440 17.690 ;
        RECT 395.090 -4.800 395.650 2.400 ;
      LAYER via2 ;
        RECT 1390.210 1905.560 1390.490 1905.840 ;
      LAYER met3 ;
        RECT 1390.185 1905.850 1390.515 1905.865 ;
        RECT 1390.185 1905.800 1400.700 1905.850 ;
        RECT 1390.185 1905.550 1404.000 1905.800 ;
        RECT 1390.185 1905.535 1390.515 1905.550 ;
        RECT 1400.000 1905.200 1404.000 1905.550 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.610 1932.120 413.930 1932.180 ;
        RECT 1389.270 1932.120 1389.590 1932.180 ;
        RECT 413.610 1931.980 1389.590 1932.120 ;
        RECT 413.610 1931.920 413.930 1931.980 ;
        RECT 1389.270 1931.920 1389.590 1931.980 ;
      LAYER via ;
        RECT 413.640 1931.920 413.900 1932.180 ;
        RECT 1389.300 1931.920 1389.560 1932.180 ;
      LAYER met2 ;
        RECT 1389.290 1937.475 1389.570 1937.845 ;
        RECT 1389.360 1932.210 1389.500 1937.475 ;
        RECT 413.640 1931.890 413.900 1932.210 ;
        RECT 1389.300 1931.890 1389.560 1932.210 ;
        RECT 413.700 17.410 413.840 1931.890 ;
        RECT 413.240 17.270 413.840 17.410 ;
        RECT 413.240 2.400 413.380 17.270 ;
        RECT 413.030 -4.800 413.590 2.400 ;
      LAYER via2 ;
        RECT 1389.290 1937.520 1389.570 1937.800 ;
      LAYER met3 ;
        RECT 1389.265 1937.810 1389.595 1937.825 ;
        RECT 1389.265 1937.760 1400.700 1937.810 ;
        RECT 1389.265 1937.510 1404.000 1937.760 ;
        RECT 1389.265 1937.495 1389.595 1937.510 ;
        RECT 1400.000 1937.160 1404.000 1937.510 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 75.510 1332.020 75.830 1332.080 ;
        RECT 1390.190 1332.020 1390.510 1332.080 ;
        RECT 75.510 1331.880 1390.510 1332.020 ;
        RECT 75.510 1331.820 75.830 1331.880 ;
        RECT 1390.190 1331.820 1390.510 1331.880 ;
      LAYER via ;
        RECT 75.540 1331.820 75.800 1332.080 ;
        RECT 1390.220 1331.820 1390.480 1332.080 ;
      LAYER met2 ;
        RECT 1390.210 1332.275 1390.490 1332.645 ;
        RECT 1390.280 1332.110 1390.420 1332.275 ;
        RECT 75.540 1331.790 75.800 1332.110 ;
        RECT 1390.220 1331.790 1390.480 1332.110 ;
        RECT 75.600 17.410 75.740 1331.790 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 1390.210 1332.320 1390.490 1332.600 ;
      LAYER met3 ;
        RECT 1390.185 1332.610 1390.515 1332.625 ;
        RECT 1390.185 1332.560 1400.700 1332.610 ;
        RECT 1390.185 1332.310 1404.000 1332.560 ;
        RECT 1390.185 1332.295 1390.515 1332.310 ;
        RECT 1400.000 1331.960 1404.000 1332.310 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.310 1966.800 434.630 1966.860 ;
        RECT 1393.410 1966.800 1393.730 1966.860 ;
        RECT 434.310 1966.660 1393.730 1966.800 ;
        RECT 434.310 1966.600 434.630 1966.660 ;
        RECT 1393.410 1966.600 1393.730 1966.660 ;
        RECT 430.630 17.920 430.950 17.980 ;
        RECT 434.310 17.920 434.630 17.980 ;
        RECT 430.630 17.780 434.630 17.920 ;
        RECT 430.630 17.720 430.950 17.780 ;
        RECT 434.310 17.720 434.630 17.780 ;
      LAYER via ;
        RECT 434.340 1966.600 434.600 1966.860 ;
        RECT 1393.440 1966.600 1393.700 1966.860 ;
        RECT 430.660 17.720 430.920 17.980 ;
        RECT 434.340 17.720 434.600 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1969.435 1393.710 1969.805 ;
        RECT 1393.500 1966.890 1393.640 1969.435 ;
        RECT 434.340 1966.570 434.600 1966.890 ;
        RECT 1393.440 1966.570 1393.700 1966.890 ;
        RECT 434.400 18.010 434.540 1966.570 ;
        RECT 430.660 17.690 430.920 18.010 ;
        RECT 434.340 17.690 434.600 18.010 ;
        RECT 430.720 2.400 430.860 17.690 ;
        RECT 430.510 -4.800 431.070 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1969.480 1393.710 1969.760 ;
      LAYER met3 ;
        RECT 1393.405 1969.770 1393.735 1969.785 ;
        RECT 1393.405 1969.720 1400.700 1969.770 ;
        RECT 1393.405 1969.470 1404.000 1969.720 ;
        RECT 1393.405 1969.455 1393.735 1969.470 ;
        RECT 1400.000 1969.120 1404.000 1969.470 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 454.550 2001.140 454.870 2001.200 ;
        RECT 1393.410 2001.140 1393.730 2001.200 ;
        RECT 454.550 2001.000 1393.730 2001.140 ;
        RECT 454.550 2000.940 454.870 2001.000 ;
        RECT 1393.410 2000.940 1393.730 2001.000 ;
        RECT 448.570 17.920 448.890 17.980 ;
        RECT 454.550 17.920 454.870 17.980 ;
        RECT 448.570 17.780 454.870 17.920 ;
        RECT 448.570 17.720 448.890 17.780 ;
        RECT 454.550 17.720 454.870 17.780 ;
      LAYER via ;
        RECT 454.580 2000.940 454.840 2001.200 ;
        RECT 1393.440 2000.940 1393.700 2001.200 ;
        RECT 448.600 17.720 448.860 17.980 ;
        RECT 454.580 17.720 454.840 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2001.395 1393.710 2001.765 ;
        RECT 1393.500 2001.230 1393.640 2001.395 ;
        RECT 454.580 2000.910 454.840 2001.230 ;
        RECT 1393.440 2000.910 1393.700 2001.230 ;
        RECT 454.640 18.010 454.780 2000.910 ;
        RECT 448.600 17.690 448.860 18.010 ;
        RECT 454.580 17.690 454.840 18.010 ;
        RECT 448.660 2.400 448.800 17.690 ;
        RECT 448.450 -4.800 449.010 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2001.440 1393.710 2001.720 ;
      LAYER met3 ;
        RECT 1393.405 2001.730 1393.735 2001.745 ;
        RECT 1393.405 2001.680 1400.700 2001.730 ;
        RECT 1393.405 2001.430 1404.000 2001.680 ;
        RECT 1393.405 2001.415 1393.735 2001.430 ;
        RECT 1400.000 2001.080 1404.000 2001.430 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 2028.680 469.130 2028.740 ;
        RECT 1393.410 2028.680 1393.730 2028.740 ;
        RECT 468.810 2028.540 1393.730 2028.680 ;
        RECT 468.810 2028.480 469.130 2028.540 ;
        RECT 1393.410 2028.480 1393.730 2028.540 ;
        RECT 466.510 17.920 466.830 17.980 ;
        RECT 468.810 17.920 469.130 17.980 ;
        RECT 466.510 17.780 469.130 17.920 ;
        RECT 466.510 17.720 466.830 17.780 ;
        RECT 468.810 17.720 469.130 17.780 ;
      LAYER via ;
        RECT 468.840 2028.480 469.100 2028.740 ;
        RECT 1393.440 2028.480 1393.700 2028.740 ;
        RECT 466.540 17.720 466.800 17.980 ;
        RECT 468.840 17.720 469.100 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2033.355 1393.710 2033.725 ;
        RECT 1393.500 2028.770 1393.640 2033.355 ;
        RECT 468.840 2028.450 469.100 2028.770 ;
        RECT 1393.440 2028.450 1393.700 2028.770 ;
        RECT 468.900 18.010 469.040 2028.450 ;
        RECT 466.540 17.690 466.800 18.010 ;
        RECT 468.840 17.690 469.100 18.010 ;
        RECT 466.600 2.400 466.740 17.690 ;
        RECT 466.390 -4.800 466.950 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2033.400 1393.710 2033.680 ;
      LAYER met3 ;
        RECT 1393.405 2033.690 1393.735 2033.705 ;
        RECT 1393.405 2033.640 1400.700 2033.690 ;
        RECT 1393.405 2033.390 1404.000 2033.640 ;
        RECT 1393.405 2033.375 1393.735 2033.390 ;
        RECT 1400.000 2033.040 1404.000 2033.390 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 489.510 2063.360 489.830 2063.420 ;
        RECT 1393.410 2063.360 1393.730 2063.420 ;
        RECT 489.510 2063.220 1393.730 2063.360 ;
        RECT 489.510 2063.160 489.830 2063.220 ;
        RECT 1393.410 2063.160 1393.730 2063.220 ;
        RECT 484.450 17.920 484.770 17.980 ;
        RECT 489.510 17.920 489.830 17.980 ;
        RECT 484.450 17.780 489.830 17.920 ;
        RECT 484.450 17.720 484.770 17.780 ;
        RECT 489.510 17.720 489.830 17.780 ;
      LAYER via ;
        RECT 489.540 2063.160 489.800 2063.420 ;
        RECT 1393.440 2063.160 1393.700 2063.420 ;
        RECT 484.480 17.720 484.740 17.980 ;
        RECT 489.540 17.720 489.800 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2065.315 1393.710 2065.685 ;
        RECT 1393.500 2063.450 1393.640 2065.315 ;
        RECT 489.540 2063.130 489.800 2063.450 ;
        RECT 1393.440 2063.130 1393.700 2063.450 ;
        RECT 489.600 18.010 489.740 2063.130 ;
        RECT 484.480 17.690 484.740 18.010 ;
        RECT 489.540 17.690 489.800 18.010 ;
        RECT 484.540 2.400 484.680 17.690 ;
        RECT 484.330 -4.800 484.890 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2065.360 1393.710 2065.640 ;
      LAYER met3 ;
        RECT 1393.405 2065.650 1393.735 2065.665 ;
        RECT 1393.405 2065.600 1400.700 2065.650 ;
        RECT 1393.405 2065.350 1404.000 2065.600 ;
        RECT 1393.405 2065.335 1393.735 2065.350 ;
        RECT 1400.000 2065.000 1404.000 2065.350 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 2090.900 503.630 2090.960 ;
        RECT 1393.410 2090.900 1393.730 2090.960 ;
        RECT 503.310 2090.760 1393.730 2090.900 ;
        RECT 503.310 2090.700 503.630 2090.760 ;
        RECT 1393.410 2090.700 1393.730 2090.760 ;
      LAYER via ;
        RECT 503.340 2090.700 503.600 2090.960 ;
        RECT 1393.440 2090.700 1393.700 2090.960 ;
      LAYER met2 ;
        RECT 1393.430 2097.275 1393.710 2097.645 ;
        RECT 1393.500 2090.990 1393.640 2097.275 ;
        RECT 503.340 2090.670 503.600 2090.990 ;
        RECT 1393.440 2090.670 1393.700 2090.990 ;
        RECT 503.400 17.410 503.540 2090.670 ;
        RECT 502.480 17.270 503.540 17.410 ;
        RECT 502.480 2.400 502.620 17.270 ;
        RECT 502.270 -4.800 502.830 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2097.320 1393.710 2097.600 ;
      LAYER met3 ;
        RECT 1393.405 2097.610 1393.735 2097.625 ;
        RECT 1393.405 2097.560 1400.700 2097.610 ;
        RECT 1393.405 2097.310 1404.000 2097.560 ;
        RECT 1393.405 2097.295 1393.735 2097.310 ;
        RECT 1400.000 2096.960 1404.000 2097.310 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 2125.580 524.330 2125.640 ;
        RECT 1393.410 2125.580 1393.730 2125.640 ;
        RECT 524.010 2125.440 1393.730 2125.580 ;
        RECT 524.010 2125.380 524.330 2125.440 ;
        RECT 1393.410 2125.380 1393.730 2125.440 ;
        RECT 519.870 17.920 520.190 17.980 ;
        RECT 524.010 17.920 524.330 17.980 ;
        RECT 519.870 17.780 524.330 17.920 ;
        RECT 519.870 17.720 520.190 17.780 ;
        RECT 524.010 17.720 524.330 17.780 ;
      LAYER via ;
        RECT 524.040 2125.380 524.300 2125.640 ;
        RECT 1393.440 2125.380 1393.700 2125.640 ;
        RECT 519.900 17.720 520.160 17.980 ;
        RECT 524.040 17.720 524.300 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2128.555 1393.710 2128.925 ;
        RECT 1393.500 2125.670 1393.640 2128.555 ;
        RECT 524.040 2125.350 524.300 2125.670 ;
        RECT 1393.440 2125.350 1393.700 2125.670 ;
        RECT 524.100 18.010 524.240 2125.350 ;
        RECT 519.900 17.690 520.160 18.010 ;
        RECT 524.040 17.690 524.300 18.010 ;
        RECT 519.960 2.400 520.100 17.690 ;
        RECT 519.750 -4.800 520.310 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2128.600 1393.710 2128.880 ;
      LAYER met3 ;
        RECT 1393.405 2128.890 1393.735 2128.905 ;
        RECT 1393.405 2128.840 1400.700 2128.890 ;
        RECT 1393.405 2128.590 1404.000 2128.840 ;
        RECT 1393.405 2128.575 1393.735 2128.590 ;
        RECT 1400.000 2128.240 1404.000 2128.590 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 2159.920 538.130 2159.980 ;
        RECT 1393.410 2159.920 1393.730 2159.980 ;
        RECT 537.810 2159.780 1393.730 2159.920 ;
        RECT 537.810 2159.720 538.130 2159.780 ;
        RECT 1393.410 2159.720 1393.730 2159.780 ;
      LAYER via ;
        RECT 537.840 2159.720 538.100 2159.980 ;
        RECT 1393.440 2159.720 1393.700 2159.980 ;
      LAYER met2 ;
        RECT 1393.430 2160.515 1393.710 2160.885 ;
        RECT 1393.500 2160.010 1393.640 2160.515 ;
        RECT 537.840 2159.690 538.100 2160.010 ;
        RECT 1393.440 2159.690 1393.700 2160.010 ;
        RECT 537.900 2.400 538.040 2159.690 ;
        RECT 537.690 -4.800 538.250 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2160.560 1393.710 2160.840 ;
      LAYER met3 ;
        RECT 1393.405 2160.850 1393.735 2160.865 ;
        RECT 1393.405 2160.800 1400.700 2160.850 ;
        RECT 1393.405 2160.550 1404.000 2160.800 ;
        RECT 1393.405 2160.535 1393.735 2160.550 ;
        RECT 1400.000 2160.200 1404.000 2160.550 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 558.510 2187.460 558.830 2187.520 ;
        RECT 1393.410 2187.460 1393.730 2187.520 ;
        RECT 558.510 2187.320 1393.730 2187.460 ;
        RECT 558.510 2187.260 558.830 2187.320 ;
        RECT 1393.410 2187.260 1393.730 2187.320 ;
        RECT 555.750 17.920 556.070 17.980 ;
        RECT 558.510 17.920 558.830 17.980 ;
        RECT 555.750 17.780 558.830 17.920 ;
        RECT 555.750 17.720 556.070 17.780 ;
        RECT 558.510 17.720 558.830 17.780 ;
      LAYER via ;
        RECT 558.540 2187.260 558.800 2187.520 ;
        RECT 1393.440 2187.260 1393.700 2187.520 ;
        RECT 555.780 17.720 556.040 17.980 ;
        RECT 558.540 17.720 558.800 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2192.475 1393.710 2192.845 ;
        RECT 1393.500 2187.550 1393.640 2192.475 ;
        RECT 558.540 2187.230 558.800 2187.550 ;
        RECT 1393.440 2187.230 1393.700 2187.550 ;
        RECT 558.600 18.010 558.740 2187.230 ;
        RECT 555.780 17.690 556.040 18.010 ;
        RECT 558.540 17.690 558.800 18.010 ;
        RECT 555.840 2.400 555.980 17.690 ;
        RECT 555.630 -4.800 556.190 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2192.520 1393.710 2192.800 ;
      LAYER met3 ;
        RECT 1393.405 2192.810 1393.735 2192.825 ;
        RECT 1393.405 2192.760 1400.700 2192.810 ;
        RECT 1393.405 2192.510 1404.000 2192.760 ;
        RECT 1393.405 2192.495 1393.735 2192.510 ;
        RECT 1400.000 2192.160 1404.000 2192.510 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 579.210 2222.140 579.530 2222.200 ;
        RECT 1393.410 2222.140 1393.730 2222.200 ;
        RECT 579.210 2222.000 1393.730 2222.140 ;
        RECT 579.210 2221.940 579.530 2222.000 ;
        RECT 1393.410 2221.940 1393.730 2222.000 ;
        RECT 573.690 17.920 574.010 17.980 ;
        RECT 579.210 17.920 579.530 17.980 ;
        RECT 573.690 17.780 579.530 17.920 ;
        RECT 573.690 17.720 574.010 17.780 ;
        RECT 579.210 17.720 579.530 17.780 ;
      LAYER via ;
        RECT 579.240 2221.940 579.500 2222.200 ;
        RECT 1393.440 2221.940 1393.700 2222.200 ;
        RECT 573.720 17.720 573.980 17.980 ;
        RECT 579.240 17.720 579.500 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2224.435 1393.710 2224.805 ;
        RECT 1393.500 2222.230 1393.640 2224.435 ;
        RECT 579.240 2221.910 579.500 2222.230 ;
        RECT 1393.440 2221.910 1393.700 2222.230 ;
        RECT 579.300 18.010 579.440 2221.910 ;
        RECT 573.720 17.690 573.980 18.010 ;
        RECT 579.240 17.690 579.500 18.010 ;
        RECT 573.780 2.400 573.920 17.690 ;
        RECT 573.570 -4.800 574.130 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2224.480 1393.710 2224.760 ;
      LAYER met3 ;
        RECT 1393.405 2224.770 1393.735 2224.785 ;
        RECT 1393.405 2224.720 1400.700 2224.770 ;
        RECT 1393.405 2224.470 1404.000 2224.720 ;
        RECT 1393.405 2224.455 1393.735 2224.470 ;
        RECT 1400.000 2224.120 1404.000 2224.470 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 2256.480 593.330 2256.540 ;
        RECT 1393.410 2256.480 1393.730 2256.540 ;
        RECT 593.010 2256.340 1393.730 2256.480 ;
        RECT 593.010 2256.280 593.330 2256.340 ;
        RECT 1393.410 2256.280 1393.730 2256.340 ;
      LAYER via ;
        RECT 593.040 2256.280 593.300 2256.540 ;
        RECT 1393.440 2256.280 1393.700 2256.540 ;
      LAYER met2 ;
        RECT 593.040 2256.250 593.300 2256.570 ;
        RECT 1393.430 2256.395 1393.710 2256.765 ;
        RECT 1393.440 2256.250 1393.700 2256.395 ;
        RECT 593.100 17.410 593.240 2256.250 ;
        RECT 591.260 17.270 593.240 17.410 ;
        RECT 591.260 2.400 591.400 17.270 ;
        RECT 591.050 -4.800 591.610 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2256.440 1393.710 2256.720 ;
      LAYER met3 ;
        RECT 1393.405 2256.730 1393.735 2256.745 ;
        RECT 1393.405 2256.680 1400.700 2256.730 ;
        RECT 1393.405 2256.430 1404.000 2256.680 ;
        RECT 1393.405 2256.415 1393.735 2256.430 ;
        RECT 1400.000 2256.080 1404.000 2256.430 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 103.110 1373.500 103.430 1373.560 ;
        RECT 1390.190 1373.500 1390.510 1373.560 ;
        RECT 103.110 1373.360 1390.510 1373.500 ;
        RECT 103.110 1373.300 103.430 1373.360 ;
        RECT 1390.190 1373.300 1390.510 1373.360 ;
        RECT 97.590 17.920 97.910 17.980 ;
        RECT 103.110 17.920 103.430 17.980 ;
        RECT 97.590 17.780 103.430 17.920 ;
        RECT 97.590 17.720 97.910 17.780 ;
        RECT 103.110 17.720 103.430 17.780 ;
      LAYER via ;
        RECT 103.140 1373.300 103.400 1373.560 ;
        RECT 1390.220 1373.300 1390.480 1373.560 ;
        RECT 97.620 17.720 97.880 17.980 ;
        RECT 103.140 17.720 103.400 17.980 ;
      LAYER met2 ;
        RECT 1390.210 1374.435 1390.490 1374.805 ;
        RECT 1390.280 1373.590 1390.420 1374.435 ;
        RECT 103.140 1373.270 103.400 1373.590 ;
        RECT 1390.220 1373.270 1390.480 1373.590 ;
        RECT 103.200 18.010 103.340 1373.270 ;
        RECT 97.620 17.690 97.880 18.010 ;
        RECT 103.140 17.690 103.400 18.010 ;
        RECT 97.680 2.400 97.820 17.690 ;
        RECT 97.470 -4.800 98.030 2.400 ;
      LAYER via2 ;
        RECT 1390.210 1374.480 1390.490 1374.760 ;
      LAYER met3 ;
        RECT 1390.185 1374.770 1390.515 1374.785 ;
        RECT 1390.185 1374.720 1400.700 1374.770 ;
        RECT 1390.185 1374.470 1404.000 1374.720 ;
        RECT 1390.185 1374.455 1390.515 1374.470 ;
        RECT 1400.000 1374.120 1404.000 1374.470 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 613.710 2284.020 614.030 2284.080 ;
        RECT 1393.410 2284.020 1393.730 2284.080 ;
        RECT 613.710 2283.880 1393.730 2284.020 ;
        RECT 613.710 2283.820 614.030 2283.880 ;
        RECT 1393.410 2283.820 1393.730 2283.880 ;
        RECT 609.110 17.920 609.430 17.980 ;
        RECT 613.710 17.920 614.030 17.980 ;
        RECT 609.110 17.780 614.030 17.920 ;
        RECT 609.110 17.720 609.430 17.780 ;
        RECT 613.710 17.720 614.030 17.780 ;
      LAYER via ;
        RECT 613.740 2283.820 614.000 2284.080 ;
        RECT 1393.440 2283.820 1393.700 2284.080 ;
        RECT 609.140 17.720 609.400 17.980 ;
        RECT 613.740 17.720 614.000 17.980 ;
      LAYER met2 ;
        RECT 1393.430 2288.355 1393.710 2288.725 ;
        RECT 1393.500 2284.110 1393.640 2288.355 ;
        RECT 613.740 2283.790 614.000 2284.110 ;
        RECT 1393.440 2283.790 1393.700 2284.110 ;
        RECT 613.800 18.010 613.940 2283.790 ;
        RECT 609.140 17.690 609.400 18.010 ;
        RECT 613.740 17.690 614.000 18.010 ;
        RECT 609.200 2.400 609.340 17.690 ;
        RECT 608.990 -4.800 609.550 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2288.400 1393.710 2288.680 ;
      LAYER met3 ;
        RECT 1393.405 2288.690 1393.735 2288.705 ;
        RECT 1393.405 2288.640 1400.700 2288.690 ;
        RECT 1393.405 2288.390 1404.000 2288.640 ;
        RECT 1393.405 2288.375 1393.735 2288.390 ;
        RECT 1400.000 2288.040 1404.000 2288.390 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 2318.700 627.830 2318.760 ;
        RECT 1393.410 2318.700 1393.730 2318.760 ;
        RECT 627.510 2318.560 1393.730 2318.700 ;
        RECT 627.510 2318.500 627.830 2318.560 ;
        RECT 1393.410 2318.500 1393.730 2318.560 ;
      LAYER via ;
        RECT 627.540 2318.500 627.800 2318.760 ;
        RECT 1393.440 2318.500 1393.700 2318.760 ;
      LAYER met2 ;
        RECT 1393.430 2320.315 1393.710 2320.685 ;
        RECT 1393.500 2318.790 1393.640 2320.315 ;
        RECT 627.540 2318.470 627.800 2318.790 ;
        RECT 1393.440 2318.470 1393.700 2318.790 ;
        RECT 627.600 17.410 627.740 2318.470 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
      LAYER via2 ;
        RECT 1393.430 2320.360 1393.710 2320.640 ;
      LAYER met3 ;
        RECT 1393.405 2320.650 1393.735 2320.665 ;
        RECT 1393.405 2320.600 1400.700 2320.650 ;
        RECT 1393.405 2320.350 1404.000 2320.600 ;
        RECT 1393.405 2320.335 1393.735 2320.350 ;
        RECT 1400.000 2320.000 1404.000 2320.350 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 123.810 1414.640 124.130 1414.700 ;
        RECT 1393.410 1414.640 1393.730 1414.700 ;
        RECT 123.810 1414.500 1393.730 1414.640 ;
        RECT 123.810 1414.440 124.130 1414.500 ;
        RECT 1393.410 1414.440 1393.730 1414.500 ;
        RECT 121.510 17.920 121.830 17.980 ;
        RECT 123.810 17.920 124.130 17.980 ;
        RECT 121.510 17.780 124.130 17.920 ;
        RECT 121.510 17.720 121.830 17.780 ;
        RECT 123.810 17.720 124.130 17.780 ;
      LAYER via ;
        RECT 123.840 1414.440 124.100 1414.700 ;
        RECT 1393.440 1414.440 1393.700 1414.700 ;
        RECT 121.540 17.720 121.800 17.980 ;
        RECT 123.840 17.720 124.100 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1417.275 1393.710 1417.645 ;
        RECT 1393.500 1414.730 1393.640 1417.275 ;
        RECT 123.840 1414.410 124.100 1414.730 ;
        RECT 1393.440 1414.410 1393.700 1414.730 ;
        RECT 123.900 18.010 124.040 1414.410 ;
        RECT 121.540 17.690 121.800 18.010 ;
        RECT 123.840 17.690 124.100 18.010 ;
        RECT 121.600 2.400 121.740 17.690 ;
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1417.320 1393.710 1417.600 ;
      LAYER met3 ;
        RECT 1393.405 1417.610 1393.735 1417.625 ;
        RECT 1393.405 1417.560 1400.700 1417.610 ;
        RECT 1393.405 1417.310 1404.000 1417.560 ;
        RECT 1393.405 1417.295 1393.735 1417.310 ;
        RECT 1400.000 1416.960 1404.000 1417.310 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 150.950 1456.120 151.270 1456.180 ;
        RECT 1393.410 1456.120 1393.730 1456.180 ;
        RECT 150.950 1455.980 1393.730 1456.120 ;
        RECT 150.950 1455.920 151.270 1455.980 ;
        RECT 1393.410 1455.920 1393.730 1455.980 ;
        RECT 145.430 17.920 145.750 17.980 ;
        RECT 150.950 17.920 151.270 17.980 ;
        RECT 145.430 17.780 151.270 17.920 ;
        RECT 145.430 17.720 145.750 17.780 ;
        RECT 150.950 17.720 151.270 17.780 ;
      LAYER via ;
        RECT 150.980 1455.920 151.240 1456.180 ;
        RECT 1393.440 1455.920 1393.700 1456.180 ;
        RECT 145.460 17.720 145.720 17.980 ;
        RECT 150.980 17.720 151.240 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1459.435 1393.710 1459.805 ;
        RECT 1393.500 1456.210 1393.640 1459.435 ;
        RECT 150.980 1455.890 151.240 1456.210 ;
        RECT 1393.440 1455.890 1393.700 1456.210 ;
        RECT 151.040 18.010 151.180 1455.890 ;
        RECT 145.460 17.690 145.720 18.010 ;
        RECT 150.980 17.690 151.240 18.010 ;
        RECT 145.520 2.400 145.660 17.690 ;
        RECT 145.310 -4.800 145.870 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1459.480 1393.710 1459.760 ;
      LAYER met3 ;
        RECT 1393.405 1459.770 1393.735 1459.785 ;
        RECT 1393.405 1459.720 1400.700 1459.770 ;
        RECT 1393.405 1459.470 1404.000 1459.720 ;
        RECT 1393.405 1459.455 1393.735 1459.470 ;
        RECT 1400.000 1459.120 1404.000 1459.470 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 165.210 1490.800 165.530 1490.860 ;
        RECT 1393.410 1490.800 1393.730 1490.860 ;
        RECT 165.210 1490.660 1393.730 1490.800 ;
        RECT 165.210 1490.600 165.530 1490.660 ;
        RECT 1393.410 1490.600 1393.730 1490.660 ;
      LAYER via ;
        RECT 165.240 1490.600 165.500 1490.860 ;
        RECT 1393.440 1490.600 1393.700 1490.860 ;
      LAYER met2 ;
        RECT 1393.430 1491.395 1393.710 1491.765 ;
        RECT 1393.500 1490.890 1393.640 1491.395 ;
        RECT 165.240 1490.570 165.500 1490.890 ;
        RECT 1393.440 1490.570 1393.700 1490.890 ;
        RECT 165.300 17.410 165.440 1490.570 ;
        RECT 163.460 17.270 165.440 17.410 ;
        RECT 163.460 2.400 163.600 17.270 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1491.440 1393.710 1491.720 ;
      LAYER met3 ;
        RECT 1393.405 1491.730 1393.735 1491.745 ;
        RECT 1393.405 1491.680 1400.700 1491.730 ;
        RECT 1393.405 1491.430 1404.000 1491.680 ;
        RECT 1393.405 1491.415 1393.735 1491.430 ;
        RECT 1400.000 1491.080 1404.000 1491.430 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 185.910 1518.340 186.230 1518.400 ;
        RECT 1393.410 1518.340 1393.730 1518.400 ;
        RECT 185.910 1518.200 1393.730 1518.340 ;
        RECT 185.910 1518.140 186.230 1518.200 ;
        RECT 1393.410 1518.140 1393.730 1518.200 ;
        RECT 180.850 17.920 181.170 17.980 ;
        RECT 185.910 17.920 186.230 17.980 ;
        RECT 180.850 17.780 186.230 17.920 ;
        RECT 180.850 17.720 181.170 17.780 ;
        RECT 185.910 17.720 186.230 17.780 ;
      LAYER via ;
        RECT 185.940 1518.140 186.200 1518.400 ;
        RECT 1393.440 1518.140 1393.700 1518.400 ;
        RECT 180.880 17.720 181.140 17.980 ;
        RECT 185.940 17.720 186.200 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1523.355 1393.710 1523.725 ;
        RECT 1393.500 1518.430 1393.640 1523.355 ;
        RECT 185.940 1518.110 186.200 1518.430 ;
        RECT 1393.440 1518.110 1393.700 1518.430 ;
        RECT 186.000 18.010 186.140 1518.110 ;
        RECT 180.880 17.690 181.140 18.010 ;
        RECT 185.940 17.690 186.200 18.010 ;
        RECT 180.940 2.400 181.080 17.690 ;
        RECT 180.730 -4.800 181.290 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1523.400 1393.710 1523.680 ;
      LAYER met3 ;
        RECT 1393.405 1523.690 1393.735 1523.705 ;
        RECT 1393.405 1523.640 1400.700 1523.690 ;
        RECT 1393.405 1523.390 1404.000 1523.640 ;
        RECT 1393.405 1523.375 1393.735 1523.390 ;
        RECT 1400.000 1523.040 1404.000 1523.390 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 199.710 1552.680 200.030 1552.740 ;
        RECT 1393.410 1552.680 1393.730 1552.740 ;
        RECT 199.710 1552.540 1393.730 1552.680 ;
        RECT 199.710 1552.480 200.030 1552.540 ;
        RECT 1393.410 1552.480 1393.730 1552.540 ;
      LAYER via ;
        RECT 199.740 1552.480 200.000 1552.740 ;
        RECT 1393.440 1552.480 1393.700 1552.740 ;
      LAYER met2 ;
        RECT 1393.430 1555.315 1393.710 1555.685 ;
        RECT 1393.500 1552.770 1393.640 1555.315 ;
        RECT 199.740 1552.450 200.000 1552.770 ;
        RECT 1393.440 1552.450 1393.700 1552.770 ;
        RECT 199.800 17.410 199.940 1552.450 ;
        RECT 198.880 17.270 199.940 17.410 ;
        RECT 198.880 2.400 199.020 17.270 ;
        RECT 198.670 -4.800 199.230 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1555.360 1393.710 1555.640 ;
      LAYER met3 ;
        RECT 1393.405 1555.650 1393.735 1555.665 ;
        RECT 1393.405 1555.600 1400.700 1555.650 ;
        RECT 1393.405 1555.350 1404.000 1555.600 ;
        RECT 1393.405 1555.335 1393.735 1555.350 ;
        RECT 1400.000 1555.000 1404.000 1555.350 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 220.410 1587.360 220.730 1587.420 ;
        RECT 1393.410 1587.360 1393.730 1587.420 ;
        RECT 220.410 1587.220 1393.730 1587.360 ;
        RECT 220.410 1587.160 220.730 1587.220 ;
        RECT 1393.410 1587.160 1393.730 1587.220 ;
        RECT 216.730 17.920 217.050 17.980 ;
        RECT 220.410 17.920 220.730 17.980 ;
        RECT 216.730 17.780 220.730 17.920 ;
        RECT 216.730 17.720 217.050 17.780 ;
        RECT 220.410 17.720 220.730 17.780 ;
      LAYER via ;
        RECT 220.440 1587.160 220.700 1587.420 ;
        RECT 1393.440 1587.160 1393.700 1587.420 ;
        RECT 216.760 17.720 217.020 17.980 ;
        RECT 220.440 17.720 220.700 17.980 ;
      LAYER met2 ;
        RECT 220.440 1587.130 220.700 1587.450 ;
        RECT 1393.430 1587.275 1393.710 1587.645 ;
        RECT 1393.440 1587.130 1393.700 1587.275 ;
        RECT 220.500 18.010 220.640 1587.130 ;
        RECT 216.760 17.690 217.020 18.010 ;
        RECT 220.440 17.690 220.700 18.010 ;
        RECT 216.820 2.400 216.960 17.690 ;
        RECT 216.610 -4.800 217.170 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1587.320 1393.710 1587.600 ;
      LAYER met3 ;
        RECT 1393.405 1587.610 1393.735 1587.625 ;
        RECT 1393.405 1587.560 1400.700 1587.610 ;
        RECT 1393.405 1587.310 1404.000 1587.560 ;
        RECT 1393.405 1587.295 1393.735 1587.310 ;
        RECT 1400.000 1586.960 1404.000 1587.310 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 240.650 1614.900 240.970 1614.960 ;
        RECT 1388.350 1614.900 1388.670 1614.960 ;
        RECT 240.650 1614.760 1388.670 1614.900 ;
        RECT 240.650 1614.700 240.970 1614.760 ;
        RECT 1388.350 1614.700 1388.670 1614.760 ;
        RECT 234.670 17.920 234.990 17.980 ;
        RECT 240.650 17.920 240.970 17.980 ;
        RECT 234.670 17.780 240.970 17.920 ;
        RECT 234.670 17.720 234.990 17.780 ;
        RECT 240.650 17.720 240.970 17.780 ;
      LAYER via ;
        RECT 240.680 1614.700 240.940 1614.960 ;
        RECT 1388.380 1614.700 1388.640 1614.960 ;
        RECT 234.700 17.720 234.960 17.980 ;
        RECT 240.680 17.720 240.940 17.980 ;
      LAYER met2 ;
        RECT 1388.370 1619.235 1388.650 1619.605 ;
        RECT 1388.440 1614.990 1388.580 1619.235 ;
        RECT 240.680 1614.670 240.940 1614.990 ;
        RECT 1388.380 1614.670 1388.640 1614.990 ;
        RECT 240.740 18.010 240.880 1614.670 ;
        RECT 234.700 17.690 234.960 18.010 ;
        RECT 240.680 17.690 240.940 18.010 ;
        RECT 234.760 2.400 234.900 17.690 ;
        RECT 234.550 -4.800 235.110 2.400 ;
      LAYER via2 ;
        RECT 1388.370 1619.280 1388.650 1619.560 ;
      LAYER met3 ;
        RECT 1388.345 1619.570 1388.675 1619.585 ;
        RECT 1388.345 1619.520 1400.700 1619.570 ;
        RECT 1388.345 1619.270 1404.000 1619.520 ;
        RECT 1388.345 1619.255 1388.675 1619.270 ;
        RECT 1400.000 1618.920 1404.000 1619.270 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 61.710 1297.340 62.030 1297.400 ;
        RECT 1391.570 1297.340 1391.890 1297.400 ;
        RECT 61.710 1297.200 1391.890 1297.340 ;
        RECT 61.710 1297.140 62.030 1297.200 ;
        RECT 1391.570 1297.140 1391.890 1297.200 ;
        RECT 56.190 17.920 56.510 17.980 ;
        RECT 61.710 17.920 62.030 17.980 ;
        RECT 56.190 17.780 62.030 17.920 ;
        RECT 56.190 17.720 56.510 17.780 ;
        RECT 61.710 17.720 62.030 17.780 ;
      LAYER via ;
        RECT 61.740 1297.140 62.000 1297.400 ;
        RECT 1391.600 1297.140 1391.860 1297.400 ;
        RECT 56.220 17.720 56.480 17.980 ;
        RECT 61.740 17.720 62.000 17.980 ;
      LAYER met2 ;
        RECT 1391.590 1300.315 1391.870 1300.685 ;
        RECT 1391.660 1297.430 1391.800 1300.315 ;
        RECT 61.740 1297.110 62.000 1297.430 ;
        RECT 1391.600 1297.110 1391.860 1297.430 ;
        RECT 61.800 18.010 61.940 1297.110 ;
        RECT 56.220 17.690 56.480 18.010 ;
        RECT 61.740 17.690 62.000 18.010 ;
        RECT 56.280 2.400 56.420 17.690 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 1391.590 1300.360 1391.870 1300.640 ;
      LAYER met3 ;
        RECT 1391.565 1300.650 1391.895 1300.665 ;
        RECT 1391.565 1300.600 1400.700 1300.650 ;
        RECT 1391.565 1300.350 1404.000 1300.600 ;
        RECT 1391.565 1300.335 1391.895 1300.350 ;
        RECT 1400.000 1300.000 1404.000 1300.350 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 1338.820 82.730 1338.880 ;
        RECT 1393.410 1338.820 1393.730 1338.880 ;
        RECT 82.410 1338.680 1393.730 1338.820 ;
        RECT 82.410 1338.620 82.730 1338.680 ;
        RECT 1393.410 1338.620 1393.730 1338.680 ;
        RECT 80.110 17.920 80.430 17.980 ;
        RECT 82.410 17.920 82.730 17.980 ;
        RECT 80.110 17.780 82.730 17.920 ;
        RECT 80.110 17.720 80.430 17.780 ;
        RECT 82.410 17.720 82.730 17.780 ;
      LAYER via ;
        RECT 82.440 1338.620 82.700 1338.880 ;
        RECT 1393.440 1338.620 1393.700 1338.880 ;
        RECT 80.140 17.720 80.400 17.980 ;
        RECT 82.440 17.720 82.700 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1343.155 1393.710 1343.525 ;
        RECT 1393.500 1338.910 1393.640 1343.155 ;
        RECT 82.440 1338.590 82.700 1338.910 ;
        RECT 1393.440 1338.590 1393.700 1338.910 ;
        RECT 82.500 18.010 82.640 1338.590 ;
        RECT 80.140 17.690 80.400 18.010 ;
        RECT 82.440 17.690 82.700 18.010 ;
        RECT 80.200 2.400 80.340 17.690 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1343.200 1393.710 1343.480 ;
      LAYER met3 ;
        RECT 1393.405 1343.490 1393.735 1343.505 ;
        RECT 1393.405 1343.440 1400.700 1343.490 ;
        RECT 1393.405 1343.190 1404.000 1343.440 ;
        RECT 1393.405 1343.175 1393.735 1343.190 ;
        RECT 1400.000 1342.840 1404.000 1343.190 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 1380.300 109.870 1380.360 ;
        RECT 1393.410 1380.300 1393.730 1380.360 ;
        RECT 109.550 1380.160 1393.730 1380.300 ;
        RECT 109.550 1380.100 109.870 1380.160 ;
        RECT 1393.410 1380.100 1393.730 1380.160 ;
        RECT 103.570 17.920 103.890 17.980 ;
        RECT 109.550 17.920 109.870 17.980 ;
        RECT 103.570 17.780 109.870 17.920 ;
        RECT 103.570 17.720 103.890 17.780 ;
        RECT 109.550 17.720 109.870 17.780 ;
      LAYER via ;
        RECT 109.580 1380.100 109.840 1380.360 ;
        RECT 1393.440 1380.100 1393.700 1380.360 ;
        RECT 103.600 17.720 103.860 17.980 ;
        RECT 109.580 17.720 109.840 17.980 ;
      LAYER met2 ;
        RECT 1393.430 1385.315 1393.710 1385.685 ;
        RECT 1393.500 1380.390 1393.640 1385.315 ;
        RECT 109.580 1380.070 109.840 1380.390 ;
        RECT 1393.440 1380.070 1393.700 1380.390 ;
        RECT 109.640 18.010 109.780 1380.070 ;
        RECT 103.600 17.690 103.860 18.010 ;
        RECT 109.580 17.690 109.840 18.010 ;
        RECT 103.660 2.400 103.800 17.690 ;
        RECT 103.450 -4.800 104.010 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1385.360 1393.710 1385.640 ;
      LAYER met3 ;
        RECT 1393.405 1385.650 1393.735 1385.665 ;
        RECT 1393.405 1385.600 1400.700 1385.650 ;
        RECT 1393.405 1385.350 1404.000 1385.600 ;
        RECT 1393.405 1385.335 1393.735 1385.350 ;
        RECT 1400.000 1385.000 1404.000 1385.350 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 130.710 1428.580 131.030 1428.640 ;
        RECT 1393.410 1428.580 1393.730 1428.640 ;
        RECT 130.710 1428.440 1393.730 1428.580 ;
        RECT 130.710 1428.380 131.030 1428.440 ;
        RECT 1393.410 1428.380 1393.730 1428.440 ;
        RECT 127.490 17.920 127.810 17.980 ;
        RECT 130.710 17.920 131.030 17.980 ;
        RECT 127.490 17.780 131.030 17.920 ;
        RECT 127.490 17.720 127.810 17.780 ;
        RECT 130.710 17.720 131.030 17.780 ;
      LAYER via ;
        RECT 130.740 1428.380 131.000 1428.640 ;
        RECT 1393.440 1428.380 1393.700 1428.640 ;
        RECT 127.520 17.720 127.780 17.980 ;
        RECT 130.740 17.720 131.000 17.980 ;
      LAYER met2 ;
        RECT 130.740 1428.350 131.000 1428.670 ;
        RECT 1393.440 1428.525 1393.700 1428.670 ;
        RECT 130.800 18.010 130.940 1428.350 ;
        RECT 1393.430 1428.155 1393.710 1428.525 ;
        RECT 127.520 17.690 127.780 18.010 ;
        RECT 130.740 17.690 131.000 18.010 ;
        RECT 127.580 2.400 127.720 17.690 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1428.200 1393.710 1428.480 ;
      LAYER met3 ;
        RECT 1393.405 1428.490 1393.735 1428.505 ;
        RECT 1393.405 1428.440 1400.700 1428.490 ;
        RECT 1393.405 1428.190 1404.000 1428.440 ;
        RECT 1393.405 1428.175 1393.735 1428.190 ;
        RECT 1400.000 1427.840 1404.000 1428.190 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.210 1242.260 27.530 1242.320 ;
        RECT 1393.410 1242.260 1393.730 1242.320 ;
        RECT 27.210 1242.120 1393.730 1242.260 ;
        RECT 27.210 1242.060 27.530 1242.120 ;
        RECT 1393.410 1242.060 1393.730 1242.120 ;
        RECT 26.290 2.960 26.610 3.020 ;
        RECT 27.210 2.960 27.530 3.020 ;
        RECT 26.290 2.820 27.530 2.960 ;
        RECT 26.290 2.760 26.610 2.820 ;
        RECT 27.210 2.760 27.530 2.820 ;
      LAYER via ;
        RECT 27.240 1242.060 27.500 1242.320 ;
        RECT 1393.440 1242.060 1393.700 1242.320 ;
        RECT 26.320 2.760 26.580 3.020 ;
        RECT 27.240 2.760 27.500 3.020 ;
      LAYER met2 ;
        RECT 1393.430 1247.275 1393.710 1247.645 ;
        RECT 1393.500 1242.350 1393.640 1247.275 ;
        RECT 27.240 1242.030 27.500 1242.350 ;
        RECT 1393.440 1242.030 1393.700 1242.350 ;
        RECT 27.300 3.050 27.440 1242.030 ;
        RECT 26.320 2.730 26.580 3.050 ;
        RECT 27.240 2.730 27.500 3.050 ;
        RECT 26.380 2.400 26.520 2.730 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1247.320 1393.710 1247.600 ;
      LAYER met3 ;
        RECT 1393.405 1247.610 1393.735 1247.625 ;
        RECT 1393.405 1247.560 1400.700 1247.610 ;
        RECT 1393.405 1247.310 1404.000 1247.560 ;
        RECT 1393.405 1247.295 1393.735 1247.310 ;
        RECT 1400.000 1246.960 1404.000 1247.310 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.110 1256.200 34.430 1256.260 ;
        RECT 1393.410 1256.200 1393.730 1256.260 ;
        RECT 34.110 1256.060 1393.730 1256.200 ;
        RECT 34.110 1256.000 34.430 1256.060 ;
        RECT 1393.410 1256.000 1393.730 1256.060 ;
      LAYER via ;
        RECT 34.140 1256.000 34.400 1256.260 ;
        RECT 1393.440 1256.000 1393.700 1256.260 ;
      LAYER met2 ;
        RECT 1393.430 1258.155 1393.710 1258.525 ;
        RECT 1393.500 1256.290 1393.640 1258.155 ;
        RECT 34.140 1255.970 34.400 1256.290 ;
        RECT 1393.440 1255.970 1393.700 1256.290 ;
        RECT 34.200 3.130 34.340 1255.970 ;
        RECT 32.360 2.990 34.340 3.130 ;
        RECT 32.360 2.400 32.500 2.990 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 1393.430 1258.200 1393.710 1258.480 ;
      LAYER met3 ;
        RECT 1393.405 1258.490 1393.735 1258.505 ;
        RECT 1393.405 1258.440 1400.700 1258.490 ;
        RECT 1393.405 1258.190 1404.000 1258.440 ;
        RECT 1393.405 1258.175 1393.735 1258.190 ;
        RECT 1400.000 1257.840 1404.000 1258.190 ;
    END
  END wbs_we_i
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1406.750 1190.580 1407.070 1190.640 ;
        RECT 1486.790 1190.580 1487.110 1190.640 ;
        RECT 1406.750 1190.440 1487.110 1190.580 ;
        RECT 1406.750 1190.380 1407.070 1190.440 ;
        RECT 1486.790 1190.380 1487.110 1190.440 ;
        RECT 1486.790 1014.120 1487.110 1014.180 ;
        RECT 1489.550 1014.120 1489.870 1014.180 ;
        RECT 1486.790 1013.980 1489.870 1014.120 ;
        RECT 1486.790 1013.920 1487.110 1013.980 ;
        RECT 1489.550 1013.920 1489.870 1013.980 ;
        RECT 1489.550 1007.660 1489.870 1007.720 ;
        RECT 2087.090 1007.660 2087.410 1007.720 ;
        RECT 1489.550 1007.520 2087.410 1007.660 ;
        RECT 1489.550 1007.460 1489.870 1007.520 ;
        RECT 2087.090 1007.460 2087.410 1007.520 ;
        RECT 1489.550 544.920 1489.870 544.980 ;
        RECT 1518.070 544.920 1518.390 544.980 ;
        RECT 1528.190 544.920 1528.510 544.980 ;
        RECT 1538.770 544.920 1539.090 544.980 ;
        RECT 1489.550 544.780 1539.090 544.920 ;
        RECT 1489.550 544.720 1489.870 544.780 ;
        RECT 1518.070 544.720 1518.390 544.780 ;
        RECT 1528.190 544.720 1528.510 544.780 ;
        RECT 1538.770 544.720 1539.090 544.780 ;
        RECT 2090.310 544.920 2090.630 544.980 ;
        RECT 2121.130 544.920 2121.450 544.980 ;
        RECT 2139.070 544.920 2139.390 544.980 ;
        RECT 2090.310 544.780 2139.390 544.920 ;
        RECT 2090.310 544.720 2090.630 544.780 ;
        RECT 2121.130 544.720 2121.450 544.780 ;
        RECT 2139.070 544.720 2139.390 544.780 ;
        RECT 710.310 14.180 710.630 14.240 ;
        RECT 728.250 14.180 728.570 14.240 ;
        RECT 746.190 14.180 746.510 14.240 ;
        RECT 763.670 14.180 763.990 14.240 ;
        RECT 781.610 14.180 781.930 14.240 ;
        RECT 799.550 14.180 799.870 14.240 ;
        RECT 817.490 14.180 817.810 14.240 ;
        RECT 835.430 14.180 835.750 14.240 ;
        RECT 852.910 14.180 853.230 14.240 ;
        RECT 870.850 14.180 871.170 14.240 ;
        RECT 888.790 14.180 889.110 14.240 ;
        RECT 906.730 14.180 907.050 14.240 ;
        RECT 924.210 14.180 924.530 14.240 ;
        RECT 942.150 14.180 942.470 14.240 ;
        RECT 960.090 14.180 960.410 14.240 ;
        RECT 978.030 14.180 978.350 14.240 ;
        RECT 995.970 14.180 996.290 14.240 ;
        RECT 1013.450 14.180 1013.770 14.240 ;
        RECT 1031.390 14.180 1031.710 14.240 ;
        RECT 1049.330 14.180 1049.650 14.240 ;
        RECT 1067.270 14.180 1067.590 14.240 ;
        RECT 1085.210 14.180 1085.530 14.240 ;
        RECT 1102.690 14.180 1103.010 14.240 ;
        RECT 1120.630 14.180 1120.950 14.240 ;
        RECT 1138.570 14.180 1138.890 14.240 ;
        RECT 1156.510 14.180 1156.830 14.240 ;
        RECT 1173.990 14.180 1174.310 14.240 ;
        RECT 1191.930 14.180 1192.250 14.240 ;
        RECT 1209.870 14.180 1210.190 14.240 ;
        RECT 1227.810 14.180 1228.130 14.240 ;
        RECT 1245.750 14.180 1246.070 14.240 ;
        RECT 1263.230 14.180 1263.550 14.240 ;
        RECT 1281.170 14.180 1281.490 14.240 ;
        RECT 1299.110 14.180 1299.430 14.240 ;
        RECT 1317.050 14.180 1317.370 14.240 ;
        RECT 1334.990 14.180 1335.310 14.240 ;
        RECT 1352.470 14.180 1352.790 14.240 ;
        RECT 1370.410 14.180 1370.730 14.240 ;
        RECT 1388.350 14.180 1388.670 14.240 ;
        RECT 1406.290 14.180 1406.610 14.240 ;
        RECT 1423.770 14.180 1424.090 14.240 ;
        RECT 1441.710 14.180 1442.030 14.240 ;
        RECT 1459.650 14.180 1459.970 14.240 ;
        RECT 1477.590 14.180 1477.910 14.240 ;
        RECT 1495.530 14.180 1495.850 14.240 ;
        RECT 1513.010 14.180 1513.330 14.240 ;
        RECT 1528.190 14.180 1528.510 14.240 ;
        RECT 1530.950 14.180 1531.270 14.240 ;
        RECT 1548.890 14.180 1549.210 14.240 ;
        RECT 1566.830 14.180 1567.150 14.240 ;
        RECT 1584.770 14.180 1585.090 14.240 ;
        RECT 1602.250 14.180 1602.570 14.240 ;
        RECT 1620.190 14.180 1620.510 14.240 ;
        RECT 1638.130 14.180 1638.450 14.240 ;
        RECT 1656.070 14.180 1656.390 14.240 ;
        RECT 1673.550 14.180 1673.870 14.240 ;
        RECT 1691.490 14.180 1691.810 14.240 ;
        RECT 1709.430 14.180 1709.750 14.240 ;
        RECT 1727.370 14.180 1727.690 14.240 ;
        RECT 1745.310 14.180 1745.630 14.240 ;
        RECT 1762.790 14.180 1763.110 14.240 ;
        RECT 1780.730 14.180 1781.050 14.240 ;
        RECT 1798.670 14.180 1798.990 14.240 ;
        RECT 1816.610 14.180 1816.930 14.240 ;
        RECT 1834.550 14.180 1834.870 14.240 ;
        RECT 1852.030 14.180 1852.350 14.240 ;
        RECT 1869.970 14.180 1870.290 14.240 ;
        RECT 1887.910 14.180 1888.230 14.240 ;
        RECT 1905.850 14.180 1906.170 14.240 ;
        RECT 1923.330 14.180 1923.650 14.240 ;
        RECT 1941.270 14.180 1941.590 14.240 ;
        RECT 1959.210 14.180 1959.530 14.240 ;
        RECT 1977.150 14.180 1977.470 14.240 ;
        RECT 1995.090 14.180 1995.410 14.240 ;
        RECT 2012.570 14.180 2012.890 14.240 ;
        RECT 2030.510 14.180 2030.830 14.240 ;
        RECT 2048.450 14.180 2048.770 14.240 ;
        RECT 2066.390 14.180 2066.710 14.240 ;
        RECT 2084.330 14.180 2084.650 14.240 ;
        RECT 2101.810 14.180 2102.130 14.240 ;
        RECT 2119.750 14.180 2120.070 14.240 ;
        RECT 2137.690 14.180 2138.010 14.240 ;
        RECT 2155.630 14.180 2155.950 14.240 ;
        RECT 2173.110 14.180 2173.430 14.240 ;
        RECT 2191.050 14.180 2191.370 14.240 ;
        RECT 2208.990 14.180 2209.310 14.240 ;
        RECT 2226.930 14.180 2227.250 14.240 ;
        RECT 2244.870 14.180 2245.190 14.240 ;
        RECT 2262.350 14.180 2262.670 14.240 ;
        RECT 2280.290 14.180 2280.610 14.240 ;
        RECT 2298.230 14.180 2298.550 14.240 ;
        RECT 2316.170 14.180 2316.490 14.240 ;
        RECT 2334.110 14.180 2334.430 14.240 ;
        RECT 2351.590 14.180 2351.910 14.240 ;
        RECT 2369.530 14.180 2369.850 14.240 ;
        RECT 2387.470 14.180 2387.790 14.240 ;
        RECT 2405.410 14.180 2405.730 14.240 ;
        RECT 2422.890 14.180 2423.210 14.240 ;
        RECT 2440.830 14.180 2441.150 14.240 ;
        RECT 2458.770 14.180 2459.090 14.240 ;
        RECT 2476.710 14.180 2477.030 14.240 ;
        RECT 2494.650 14.180 2494.970 14.240 ;
        RECT 2512.130 14.180 2512.450 14.240 ;
        RECT 2530.070 14.180 2530.390 14.240 ;
        RECT 2548.010 14.180 2548.330 14.240 ;
        RECT 2565.950 14.180 2566.270 14.240 ;
        RECT 2583.890 14.180 2584.210 14.240 ;
        RECT 2601.370 14.180 2601.690 14.240 ;
        RECT 2619.310 14.180 2619.630 14.240 ;
        RECT 2637.250 14.180 2637.570 14.240 ;
        RECT 2655.190 14.180 2655.510 14.240 ;
        RECT 2672.670 14.180 2672.990 14.240 ;
        RECT 2690.610 14.180 2690.930 14.240 ;
        RECT 2708.550 14.180 2708.870 14.240 ;
        RECT 2726.490 14.180 2726.810 14.240 ;
        RECT 2744.430 14.180 2744.750 14.240 ;
        RECT 2761.910 14.180 2762.230 14.240 ;
        RECT 2779.850 14.180 2780.170 14.240 ;
        RECT 2797.790 14.180 2798.110 14.240 ;
        RECT 2815.730 14.180 2816.050 14.240 ;
        RECT 2833.670 14.180 2833.990 14.240 ;
        RECT 2851.150 14.180 2851.470 14.240 ;
        RECT 2869.090 14.180 2869.410 14.240 ;
        RECT 2887.030 14.180 2887.350 14.240 ;
        RECT 2904.970 14.180 2905.290 14.240 ;
        RECT 710.310 14.040 2905.290 14.180 ;
        RECT 710.310 13.980 710.630 14.040 ;
        RECT 728.250 13.980 728.570 14.040 ;
        RECT 746.190 13.980 746.510 14.040 ;
        RECT 763.670 13.980 763.990 14.040 ;
        RECT 781.610 13.980 781.930 14.040 ;
        RECT 799.550 13.980 799.870 14.040 ;
        RECT 817.490 13.980 817.810 14.040 ;
        RECT 835.430 13.980 835.750 14.040 ;
        RECT 852.910 13.980 853.230 14.040 ;
        RECT 870.850 13.980 871.170 14.040 ;
        RECT 888.790 13.980 889.110 14.040 ;
        RECT 906.730 13.980 907.050 14.040 ;
        RECT 924.210 13.980 924.530 14.040 ;
        RECT 942.150 13.980 942.470 14.040 ;
        RECT 960.090 13.980 960.410 14.040 ;
        RECT 978.030 13.980 978.350 14.040 ;
        RECT 995.970 13.980 996.290 14.040 ;
        RECT 1013.450 13.980 1013.770 14.040 ;
        RECT 1031.390 13.980 1031.710 14.040 ;
        RECT 1049.330 13.980 1049.650 14.040 ;
        RECT 1067.270 13.980 1067.590 14.040 ;
        RECT 1085.210 13.980 1085.530 14.040 ;
        RECT 1102.690 13.980 1103.010 14.040 ;
        RECT 1120.630 13.980 1120.950 14.040 ;
        RECT 1138.570 13.980 1138.890 14.040 ;
        RECT 1156.510 13.980 1156.830 14.040 ;
        RECT 1173.990 13.980 1174.310 14.040 ;
        RECT 1191.930 13.980 1192.250 14.040 ;
        RECT 1209.870 13.980 1210.190 14.040 ;
        RECT 1227.810 13.980 1228.130 14.040 ;
        RECT 1245.750 13.980 1246.070 14.040 ;
        RECT 1263.230 13.980 1263.550 14.040 ;
        RECT 1281.170 13.980 1281.490 14.040 ;
        RECT 1299.110 13.980 1299.430 14.040 ;
        RECT 1317.050 13.980 1317.370 14.040 ;
        RECT 1334.990 13.980 1335.310 14.040 ;
        RECT 1352.470 13.980 1352.790 14.040 ;
        RECT 1370.410 13.980 1370.730 14.040 ;
        RECT 1388.350 13.980 1388.670 14.040 ;
        RECT 1406.290 13.980 1406.610 14.040 ;
        RECT 1423.770 13.980 1424.090 14.040 ;
        RECT 1441.710 13.980 1442.030 14.040 ;
        RECT 1459.650 13.980 1459.970 14.040 ;
        RECT 1477.590 13.980 1477.910 14.040 ;
        RECT 1495.530 13.980 1495.850 14.040 ;
        RECT 1513.010 13.980 1513.330 14.040 ;
        RECT 1528.190 13.980 1528.510 14.040 ;
        RECT 1530.950 13.980 1531.270 14.040 ;
        RECT 1548.890 13.980 1549.210 14.040 ;
        RECT 1566.830 13.980 1567.150 14.040 ;
        RECT 1584.770 13.980 1585.090 14.040 ;
        RECT 1602.250 13.980 1602.570 14.040 ;
        RECT 1620.190 13.980 1620.510 14.040 ;
        RECT 1638.130 13.980 1638.450 14.040 ;
        RECT 1656.070 13.980 1656.390 14.040 ;
        RECT 1673.550 13.980 1673.870 14.040 ;
        RECT 1691.490 13.980 1691.810 14.040 ;
        RECT 1709.430 13.980 1709.750 14.040 ;
        RECT 1727.370 13.980 1727.690 14.040 ;
        RECT 1745.310 13.980 1745.630 14.040 ;
        RECT 1762.790 13.980 1763.110 14.040 ;
        RECT 1780.730 13.980 1781.050 14.040 ;
        RECT 1798.670 13.980 1798.990 14.040 ;
        RECT 1816.610 13.980 1816.930 14.040 ;
        RECT 1834.550 13.980 1834.870 14.040 ;
        RECT 1852.030 13.980 1852.350 14.040 ;
        RECT 1869.970 13.980 1870.290 14.040 ;
        RECT 1887.910 13.980 1888.230 14.040 ;
        RECT 1905.850 13.980 1906.170 14.040 ;
        RECT 1923.330 13.980 1923.650 14.040 ;
        RECT 1941.270 13.980 1941.590 14.040 ;
        RECT 1959.210 13.980 1959.530 14.040 ;
        RECT 1977.150 13.980 1977.470 14.040 ;
        RECT 1995.090 13.980 1995.410 14.040 ;
        RECT 2012.570 13.980 2012.890 14.040 ;
        RECT 2030.510 13.980 2030.830 14.040 ;
        RECT 2048.450 13.980 2048.770 14.040 ;
        RECT 2066.390 13.980 2066.710 14.040 ;
        RECT 2084.330 13.980 2084.650 14.040 ;
        RECT 2101.810 13.980 2102.130 14.040 ;
        RECT 2119.750 13.980 2120.070 14.040 ;
        RECT 2137.690 13.980 2138.010 14.040 ;
        RECT 2155.630 13.980 2155.950 14.040 ;
        RECT 2173.110 13.980 2173.430 14.040 ;
        RECT 2191.050 13.980 2191.370 14.040 ;
        RECT 2208.990 13.980 2209.310 14.040 ;
        RECT 2226.930 13.980 2227.250 14.040 ;
        RECT 2244.870 13.980 2245.190 14.040 ;
        RECT 2262.350 13.980 2262.670 14.040 ;
        RECT 2280.290 13.980 2280.610 14.040 ;
        RECT 2298.230 13.980 2298.550 14.040 ;
        RECT 2316.170 13.980 2316.490 14.040 ;
        RECT 2334.110 13.980 2334.430 14.040 ;
        RECT 2351.590 13.980 2351.910 14.040 ;
        RECT 2369.530 13.980 2369.850 14.040 ;
        RECT 2387.470 13.980 2387.790 14.040 ;
        RECT 2405.410 13.980 2405.730 14.040 ;
        RECT 2422.890 13.980 2423.210 14.040 ;
        RECT 2440.830 13.980 2441.150 14.040 ;
        RECT 2458.770 13.980 2459.090 14.040 ;
        RECT 2476.710 13.980 2477.030 14.040 ;
        RECT 2494.650 13.980 2494.970 14.040 ;
        RECT 2512.130 13.980 2512.450 14.040 ;
        RECT 2530.070 13.980 2530.390 14.040 ;
        RECT 2548.010 13.980 2548.330 14.040 ;
        RECT 2565.950 13.980 2566.270 14.040 ;
        RECT 2583.890 13.980 2584.210 14.040 ;
        RECT 2601.370 13.980 2601.690 14.040 ;
        RECT 2619.310 13.980 2619.630 14.040 ;
        RECT 2637.250 13.980 2637.570 14.040 ;
        RECT 2655.190 13.980 2655.510 14.040 ;
        RECT 2672.670 13.980 2672.990 14.040 ;
        RECT 2690.610 13.980 2690.930 14.040 ;
        RECT 2708.550 13.980 2708.870 14.040 ;
        RECT 2726.490 13.980 2726.810 14.040 ;
        RECT 2744.430 13.980 2744.750 14.040 ;
        RECT 2761.910 13.980 2762.230 14.040 ;
        RECT 2779.850 13.980 2780.170 14.040 ;
        RECT 2797.790 13.980 2798.110 14.040 ;
        RECT 2815.730 13.980 2816.050 14.040 ;
        RECT 2833.670 13.980 2833.990 14.040 ;
        RECT 2851.150 13.980 2851.470 14.040 ;
        RECT 2869.090 13.980 2869.410 14.040 ;
        RECT 2887.030 13.980 2887.350 14.040 ;
        RECT 2904.970 13.980 2905.290 14.040 ;
        RECT 692.370 2.960 692.690 3.020 ;
        RECT 710.310 2.960 710.630 3.020 ;
        RECT 692.370 2.820 710.630 2.960 ;
        RECT 692.370 2.760 692.690 2.820 ;
        RECT 710.310 2.760 710.630 2.820 ;
      LAYER via ;
        RECT 1406.780 1190.380 1407.040 1190.640 ;
        RECT 1486.820 1190.380 1487.080 1190.640 ;
        RECT 1486.820 1013.920 1487.080 1014.180 ;
        RECT 1489.580 1013.920 1489.840 1014.180 ;
        RECT 1489.580 1007.460 1489.840 1007.720 ;
        RECT 2087.120 1007.460 2087.380 1007.720 ;
        RECT 1489.580 544.720 1489.840 544.980 ;
        RECT 1518.100 544.720 1518.360 544.980 ;
        RECT 1528.220 544.720 1528.480 544.980 ;
        RECT 1538.800 544.720 1539.060 544.980 ;
        RECT 2090.340 544.720 2090.600 544.980 ;
        RECT 2121.160 544.720 2121.420 544.980 ;
        RECT 2139.100 544.720 2139.360 544.980 ;
        RECT 710.340 13.980 710.600 14.240 ;
        RECT 728.280 13.980 728.540 14.240 ;
        RECT 746.220 13.980 746.480 14.240 ;
        RECT 763.700 13.980 763.960 14.240 ;
        RECT 781.640 13.980 781.900 14.240 ;
        RECT 799.580 13.980 799.840 14.240 ;
        RECT 817.520 13.980 817.780 14.240 ;
        RECT 835.460 13.980 835.720 14.240 ;
        RECT 852.940 13.980 853.200 14.240 ;
        RECT 870.880 13.980 871.140 14.240 ;
        RECT 888.820 13.980 889.080 14.240 ;
        RECT 906.760 13.980 907.020 14.240 ;
        RECT 924.240 13.980 924.500 14.240 ;
        RECT 942.180 13.980 942.440 14.240 ;
        RECT 960.120 13.980 960.380 14.240 ;
        RECT 978.060 13.980 978.320 14.240 ;
        RECT 996.000 13.980 996.260 14.240 ;
        RECT 1013.480 13.980 1013.740 14.240 ;
        RECT 1031.420 13.980 1031.680 14.240 ;
        RECT 1049.360 13.980 1049.620 14.240 ;
        RECT 1067.300 13.980 1067.560 14.240 ;
        RECT 1085.240 13.980 1085.500 14.240 ;
        RECT 1102.720 13.980 1102.980 14.240 ;
        RECT 1120.660 13.980 1120.920 14.240 ;
        RECT 1138.600 13.980 1138.860 14.240 ;
        RECT 1156.540 13.980 1156.800 14.240 ;
        RECT 1174.020 13.980 1174.280 14.240 ;
        RECT 1191.960 13.980 1192.220 14.240 ;
        RECT 1209.900 13.980 1210.160 14.240 ;
        RECT 1227.840 13.980 1228.100 14.240 ;
        RECT 1245.780 13.980 1246.040 14.240 ;
        RECT 1263.260 13.980 1263.520 14.240 ;
        RECT 1281.200 13.980 1281.460 14.240 ;
        RECT 1299.140 13.980 1299.400 14.240 ;
        RECT 1317.080 13.980 1317.340 14.240 ;
        RECT 1335.020 13.980 1335.280 14.240 ;
        RECT 1352.500 13.980 1352.760 14.240 ;
        RECT 1370.440 13.980 1370.700 14.240 ;
        RECT 1388.380 13.980 1388.640 14.240 ;
        RECT 1406.320 13.980 1406.580 14.240 ;
        RECT 1423.800 13.980 1424.060 14.240 ;
        RECT 1441.740 13.980 1442.000 14.240 ;
        RECT 1459.680 13.980 1459.940 14.240 ;
        RECT 1477.620 13.980 1477.880 14.240 ;
        RECT 1495.560 13.980 1495.820 14.240 ;
        RECT 1513.040 13.980 1513.300 14.240 ;
        RECT 1528.220 13.980 1528.480 14.240 ;
        RECT 1530.980 13.980 1531.240 14.240 ;
        RECT 1548.920 13.980 1549.180 14.240 ;
        RECT 1566.860 13.980 1567.120 14.240 ;
        RECT 1584.800 13.980 1585.060 14.240 ;
        RECT 1602.280 13.980 1602.540 14.240 ;
        RECT 1620.220 13.980 1620.480 14.240 ;
        RECT 1638.160 13.980 1638.420 14.240 ;
        RECT 1656.100 13.980 1656.360 14.240 ;
        RECT 1673.580 13.980 1673.840 14.240 ;
        RECT 1691.520 13.980 1691.780 14.240 ;
        RECT 1709.460 13.980 1709.720 14.240 ;
        RECT 1727.400 13.980 1727.660 14.240 ;
        RECT 1745.340 13.980 1745.600 14.240 ;
        RECT 1762.820 13.980 1763.080 14.240 ;
        RECT 1780.760 13.980 1781.020 14.240 ;
        RECT 1798.700 13.980 1798.960 14.240 ;
        RECT 1816.640 13.980 1816.900 14.240 ;
        RECT 1834.580 13.980 1834.840 14.240 ;
        RECT 1852.060 13.980 1852.320 14.240 ;
        RECT 1870.000 13.980 1870.260 14.240 ;
        RECT 1887.940 13.980 1888.200 14.240 ;
        RECT 1905.880 13.980 1906.140 14.240 ;
        RECT 1923.360 13.980 1923.620 14.240 ;
        RECT 1941.300 13.980 1941.560 14.240 ;
        RECT 1959.240 13.980 1959.500 14.240 ;
        RECT 1977.180 13.980 1977.440 14.240 ;
        RECT 1995.120 13.980 1995.380 14.240 ;
        RECT 2012.600 13.980 2012.860 14.240 ;
        RECT 2030.540 13.980 2030.800 14.240 ;
        RECT 2048.480 13.980 2048.740 14.240 ;
        RECT 2066.420 13.980 2066.680 14.240 ;
        RECT 2084.360 13.980 2084.620 14.240 ;
        RECT 2101.840 13.980 2102.100 14.240 ;
        RECT 2119.780 13.980 2120.040 14.240 ;
        RECT 2137.720 13.980 2137.980 14.240 ;
        RECT 2155.660 13.980 2155.920 14.240 ;
        RECT 2173.140 13.980 2173.400 14.240 ;
        RECT 2191.080 13.980 2191.340 14.240 ;
        RECT 2209.020 13.980 2209.280 14.240 ;
        RECT 2226.960 13.980 2227.220 14.240 ;
        RECT 2244.900 13.980 2245.160 14.240 ;
        RECT 2262.380 13.980 2262.640 14.240 ;
        RECT 2280.320 13.980 2280.580 14.240 ;
        RECT 2298.260 13.980 2298.520 14.240 ;
        RECT 2316.200 13.980 2316.460 14.240 ;
        RECT 2334.140 13.980 2334.400 14.240 ;
        RECT 2351.620 13.980 2351.880 14.240 ;
        RECT 2369.560 13.980 2369.820 14.240 ;
        RECT 2387.500 13.980 2387.760 14.240 ;
        RECT 2405.440 13.980 2405.700 14.240 ;
        RECT 2422.920 13.980 2423.180 14.240 ;
        RECT 2440.860 13.980 2441.120 14.240 ;
        RECT 2458.800 13.980 2459.060 14.240 ;
        RECT 2476.740 13.980 2477.000 14.240 ;
        RECT 2494.680 13.980 2494.940 14.240 ;
        RECT 2512.160 13.980 2512.420 14.240 ;
        RECT 2530.100 13.980 2530.360 14.240 ;
        RECT 2548.040 13.980 2548.300 14.240 ;
        RECT 2565.980 13.980 2566.240 14.240 ;
        RECT 2583.920 13.980 2584.180 14.240 ;
        RECT 2601.400 13.980 2601.660 14.240 ;
        RECT 2619.340 13.980 2619.600 14.240 ;
        RECT 2637.280 13.980 2637.540 14.240 ;
        RECT 2655.220 13.980 2655.480 14.240 ;
        RECT 2672.700 13.980 2672.960 14.240 ;
        RECT 2690.640 13.980 2690.900 14.240 ;
        RECT 2708.580 13.980 2708.840 14.240 ;
        RECT 2726.520 13.980 2726.780 14.240 ;
        RECT 2744.460 13.980 2744.720 14.240 ;
        RECT 2761.940 13.980 2762.200 14.240 ;
        RECT 2779.880 13.980 2780.140 14.240 ;
        RECT 2797.820 13.980 2798.080 14.240 ;
        RECT 2815.760 13.980 2816.020 14.240 ;
        RECT 2833.700 13.980 2833.960 14.240 ;
        RECT 2851.180 13.980 2851.440 14.240 ;
        RECT 2869.120 13.980 2869.380 14.240 ;
        RECT 2887.060 13.980 2887.320 14.240 ;
        RECT 2905.000 13.980 2905.260 14.240 ;
        RECT 692.400 2.760 692.660 3.020 ;
        RECT 710.340 2.760 710.600 3.020 ;
      LAYER met2 ;
        RECT 1405.150 1200.610 1405.430 1204.000 ;
        RECT 1405.150 1200.470 1406.980 1200.610 ;
        RECT 1405.150 1200.000 1405.430 1200.470 ;
        RECT 1406.840 1190.670 1406.980 1200.470 ;
        RECT 1406.780 1190.350 1407.040 1190.670 ;
        RECT 1486.820 1190.350 1487.080 1190.670 ;
        RECT 1486.880 1014.210 1487.020 1190.350 ;
        RECT 1486.820 1013.890 1487.080 1014.210 ;
        RECT 1489.580 1013.890 1489.840 1014.210 ;
        RECT 1489.640 1007.750 1489.780 1013.890 ;
        RECT 1489.580 1007.430 1489.840 1007.750 ;
        RECT 2087.120 1007.430 2087.380 1007.750 ;
        RECT 1489.640 901.525 1489.780 1007.430 ;
        RECT 2087.180 902.885 2087.320 1007.430 ;
        RECT 2087.110 902.515 2087.390 902.885 ;
        RECT 1489.570 901.155 1489.850 901.525 ;
        RECT 1489.570 858.995 1489.850 859.365 ;
        RECT 1489.640 545.010 1489.780 858.995 ;
        RECT 2090.330 858.315 2090.610 858.685 ;
        RECT 1489.580 544.690 1489.840 545.010 ;
        RECT 1518.090 544.835 1518.370 545.205 ;
        RECT 1518.100 544.690 1518.360 544.835 ;
        RECT 1528.220 544.690 1528.480 545.010 ;
        RECT 1538.790 544.835 1539.070 545.205 ;
        RECT 2090.400 545.010 2090.540 858.315 ;
        RECT 1538.800 544.690 1539.060 544.835 ;
        RECT 2090.340 544.690 2090.600 545.010 ;
        RECT 2121.150 544.835 2121.430 545.205 ;
        RECT 2139.090 544.835 2139.370 545.205 ;
        RECT 2121.160 544.690 2121.420 544.835 ;
        RECT 2139.100 544.690 2139.360 544.835 ;
        RECT 1528.280 14.270 1528.420 544.690 ;
        RECT 710.340 13.950 710.600 14.270 ;
        RECT 728.280 13.950 728.540 14.270 ;
        RECT 746.220 13.950 746.480 14.270 ;
        RECT 763.700 13.950 763.960 14.270 ;
        RECT 781.640 13.950 781.900 14.270 ;
        RECT 799.580 13.950 799.840 14.270 ;
        RECT 817.520 13.950 817.780 14.270 ;
        RECT 835.460 13.950 835.720 14.270 ;
        RECT 852.940 13.950 853.200 14.270 ;
        RECT 870.880 13.950 871.140 14.270 ;
        RECT 888.820 13.950 889.080 14.270 ;
        RECT 906.760 13.950 907.020 14.270 ;
        RECT 924.240 13.950 924.500 14.270 ;
        RECT 942.180 13.950 942.440 14.270 ;
        RECT 960.120 13.950 960.380 14.270 ;
        RECT 978.060 13.950 978.320 14.270 ;
        RECT 996.000 13.950 996.260 14.270 ;
        RECT 1013.480 13.950 1013.740 14.270 ;
        RECT 1031.420 13.950 1031.680 14.270 ;
        RECT 1049.360 13.950 1049.620 14.270 ;
        RECT 1067.300 13.950 1067.560 14.270 ;
        RECT 1085.240 13.950 1085.500 14.270 ;
        RECT 1102.720 13.950 1102.980 14.270 ;
        RECT 1120.660 13.950 1120.920 14.270 ;
        RECT 1138.600 13.950 1138.860 14.270 ;
        RECT 1156.540 13.950 1156.800 14.270 ;
        RECT 1174.020 13.950 1174.280 14.270 ;
        RECT 1191.960 13.950 1192.220 14.270 ;
        RECT 1209.900 13.950 1210.160 14.270 ;
        RECT 1227.840 13.950 1228.100 14.270 ;
        RECT 1245.780 13.950 1246.040 14.270 ;
        RECT 1263.260 13.950 1263.520 14.270 ;
        RECT 1281.200 13.950 1281.460 14.270 ;
        RECT 1299.140 13.950 1299.400 14.270 ;
        RECT 1317.080 13.950 1317.340 14.270 ;
        RECT 1335.020 13.950 1335.280 14.270 ;
        RECT 1352.500 13.950 1352.760 14.270 ;
        RECT 1370.440 13.950 1370.700 14.270 ;
        RECT 1388.380 13.950 1388.640 14.270 ;
        RECT 1406.320 13.950 1406.580 14.270 ;
        RECT 1423.800 13.950 1424.060 14.270 ;
        RECT 1441.740 13.950 1442.000 14.270 ;
        RECT 1459.680 13.950 1459.940 14.270 ;
        RECT 1477.620 13.950 1477.880 14.270 ;
        RECT 1495.560 13.950 1495.820 14.270 ;
        RECT 1513.040 13.950 1513.300 14.270 ;
        RECT 1528.220 13.950 1528.480 14.270 ;
        RECT 1530.980 13.950 1531.240 14.270 ;
        RECT 1548.920 13.950 1549.180 14.270 ;
        RECT 1566.860 13.950 1567.120 14.270 ;
        RECT 1584.800 13.950 1585.060 14.270 ;
        RECT 1602.280 13.950 1602.540 14.270 ;
        RECT 1620.220 13.950 1620.480 14.270 ;
        RECT 1638.160 13.950 1638.420 14.270 ;
        RECT 1656.100 13.950 1656.360 14.270 ;
        RECT 1673.580 13.950 1673.840 14.270 ;
        RECT 1691.520 13.950 1691.780 14.270 ;
        RECT 1709.460 13.950 1709.720 14.270 ;
        RECT 1727.400 13.950 1727.660 14.270 ;
        RECT 1745.340 13.950 1745.600 14.270 ;
        RECT 1762.820 13.950 1763.080 14.270 ;
        RECT 1780.760 13.950 1781.020 14.270 ;
        RECT 1798.700 13.950 1798.960 14.270 ;
        RECT 1816.640 13.950 1816.900 14.270 ;
        RECT 1834.580 13.950 1834.840 14.270 ;
        RECT 1852.060 13.950 1852.320 14.270 ;
        RECT 1870.000 13.950 1870.260 14.270 ;
        RECT 1887.940 13.950 1888.200 14.270 ;
        RECT 1905.880 13.950 1906.140 14.270 ;
        RECT 1923.360 13.950 1923.620 14.270 ;
        RECT 1941.300 13.950 1941.560 14.270 ;
        RECT 1959.240 13.950 1959.500 14.270 ;
        RECT 1977.180 13.950 1977.440 14.270 ;
        RECT 1995.120 13.950 1995.380 14.270 ;
        RECT 2012.600 13.950 2012.860 14.270 ;
        RECT 2030.540 13.950 2030.800 14.270 ;
        RECT 2048.480 13.950 2048.740 14.270 ;
        RECT 2066.420 13.950 2066.680 14.270 ;
        RECT 2084.360 13.950 2084.620 14.270 ;
        RECT 2101.840 13.950 2102.100 14.270 ;
        RECT 2119.780 13.950 2120.040 14.270 ;
        RECT 2137.720 13.950 2137.980 14.270 ;
        RECT 2155.660 13.950 2155.920 14.270 ;
        RECT 2173.140 13.950 2173.400 14.270 ;
        RECT 2191.080 13.950 2191.340 14.270 ;
        RECT 2209.020 13.950 2209.280 14.270 ;
        RECT 2226.960 13.950 2227.220 14.270 ;
        RECT 2244.900 13.950 2245.160 14.270 ;
        RECT 2262.380 13.950 2262.640 14.270 ;
        RECT 2280.320 13.950 2280.580 14.270 ;
        RECT 2298.260 13.950 2298.520 14.270 ;
        RECT 2316.200 13.950 2316.460 14.270 ;
        RECT 2334.140 13.950 2334.400 14.270 ;
        RECT 2351.620 13.950 2351.880 14.270 ;
        RECT 2369.560 13.950 2369.820 14.270 ;
        RECT 2387.500 13.950 2387.760 14.270 ;
        RECT 2405.440 13.950 2405.700 14.270 ;
        RECT 2422.920 13.950 2423.180 14.270 ;
        RECT 2440.860 13.950 2441.120 14.270 ;
        RECT 2458.800 13.950 2459.060 14.270 ;
        RECT 2476.740 13.950 2477.000 14.270 ;
        RECT 2494.680 13.950 2494.940 14.270 ;
        RECT 2512.160 13.950 2512.420 14.270 ;
        RECT 2530.100 13.950 2530.360 14.270 ;
        RECT 2548.040 13.950 2548.300 14.270 ;
        RECT 2565.980 13.950 2566.240 14.270 ;
        RECT 2583.920 13.950 2584.180 14.270 ;
        RECT 2601.400 13.950 2601.660 14.270 ;
        RECT 2619.340 13.950 2619.600 14.270 ;
        RECT 2637.280 13.950 2637.540 14.270 ;
        RECT 2655.220 13.950 2655.480 14.270 ;
        RECT 2672.700 13.950 2672.960 14.270 ;
        RECT 2690.640 13.950 2690.900 14.270 ;
        RECT 2708.580 13.950 2708.840 14.270 ;
        RECT 2726.520 13.950 2726.780 14.270 ;
        RECT 2744.460 13.950 2744.720 14.270 ;
        RECT 2761.940 13.950 2762.200 14.270 ;
        RECT 2779.880 13.950 2780.140 14.270 ;
        RECT 2797.820 13.950 2798.080 14.270 ;
        RECT 2815.760 13.950 2816.020 14.270 ;
        RECT 2833.700 13.950 2833.960 14.270 ;
        RECT 2851.180 13.950 2851.440 14.270 ;
        RECT 2869.120 13.950 2869.380 14.270 ;
        RECT 2887.060 13.950 2887.320 14.270 ;
        RECT 2905.000 13.950 2905.260 14.270 ;
        RECT 710.400 3.050 710.540 13.950 ;
        RECT 692.400 2.730 692.660 3.050 ;
        RECT 710.340 2.730 710.600 3.050 ;
        RECT 692.460 2.400 692.600 2.730 ;
        RECT 710.400 2.400 710.540 2.730 ;
        RECT 728.340 2.400 728.480 13.950 ;
        RECT 746.280 2.400 746.420 13.950 ;
        RECT 763.760 2.400 763.900 13.950 ;
        RECT 781.700 2.400 781.840 13.950 ;
        RECT 799.640 2.400 799.780 13.950 ;
        RECT 817.580 2.400 817.720 13.950 ;
        RECT 835.520 2.400 835.660 13.950 ;
        RECT 853.000 2.400 853.140 13.950 ;
        RECT 870.940 2.400 871.080 13.950 ;
        RECT 888.880 2.400 889.020 13.950 ;
        RECT 906.820 2.400 906.960 13.950 ;
        RECT 924.300 2.400 924.440 13.950 ;
        RECT 942.240 2.400 942.380 13.950 ;
        RECT 960.180 2.400 960.320 13.950 ;
        RECT 978.120 2.400 978.260 13.950 ;
        RECT 996.060 2.400 996.200 13.950 ;
        RECT 1013.540 2.400 1013.680 13.950 ;
        RECT 1031.480 2.400 1031.620 13.950 ;
        RECT 1049.420 2.400 1049.560 13.950 ;
        RECT 1067.360 2.400 1067.500 13.950 ;
        RECT 1085.300 2.400 1085.440 13.950 ;
        RECT 1102.780 2.400 1102.920 13.950 ;
        RECT 1120.720 2.400 1120.860 13.950 ;
        RECT 1138.660 2.400 1138.800 13.950 ;
        RECT 1156.600 2.400 1156.740 13.950 ;
        RECT 1174.080 2.400 1174.220 13.950 ;
        RECT 1192.020 2.400 1192.160 13.950 ;
        RECT 1209.960 2.400 1210.100 13.950 ;
        RECT 1227.900 2.400 1228.040 13.950 ;
        RECT 1245.840 2.400 1245.980 13.950 ;
        RECT 1263.320 2.400 1263.460 13.950 ;
        RECT 1281.260 2.400 1281.400 13.950 ;
        RECT 1299.200 2.400 1299.340 13.950 ;
        RECT 1317.140 2.400 1317.280 13.950 ;
        RECT 1335.080 2.400 1335.220 13.950 ;
        RECT 1352.560 2.400 1352.700 13.950 ;
        RECT 1370.500 2.400 1370.640 13.950 ;
        RECT 1388.440 2.400 1388.580 13.950 ;
        RECT 1406.380 2.400 1406.520 13.950 ;
        RECT 1423.860 2.400 1424.000 13.950 ;
        RECT 1441.800 2.400 1441.940 13.950 ;
        RECT 1459.740 2.400 1459.880 13.950 ;
        RECT 1477.680 2.400 1477.820 13.950 ;
        RECT 1495.620 2.400 1495.760 13.950 ;
        RECT 1513.100 2.400 1513.240 13.950 ;
        RECT 1531.040 2.400 1531.180 13.950 ;
        RECT 1548.980 2.400 1549.120 13.950 ;
        RECT 1566.920 2.400 1567.060 13.950 ;
        RECT 1584.860 2.400 1585.000 13.950 ;
        RECT 1602.340 2.400 1602.480 13.950 ;
        RECT 1620.280 2.400 1620.420 13.950 ;
        RECT 1638.220 2.400 1638.360 13.950 ;
        RECT 1656.160 2.400 1656.300 13.950 ;
        RECT 1673.640 2.400 1673.780 13.950 ;
        RECT 1691.580 2.400 1691.720 13.950 ;
        RECT 1709.520 2.400 1709.660 13.950 ;
        RECT 1727.460 2.400 1727.600 13.950 ;
        RECT 1745.400 2.400 1745.540 13.950 ;
        RECT 1762.880 2.400 1763.020 13.950 ;
        RECT 1780.820 2.400 1780.960 13.950 ;
        RECT 1798.760 2.400 1798.900 13.950 ;
        RECT 1816.700 2.400 1816.840 13.950 ;
        RECT 1834.640 2.400 1834.780 13.950 ;
        RECT 1852.120 2.400 1852.260 13.950 ;
        RECT 1870.060 2.400 1870.200 13.950 ;
        RECT 1888.000 2.400 1888.140 13.950 ;
        RECT 1905.940 2.400 1906.080 13.950 ;
        RECT 1923.420 2.400 1923.560 13.950 ;
        RECT 1941.360 2.400 1941.500 13.950 ;
        RECT 1959.300 2.400 1959.440 13.950 ;
        RECT 1977.240 2.400 1977.380 13.950 ;
        RECT 1995.180 2.400 1995.320 13.950 ;
        RECT 2012.660 2.400 2012.800 13.950 ;
        RECT 2030.600 2.400 2030.740 13.950 ;
        RECT 2048.540 2.400 2048.680 13.950 ;
        RECT 2066.480 2.400 2066.620 13.950 ;
        RECT 2084.420 2.400 2084.560 13.950 ;
        RECT 2101.900 2.400 2102.040 13.950 ;
        RECT 2119.840 2.400 2119.980 13.950 ;
        RECT 2137.780 2.400 2137.920 13.950 ;
        RECT 2155.720 2.400 2155.860 13.950 ;
        RECT 2173.200 2.400 2173.340 13.950 ;
        RECT 2191.140 2.400 2191.280 13.950 ;
        RECT 2209.080 2.400 2209.220 13.950 ;
        RECT 2227.020 2.400 2227.160 13.950 ;
        RECT 2244.960 2.400 2245.100 13.950 ;
        RECT 2262.440 2.400 2262.580 13.950 ;
        RECT 2280.380 2.400 2280.520 13.950 ;
        RECT 2298.320 2.400 2298.460 13.950 ;
        RECT 2316.260 2.400 2316.400 13.950 ;
        RECT 2334.200 2.400 2334.340 13.950 ;
        RECT 2351.680 2.400 2351.820 13.950 ;
        RECT 2369.620 2.400 2369.760 13.950 ;
        RECT 2387.560 2.400 2387.700 13.950 ;
        RECT 2405.500 2.400 2405.640 13.950 ;
        RECT 2422.980 2.400 2423.120 13.950 ;
        RECT 2440.920 2.400 2441.060 13.950 ;
        RECT 2458.860 2.400 2459.000 13.950 ;
        RECT 2476.800 2.400 2476.940 13.950 ;
        RECT 2494.740 2.400 2494.880 13.950 ;
        RECT 2512.220 2.400 2512.360 13.950 ;
        RECT 2530.160 2.400 2530.300 13.950 ;
        RECT 2548.100 2.400 2548.240 13.950 ;
        RECT 2566.040 2.400 2566.180 13.950 ;
        RECT 2583.980 2.400 2584.120 13.950 ;
        RECT 2601.460 2.400 2601.600 13.950 ;
        RECT 2619.400 2.400 2619.540 13.950 ;
        RECT 2637.340 2.400 2637.480 13.950 ;
        RECT 2655.280 2.400 2655.420 13.950 ;
        RECT 2672.760 2.400 2672.900 13.950 ;
        RECT 2690.700 2.400 2690.840 13.950 ;
        RECT 2708.640 2.400 2708.780 13.950 ;
        RECT 2726.580 2.400 2726.720 13.950 ;
        RECT 2744.520 2.400 2744.660 13.950 ;
        RECT 2762.000 2.400 2762.140 13.950 ;
        RECT 2779.940 2.400 2780.080 13.950 ;
        RECT 2797.880 2.400 2798.020 13.950 ;
        RECT 2815.820 2.400 2815.960 13.950 ;
        RECT 2833.760 2.400 2833.900 13.950 ;
        RECT 2851.240 2.400 2851.380 13.950 ;
        RECT 2869.180 2.400 2869.320 13.950 ;
        RECT 2887.120 2.400 2887.260 13.950 ;
        RECT 2905.060 2.400 2905.200 13.950 ;
        RECT 692.250 -4.800 692.810 2.400 ;
        RECT 710.190 -4.800 710.750 2.400 ;
        RECT 728.130 -4.800 728.690 2.400 ;
        RECT 746.070 -4.800 746.630 2.400 ;
        RECT 763.550 -4.800 764.110 2.400 ;
        RECT 781.490 -4.800 782.050 2.400 ;
        RECT 799.430 -4.800 799.990 2.400 ;
        RECT 817.370 -4.800 817.930 2.400 ;
        RECT 835.310 -4.800 835.870 2.400 ;
        RECT 852.790 -4.800 853.350 2.400 ;
        RECT 870.730 -4.800 871.290 2.400 ;
        RECT 888.670 -4.800 889.230 2.400 ;
        RECT 906.610 -4.800 907.170 2.400 ;
        RECT 924.090 -4.800 924.650 2.400 ;
        RECT 942.030 -4.800 942.590 2.400 ;
        RECT 959.970 -4.800 960.530 2.400 ;
        RECT 977.910 -4.800 978.470 2.400 ;
        RECT 995.850 -4.800 996.410 2.400 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 2087.110 902.560 2087.390 902.840 ;
        RECT 1489.570 901.200 1489.850 901.480 ;
        RECT 1489.570 859.040 1489.850 859.320 ;
        RECT 2090.330 858.360 2090.610 858.640 ;
        RECT 1518.090 544.880 1518.370 545.160 ;
        RECT 1538.790 544.880 1539.070 545.160 ;
        RECT 2121.150 544.880 2121.430 545.160 ;
        RECT 2139.090 544.880 2139.370 545.160 ;
      LAYER met3 ;
        RECT 2087.085 902.850 2087.415 902.865 ;
        RECT 2087.085 902.550 2101.890 902.850 ;
        RECT 2087.085 902.535 2087.415 902.550 ;
        RECT 2101.590 901.745 2101.890 902.550 ;
        RECT 1489.545 901.490 1489.875 901.505 ;
        RECT 1500.000 901.490 1504.600 901.745 ;
        RECT 1489.545 901.445 1504.600 901.490 ;
        RECT 2100.000 901.445 2104.600 901.745 ;
        RECT 1489.545 901.190 1501.130 901.445 ;
        RECT 1489.545 901.175 1489.875 901.190 ;
        RECT 1500.830 896.105 1501.130 901.190 ;
        RECT 2101.590 896.105 2101.890 901.445 ;
        RECT 1500.000 895.805 1504.600 896.105 ;
        RECT 2100.000 895.805 2104.600 896.105 ;
        RECT 1500.830 887.605 1501.130 895.805 ;
        RECT 2101.590 887.605 2101.890 895.805 ;
        RECT 1500.000 887.305 1504.600 887.605 ;
        RECT 2100.000 887.305 2104.600 887.605 ;
        RECT 1500.830 881.965 1501.130 887.305 ;
        RECT 2101.590 881.965 2101.890 887.305 ;
        RECT 1500.000 881.665 1504.600 881.965 ;
        RECT 2100.000 881.665 2104.600 881.965 ;
        RECT 1500.830 873.465 1501.130 881.665 ;
        RECT 2101.590 873.465 2101.890 881.665 ;
        RECT 1500.000 873.165 1504.600 873.465 ;
        RECT 2100.000 873.165 2104.600 873.465 ;
        RECT 1500.830 867.825 1501.130 873.165 ;
        RECT 2101.590 867.825 2101.890 873.165 ;
        RECT 1500.000 867.525 1504.600 867.825 ;
        RECT 2100.000 867.525 2104.600 867.825 ;
        RECT 1489.545 859.330 1489.875 859.345 ;
        RECT 1489.545 859.325 1498.370 859.330 ;
        RECT 1500.830 859.325 1501.130 867.525 ;
        RECT 2101.590 859.325 2101.890 867.525 ;
        RECT 1489.545 859.030 1504.600 859.325 ;
        RECT 1489.545 859.015 1489.875 859.030 ;
        RECT 1498.070 859.025 1504.600 859.030 ;
        RECT 2100.000 859.025 2104.600 859.325 ;
        RECT 2090.305 858.650 2090.635 858.665 ;
        RECT 2100.670 858.650 2100.970 859.025 ;
        RECT 2090.305 858.350 2100.970 858.650 ;
        RECT 2090.305 858.335 2090.635 858.350 ;
        RECT 1518.065 545.180 1518.395 545.185 ;
        RECT 1518.065 545.170 1518.650 545.180 ;
        RECT 1538.765 545.170 1539.095 545.185 ;
        RECT 2121.125 545.180 2121.455 545.185 ;
        RECT 1540.350 545.170 1540.730 545.180 ;
        RECT 2120.870 545.170 2121.455 545.180 ;
        RECT 1518.065 544.870 1518.850 545.170 ;
        RECT 1538.765 544.870 1540.730 545.170 ;
        RECT 2120.670 544.870 2121.455 545.170 ;
        RECT 1518.065 544.860 1518.650 544.870 ;
        RECT 1518.065 544.855 1518.395 544.860 ;
        RECT 1538.765 544.855 1539.095 544.870 ;
        RECT 1540.350 544.860 1540.730 544.870 ;
        RECT 2120.870 544.860 2121.455 544.870 ;
        RECT 2121.125 544.855 2121.455 544.860 ;
        RECT 2139.065 545.170 2139.395 545.185 ;
        RECT 2140.190 545.170 2140.570 545.180 ;
        RECT 2139.065 544.870 2140.570 545.170 ;
        RECT 2139.065 544.855 2139.395 544.870 ;
        RECT 2140.190 544.860 2140.570 544.870 ;
      LAYER via3 ;
        RECT 1518.300 544.860 1518.620 545.180 ;
        RECT 1540.380 544.860 1540.700 545.180 ;
        RECT 2120.900 544.860 2121.220 545.180 ;
        RECT 2140.220 544.860 2140.540 545.180 ;
      LAYER met4 ;
        RECT 1518.315 550.950 1518.615 554.600 ;
        RECT 1543.290 550.950 1543.590 554.600 ;
        RECT 1518.310 550.000 1518.615 550.950 ;
        RECT 1540.390 550.650 1543.590 550.950 ;
        RECT 1518.310 545.185 1518.610 550.000 ;
        RECT 1540.390 545.185 1540.690 550.650 ;
        RECT 1543.290 550.000 1543.590 550.650 ;
        RECT 2118.315 550.950 2118.615 554.600 ;
        RECT 2143.290 550.950 2143.590 554.600 ;
        RECT 2118.315 550.650 2121.210 550.950 ;
        RECT 2118.315 550.000 2118.615 550.650 ;
        RECT 2120.910 545.185 2121.210 550.650 ;
        RECT 2140.230 550.650 2143.590 550.950 ;
        RECT 2140.230 545.185 2140.530 550.650 ;
        RECT 2143.290 550.000 2143.590 550.650 ;
        RECT 1518.295 544.855 1518.625 545.185 ;
        RECT 1540.375 544.855 1540.705 545.185 ;
        RECT 2120.895 544.855 2121.225 545.185 ;
        RECT 2140.215 544.855 2140.545 545.185 ;
    END
  END la_data_out[100]
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1881.480 3043.600 1884.050 3044.660 ;
        RECT 2481.480 3043.600 2484.050 3044.660 ;
        RECT 1502.430 561.575 1505.000 562.635 ;
        RECT 2102.430 561.575 2105.000 562.635 ;
      LAYER via3 ;
        RECT 1882.500 3043.620 1884.020 3044.630 ;
        RECT 2482.500 3043.620 2484.020 3044.630 ;
        RECT 1502.460 561.605 1503.980 562.615 ;
        RECT 2102.460 561.605 2103.980 562.615 ;
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 -9.320 367.020 3529.000 ;
        RECT 544.020 -9.320 547.020 3529.000 ;
        RECT 724.020 -9.320 727.020 3529.000 ;
        RECT 904.020 -9.320 907.020 3529.000 ;
        RECT 1084.020 -9.320 1087.020 3529.000 ;
        RECT 1264.020 -9.320 1267.020 3529.000 ;
        RECT 1444.020 2415.000 1447.020 3529.000 ;
        RECT 1624.020 3071.235 1627.020 3529.000 ;
        RECT 1804.020 3071.235 1807.020 3529.000 ;
        RECT 1882.470 2603.670 1884.070 3044.680 ;
        RECT 1624.020 2415.000 1627.020 2585.000 ;
        RECT 1804.020 2415.000 1807.020 2585.000 ;
        RECT 1984.020 2415.000 1987.020 3529.000 ;
        RECT 2164.020 3071.235 2167.020 3529.000 ;
        RECT 2344.020 3071.235 2347.020 3529.000 ;
        RECT 2482.470 2603.670 2484.070 3044.680 ;
        RECT 2164.020 2415.000 2167.020 2585.000 ;
        RECT 2344.020 2415.000 2347.020 2585.000 ;
        RECT 2524.020 2415.000 2527.020 3529.000 ;
        RECT 1421.040 1210.640 1422.640 2388.880 ;
        RECT 1444.020 -9.320 1447.020 1185.000 ;
        RECT 1624.020 1021.235 1627.020 1185.000 ;
        RECT 1804.020 1021.235 1807.020 1185.000 ;
        RECT 1502.410 561.555 1504.010 1002.565 ;
        RECT 1624.020 -9.320 1627.020 535.000 ;
        RECT 1804.020 -9.320 1807.020 535.000 ;
        RECT 1984.020 -9.320 1987.020 1185.000 ;
        RECT 2164.020 1021.235 2167.020 1185.000 ;
        RECT 2344.020 1021.235 2347.020 1185.000 ;
        RECT 2102.410 561.555 2104.010 1002.565 ;
        RECT 2164.020 -9.320 2167.020 535.000 ;
        RECT 2344.020 -9.320 2347.020 535.000 ;
        RECT 2524.020 -9.320 2527.020 1185.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1882.680 2891.090 1883.860 2892.270 ;
        RECT 1882.680 2889.490 1883.860 2890.670 ;
        RECT 1882.680 2711.090 1883.860 2712.270 ;
        RECT 1882.680 2709.490 1883.860 2710.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 2482.680 2891.090 2483.860 2892.270 ;
        RECT 2482.680 2889.490 2483.860 2890.670 ;
        RECT 2482.680 2711.090 2483.860 2712.270 ;
        RECT 2482.680 2709.490 2483.860 2710.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1421.250 2351.090 1422.430 2352.270 ;
        RECT 1421.250 2349.490 1422.430 2350.670 ;
        RECT 1421.250 2171.090 1422.430 2172.270 ;
        RECT 1421.250 2169.490 1422.430 2170.670 ;
        RECT 1421.250 1991.090 1422.430 1992.270 ;
        RECT 1421.250 1989.490 1422.430 1990.670 ;
        RECT 1421.250 1811.090 1422.430 1812.270 ;
        RECT 1421.250 1809.490 1422.430 1810.670 ;
        RECT 1421.250 1631.090 1422.430 1632.270 ;
        RECT 1421.250 1629.490 1422.430 1630.670 ;
        RECT 1421.250 1451.090 1422.430 1452.270 ;
        RECT 1421.250 1449.490 1422.430 1450.670 ;
        RECT 1421.250 1271.090 1422.430 1272.270 ;
        RECT 1421.250 1269.490 1422.430 1270.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1502.620 911.090 1503.800 912.270 ;
        RECT 1502.620 909.490 1503.800 910.670 ;
        RECT 1502.620 731.090 1503.800 732.270 ;
        RECT 1502.620 729.490 1503.800 730.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 2102.620 911.090 2103.800 912.270 ;
        RECT 2102.620 909.490 2103.800 910.670 ;
        RECT 2102.620 731.090 2103.800 732.270 ;
        RECT 2102.620 729.490 2103.800 730.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1882.470 2892.380 1884.070 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2482.470 2892.380 2484.070 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1882.470 2889.370 1884.070 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2482.470 2889.370 2484.070 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1882.470 2712.380 1884.070 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2482.470 2712.380 2484.070 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1882.470 2709.370 1884.070 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2482.470 2709.370 2484.070 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1421.040 2352.380 1422.640 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1421.040 2349.370 1422.640 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1421.040 2172.380 1422.640 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1421.040 2169.370 1422.640 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1421.040 1992.380 1422.640 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1421.040 1989.370 1422.640 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1421.040 1812.380 1422.640 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1421.040 1809.370 1422.640 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1421.040 1632.380 1422.640 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1421.040 1629.370 1422.640 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1421.040 1452.380 1422.640 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1421.040 1449.370 1422.640 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1421.040 1272.380 1422.640 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1421.040 1269.370 1422.640 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1502.410 912.380 1504.010 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2102.410 912.380 2104.010 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1502.410 909.370 1504.010 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2102.410 909.370 2104.010 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1502.410 732.380 1504.010 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2102.410 732.380 2104.010 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1502.410 729.370 1504.010 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2102.410 729.370 2104.010 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1881.040 3051.235 1886.300 3052.140 ;
        RECT 2481.040 3051.235 2486.300 3052.140 ;
        RECT 1881.480 3050.400 1886.300 3051.235 ;
        RECT 2481.480 3050.400 2486.300 3051.235 ;
        RECT 1500.180 555.000 1505.000 555.835 ;
        RECT 2100.180 555.000 2105.000 555.835 ;
        RECT 1500.180 554.095 1505.440 555.000 ;
        RECT 2100.180 554.095 2105.440 555.000 ;
      LAYER via3 ;
        RECT 1884.720 3050.440 1886.240 3052.050 ;
        RECT 2484.720 3050.440 2486.240 3052.050 ;
        RECT 1500.240 554.185 1501.760 555.795 ;
        RECT 2100.240 554.185 2101.760 555.795 ;
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 -9.320 457.020 3529.000 ;
        RECT 634.020 -9.320 637.020 3529.000 ;
        RECT 814.020 -9.320 817.020 3529.000 ;
        RECT 994.020 -9.320 997.020 3529.000 ;
        RECT 1174.020 -9.320 1177.020 3529.000 ;
        RECT 1354.020 -9.320 1357.020 3529.000 ;
        RECT 1534.020 3071.235 1537.020 3529.000 ;
        RECT 1714.020 3071.235 1717.020 3529.000 ;
        RECT 1894.020 3071.235 1897.020 3529.000 ;
        RECT 1884.690 2604.060 1886.310 3052.140 ;
        RECT 1534.020 2415.000 1537.020 2585.000 ;
        RECT 1714.020 2415.000 1717.020 2585.000 ;
        RECT 1894.020 2415.000 1897.020 2585.000 ;
        RECT 2074.020 2415.000 2077.020 3529.000 ;
        RECT 2254.020 3071.235 2257.020 3529.000 ;
        RECT 2434.020 3071.235 2437.020 3529.000 ;
        RECT 2484.690 2604.060 2486.310 3052.140 ;
        RECT 2254.020 2415.000 2257.020 2585.000 ;
        RECT 2434.020 2415.000 2437.020 2585.000 ;
        RECT 2614.020 2415.000 2617.020 3529.000 ;
        RECT 1497.840 1210.640 1499.440 2388.880 ;
        RECT 1534.020 1021.235 1537.020 1185.000 ;
        RECT 1714.020 1021.235 1717.020 1185.000 ;
        RECT 1894.020 1021.235 1897.020 1185.000 ;
        RECT 1500.170 554.095 1501.790 1002.175 ;
        RECT 1534.020 -9.320 1537.020 535.000 ;
        RECT 1714.020 -9.320 1717.020 535.000 ;
        RECT 1894.020 -9.320 1897.020 535.000 ;
        RECT 2074.020 -9.320 2077.020 1185.000 ;
        RECT 2254.020 1021.235 2257.020 1185.000 ;
        RECT 2434.020 1021.235 2437.020 1185.000 ;
        RECT 2100.170 554.095 2101.790 1002.175 ;
        RECT 2254.020 -9.320 2257.020 535.000 ;
        RECT 2434.020 -9.320 2437.020 535.000 ;
        RECT 2614.020 -9.320 2617.020 1185.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1884.910 2981.090 1886.090 2982.270 ;
        RECT 1884.910 2979.490 1886.090 2980.670 ;
        RECT 1884.910 2801.090 1886.090 2802.270 ;
        RECT 1884.910 2799.490 1886.090 2800.670 ;
        RECT 1884.910 2621.090 1886.090 2622.270 ;
        RECT 1884.910 2619.490 1886.090 2620.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 2484.910 2981.090 2486.090 2982.270 ;
        RECT 2484.910 2979.490 2486.090 2980.670 ;
        RECT 2484.910 2801.090 2486.090 2802.270 ;
        RECT 2484.910 2799.490 2486.090 2800.670 ;
        RECT 2484.910 2621.090 2486.090 2622.270 ;
        RECT 2484.910 2619.490 2486.090 2620.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1498.050 2261.090 1499.230 2262.270 ;
        RECT 1498.050 2259.490 1499.230 2260.670 ;
        RECT 1498.050 2081.090 1499.230 2082.270 ;
        RECT 1498.050 2079.490 1499.230 2080.670 ;
        RECT 1498.050 1901.090 1499.230 1902.270 ;
        RECT 1498.050 1899.490 1499.230 1900.670 ;
        RECT 1498.050 1721.090 1499.230 1722.270 ;
        RECT 1498.050 1719.490 1499.230 1720.670 ;
        RECT 1498.050 1541.090 1499.230 1542.270 ;
        RECT 1498.050 1539.490 1499.230 1540.670 ;
        RECT 1498.050 1361.090 1499.230 1362.270 ;
        RECT 1498.050 1359.490 1499.230 1360.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1500.390 821.090 1501.570 822.270 ;
        RECT 1500.390 819.490 1501.570 820.670 ;
        RECT 1500.390 641.090 1501.570 642.270 ;
        RECT 1500.390 639.490 1501.570 640.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2100.390 821.090 2101.570 822.270 ;
        RECT 2100.390 819.490 2101.570 820.670 ;
        RECT 2100.390 641.090 2101.570 642.270 ;
        RECT 2100.390 639.490 2101.570 640.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1884.690 2982.380 1886.310 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2484.690 2982.380 2486.310 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1884.690 2979.370 1886.310 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2484.690 2979.370 2486.310 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1884.690 2802.380 1886.310 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2484.690 2802.380 2486.310 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1884.690 2799.370 1886.310 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2484.690 2799.370 2486.310 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1884.690 2622.380 1886.310 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2484.690 2622.380 2486.310 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1884.690 2619.370 1886.310 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2484.690 2619.370 2486.310 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1497.840 2262.380 1499.440 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1497.840 2259.370 1499.440 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1497.840 2082.380 1499.440 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1497.840 2079.370 1499.440 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1497.840 1902.380 1499.440 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1497.840 1899.370 1499.440 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1497.840 1722.380 1499.440 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1497.840 1719.370 1499.440 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1497.840 1542.380 1499.440 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1497.840 1539.370 1499.440 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1497.840 1362.380 1499.440 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1497.840 1359.370 1499.440 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1500.170 822.380 1501.790 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2100.170 822.380 2101.790 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1500.170 819.370 1501.790 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2100.170 819.370 2101.790 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1500.170 642.380 1501.790 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2100.170 642.380 2101.790 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1500.170 639.370 1501.790 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2100.170 639.370 2101.790 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 382.020 -18.720 385.020 3538.400 ;
        RECT 562.020 -18.720 565.020 3538.400 ;
        RECT 742.020 -18.720 745.020 3538.400 ;
        RECT 922.020 -18.720 925.020 3538.400 ;
        RECT 1102.020 -18.720 1105.020 3538.400 ;
        RECT 1282.020 -18.720 1285.020 3538.400 ;
        RECT 1462.020 2415.000 1465.020 3538.400 ;
        RECT 1642.020 3071.235 1645.020 3538.400 ;
        RECT 1822.020 3071.235 1825.020 3538.400 ;
        RECT 1642.020 2415.000 1645.020 2585.000 ;
        RECT 1822.020 2415.000 1825.020 2585.000 ;
        RECT 2002.020 2415.000 2005.020 3538.400 ;
        RECT 2182.020 3071.235 2185.020 3538.400 ;
        RECT 2362.020 3071.235 2365.020 3538.400 ;
        RECT 2182.020 2415.000 2185.020 2585.000 ;
        RECT 2362.020 2415.000 2365.020 2585.000 ;
        RECT 2542.020 2415.000 2545.020 3538.400 ;
        RECT 1462.020 -18.720 1465.020 1185.000 ;
        RECT 1642.020 1021.235 1645.020 1185.000 ;
        RECT 1822.020 1021.235 1825.020 1185.000 ;
        RECT 1642.020 -18.720 1645.020 535.000 ;
        RECT 1822.020 -18.720 1825.020 535.000 ;
        RECT 2002.020 -18.720 2005.020 1185.000 ;
        RECT 2182.020 1021.235 2185.020 1185.000 ;
        RECT 2362.020 1021.235 2365.020 1185.000 ;
        RECT 2182.020 -18.720 2185.020 535.000 ;
        RECT 2362.020 -18.720 2365.020 535.000 ;
        RECT 2542.020 -18.720 2545.020 1185.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 292.020 -18.720 295.020 3538.400 ;
        RECT 472.020 -18.720 475.020 3538.400 ;
        RECT 652.020 -18.720 655.020 3538.400 ;
        RECT 832.020 -18.720 835.020 3538.400 ;
        RECT 1012.020 -18.720 1015.020 3538.400 ;
        RECT 1192.020 -18.720 1195.020 3538.400 ;
        RECT 1372.020 -18.720 1375.020 3538.400 ;
        RECT 1552.020 3071.235 1555.020 3538.400 ;
        RECT 1732.020 3071.235 1735.020 3538.400 ;
        RECT 1552.020 2415.000 1555.020 2585.000 ;
        RECT 1732.020 2415.000 1735.020 2585.000 ;
        RECT 1912.020 2415.000 1915.020 3538.400 ;
        RECT 2092.020 3071.235 2095.020 3538.400 ;
        RECT 2272.020 3071.235 2275.020 3538.400 ;
        RECT 2452.020 3071.235 2455.020 3538.400 ;
        RECT 2092.020 2415.000 2095.020 2585.000 ;
        RECT 2272.020 2415.000 2275.020 2585.000 ;
        RECT 2452.020 2415.000 2455.020 2585.000 ;
        RECT 1552.020 -18.720 1555.020 535.000 ;
        RECT 1732.020 -18.720 1735.020 535.000 ;
        RECT 1912.020 -18.720 1915.020 1185.000 ;
        RECT 2092.020 -18.720 2095.020 535.000 ;
        RECT 2272.020 -18.720 2275.020 535.000 ;
        RECT 2452.020 -18.720 2455.020 535.000 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 400.020 -28.120 403.020 3547.800 ;
        RECT 580.020 -28.120 583.020 3547.800 ;
        RECT 760.020 -28.120 763.020 3547.800 ;
        RECT 940.020 -28.120 943.020 3547.800 ;
        RECT 1120.020 -28.120 1123.020 3547.800 ;
        RECT 1300.020 -28.120 1303.020 3547.800 ;
        RECT 1480.020 2415.000 1483.020 3547.800 ;
        RECT 1660.020 3071.235 1663.020 3547.800 ;
        RECT 1840.020 3071.235 1843.020 3547.800 ;
        RECT 1660.020 2415.000 1663.020 2585.000 ;
        RECT 1840.020 2415.000 1843.020 2585.000 ;
        RECT 2020.020 2415.000 2023.020 3547.800 ;
        RECT 2200.020 3071.235 2203.020 3547.800 ;
        RECT 2380.020 3071.235 2383.020 3547.800 ;
        RECT 2200.020 2415.000 2203.020 2585.000 ;
        RECT 2380.020 2415.000 2383.020 2585.000 ;
        RECT 2560.020 2415.000 2563.020 3547.800 ;
        RECT 1480.020 -28.120 1483.020 1185.000 ;
        RECT 1660.020 1021.235 1663.020 1185.000 ;
        RECT 1840.020 1021.235 1843.020 1185.000 ;
        RECT 1660.020 -28.120 1663.020 535.000 ;
        RECT 1840.020 -28.120 1843.020 535.000 ;
        RECT 2020.020 -28.120 2023.020 1185.000 ;
        RECT 2200.020 1021.235 2203.020 1185.000 ;
        RECT 2380.020 1021.235 2383.020 1185.000 ;
        RECT 2200.020 -28.120 2203.020 535.000 ;
        RECT 2380.020 -28.120 2383.020 535.000 ;
        RECT 2560.020 -28.120 2563.020 1185.000 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 310.020 -28.120 313.020 3547.800 ;
        RECT 490.020 -28.120 493.020 3547.800 ;
        RECT 670.020 -28.120 673.020 3547.800 ;
        RECT 850.020 -28.120 853.020 3547.800 ;
        RECT 1030.020 -28.120 1033.020 3547.800 ;
        RECT 1210.020 -28.120 1213.020 3547.800 ;
        RECT 1390.020 2415.000 1393.020 3547.800 ;
        RECT 1570.020 3071.235 1573.020 3547.800 ;
        RECT 1750.020 3071.235 1753.020 3547.800 ;
        RECT 1570.020 2415.000 1573.020 2585.000 ;
        RECT 1750.020 2415.000 1753.020 2585.000 ;
        RECT 1930.020 2415.000 1933.020 3547.800 ;
        RECT 2110.020 3071.235 2113.020 3547.800 ;
        RECT 2290.020 3071.235 2293.020 3547.800 ;
        RECT 2470.020 3071.235 2473.020 3547.800 ;
        RECT 2110.020 2415.000 2113.020 2585.000 ;
        RECT 2290.020 2415.000 2293.020 2585.000 ;
        RECT 2470.020 2415.000 2473.020 2585.000 ;
        RECT 1390.020 -28.120 1393.020 1185.000 ;
        RECT 1570.020 1021.235 1573.020 1185.000 ;
        RECT 1750.020 1021.235 1753.020 1185.000 ;
        RECT 1570.020 -28.120 1573.020 535.000 ;
        RECT 1750.020 -28.120 1753.020 535.000 ;
        RECT 1930.020 -28.120 1933.020 1185.000 ;
        RECT 2110.020 1021.235 2113.020 1185.000 ;
        RECT 2290.020 1021.235 2293.020 1185.000 ;
        RECT 2470.020 1021.235 2473.020 1185.000 ;
        RECT 2110.020 -28.120 2113.020 535.000 ;
        RECT 2290.020 -28.120 2293.020 535.000 ;
        RECT 2470.020 -28.120 2473.020 535.000 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 418.020 -37.520 421.020 3557.200 ;
        RECT 598.020 -37.520 601.020 3557.200 ;
        RECT 778.020 -37.520 781.020 3557.200 ;
        RECT 958.020 -37.520 961.020 3557.200 ;
        RECT 1138.020 -37.520 1141.020 3557.200 ;
        RECT 1318.020 -37.520 1321.020 3557.200 ;
        RECT 1498.020 3071.235 1501.020 3557.200 ;
        RECT 1678.020 3071.235 1681.020 3557.200 ;
        RECT 1858.020 3071.235 1861.020 3557.200 ;
        RECT 2038.020 2415.000 2041.020 3557.200 ;
        RECT 2218.020 3071.235 2221.020 3557.200 ;
        RECT 2398.020 3071.235 2401.020 3557.200 ;
        RECT 2578.020 2415.000 2581.020 3557.200 ;
        RECT 1498.020 1021.235 1501.020 1185.000 ;
        RECT 1678.020 1021.235 1681.020 1185.000 ;
        RECT 1858.020 1021.235 1861.020 1185.000 ;
        RECT 1498.020 -37.520 1501.020 535.000 ;
        RECT 1678.020 -37.520 1681.020 535.000 ;
        RECT 1858.020 -37.520 1861.020 535.000 ;
        RECT 2038.020 -37.520 2041.020 1185.000 ;
        RECT 2218.020 1021.235 2221.020 1185.000 ;
        RECT 2398.020 1021.235 2401.020 1185.000 ;
        RECT 2218.020 -37.520 2221.020 535.000 ;
        RECT 2398.020 -37.520 2401.020 535.000 ;
        RECT 2578.020 -37.520 2581.020 1185.000 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 328.020 -37.520 331.020 3557.200 ;
        RECT 508.020 -37.520 511.020 3557.200 ;
        RECT 688.020 -37.520 691.020 3557.200 ;
        RECT 868.020 -37.520 871.020 3557.200 ;
        RECT 1048.020 -37.520 1051.020 3557.200 ;
        RECT 1228.020 -37.520 1231.020 3557.200 ;
        RECT 1408.020 2415.000 1411.020 3557.200 ;
        RECT 1588.020 3071.235 1591.020 3557.200 ;
        RECT 1768.020 3071.235 1771.020 3557.200 ;
        RECT 1588.020 2415.000 1591.020 2585.000 ;
        RECT 1768.020 2415.000 1771.020 2585.000 ;
        RECT 1948.020 2415.000 1951.020 3557.200 ;
        RECT 2128.020 3071.235 2131.020 3557.200 ;
        RECT 2308.020 3071.235 2311.020 3557.200 ;
        RECT 2488.020 3071.235 2491.020 3557.200 ;
        RECT 2128.020 2415.000 2131.020 2585.000 ;
        RECT 2308.020 2415.000 2311.020 2585.000 ;
        RECT 2488.020 2415.000 2491.020 2585.000 ;
        RECT 1408.020 -37.520 1411.020 1185.000 ;
        RECT 1588.020 1021.235 1591.020 1185.000 ;
        RECT 1768.020 1021.235 1771.020 1185.000 ;
        RECT 1588.020 -37.520 1591.020 535.000 ;
        RECT 1768.020 -37.520 1771.020 535.000 ;
        RECT 1948.020 -37.520 1951.020 1185.000 ;
        RECT 2128.020 1021.235 2131.020 1185.000 ;
        RECT 2308.020 1021.235 2311.020 1185.000 ;
        RECT 2488.020 1021.235 2491.020 1185.000 ;
        RECT 2128.020 -37.520 2131.020 535.000 ;
        RECT 2308.020 -37.520 2311.020 535.000 ;
        RECT 2488.020 -37.520 2491.020 535.000 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
        RECT 1405.520 1210.795 2594.935 2388.725 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met1 ;
        RECT 2442.670 3067.040 2442.990 3067.100 ;
        RECT 2469.810 3067.040 2470.130 3067.100 ;
        RECT 2442.670 3066.900 2470.130 3067.040 ;
        RECT 2442.670 3066.840 2442.990 3066.900 ;
        RECT 2469.810 3066.840 2470.130 3066.900 ;
        RECT 1868.130 3063.980 1868.450 3064.040 ;
        RECT 1898.030 3063.980 1898.350 3064.040 ;
        RECT 2442.670 3063.980 2442.990 3064.040 ;
        RECT 1868.130 3063.840 2442.990 3063.980 ;
        RECT 1868.130 3063.780 1868.450 3063.840 ;
        RECT 1898.030 3063.780 1898.350 3063.840 ;
        RECT 2442.670 3063.780 2442.990 3063.840 ;
        RECT 2469.810 3063.980 2470.130 3064.040 ;
        RECT 2497.870 3063.980 2498.190 3064.040 ;
        RECT 2469.810 3063.840 2498.190 3063.980 ;
        RECT 2469.810 3063.780 2470.130 3063.840 ;
        RECT 2497.870 3063.780 2498.190 3063.840 ;
        RECT 1899.870 3052.080 1900.190 3052.140 ;
        RECT 2482.230 3052.080 2482.550 3052.140 ;
        RECT 1899.870 3051.940 2482.550 3052.080 ;
        RECT 1899.870 3051.880 1900.190 3051.940 ;
        RECT 2482.230 3051.880 2482.550 3051.940 ;
      LAYER met1 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
      LAYER met1 ;
        RECT 2048.910 2698.140 2049.230 2698.200 ;
        RECT 2083.870 2698.140 2084.190 2698.200 ;
        RECT 2048.910 2698.000 2084.190 2698.140 ;
        RECT 2048.910 2697.940 2049.230 2698.000 ;
        RECT 2083.870 2697.940 2084.190 2698.000 ;
      LAYER met1 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
      LAYER met1 ;
        RECT 1486.330 2604.640 1486.650 2604.700 ;
        RECT 2090.310 2604.640 2090.630 2604.700 ;
        RECT 1486.330 2604.500 2090.630 2604.640 ;
        RECT 1486.330 2604.440 1486.650 2604.500 ;
        RECT 2090.310 2604.440 2090.630 2604.500 ;
        RECT 1614.670 2594.440 1614.990 2594.500 ;
        RECT 1661.590 2594.440 1661.910 2594.500 ;
        RECT 1614.670 2594.300 1661.910 2594.440 ;
        RECT 1614.670 2594.240 1614.990 2594.300 ;
        RECT 1661.590 2594.240 1661.910 2594.300 ;
        RECT 1537.850 2594.100 1538.170 2594.160 ;
        RECT 1621.570 2594.100 1621.890 2594.160 ;
        RECT 1537.850 2593.960 1621.890 2594.100 ;
        RECT 1537.850 2593.900 1538.170 2593.960 ;
        RECT 1621.570 2593.900 1621.890 2593.960 ;
        RECT 1656.070 2594.100 1656.390 2594.160 ;
        RECT 1702.530 2594.100 1702.850 2594.160 ;
        RECT 1656.070 2593.960 1702.850 2594.100 ;
        RECT 1656.070 2593.900 1656.390 2593.960 ;
        RECT 1702.530 2593.900 1702.850 2593.960 ;
        RECT 1586.610 2593.760 1586.930 2593.820 ;
        RECT 1626.630 2593.760 1626.950 2593.820 ;
        RECT 1669.870 2593.760 1670.190 2593.820 ;
        RECT 1586.610 2593.620 1670.190 2593.760 ;
        RECT 1586.610 2593.560 1586.930 2593.620 ;
        RECT 1626.630 2593.560 1626.950 2593.620 ;
        RECT 1669.870 2593.560 1670.190 2593.620 ;
        RECT 1690.570 2593.760 1690.890 2593.820 ;
        RECT 1738.410 2593.760 1738.730 2593.820 ;
        RECT 1690.570 2593.620 1738.730 2593.760 ;
        RECT 1690.570 2593.560 1690.890 2593.620 ;
        RECT 1738.410 2593.560 1738.730 2593.620 ;
        RECT 2256.370 2593.760 2256.690 2593.820 ;
        RECT 2297.770 2593.760 2298.090 2593.820 ;
        RECT 2256.370 2593.620 2298.090 2593.760 ;
        RECT 2256.370 2593.560 2256.690 2593.620 ;
        RECT 2297.770 2593.560 2298.090 2593.620 ;
        RECT 1598.570 2593.420 1598.890 2593.480 ;
        RECT 1644.570 2593.420 1644.890 2593.480 ;
        RECT 1598.570 2593.280 1644.890 2593.420 ;
        RECT 1598.570 2593.220 1598.890 2593.280 ;
        RECT 1644.570 2593.220 1644.890 2593.280 ;
        RECT 1651.010 2593.420 1651.330 2593.480 ;
        RECT 1697.930 2593.420 1698.250 2593.480 ;
        RECT 1743.930 2593.420 1744.250 2593.480 ;
        RECT 1651.010 2593.280 1744.250 2593.420 ;
        RECT 1651.010 2593.220 1651.330 2593.280 ;
        RECT 1697.930 2593.220 1698.250 2593.280 ;
        RECT 1743.930 2593.220 1744.250 2593.280 ;
        RECT 2215.890 2593.420 2216.210 2593.480 ;
        RECT 2262.810 2593.420 2263.130 2593.480 ;
        RECT 2305.130 2593.420 2305.450 2593.480 ;
        RECT 2215.890 2593.280 2305.450 2593.420 ;
        RECT 2215.890 2593.220 2216.210 2593.280 ;
        RECT 2262.810 2593.220 2263.130 2593.280 ;
        RECT 2305.130 2593.220 2305.450 2593.280 ;
        RECT 1476.210 2593.080 1476.530 2593.140 ;
        RECT 1587.070 2593.080 1587.390 2593.140 ;
        RECT 1476.210 2592.940 1587.390 2593.080 ;
        RECT 1476.210 2592.880 1476.530 2592.940 ;
        RECT 1587.070 2592.880 1587.390 2592.940 ;
        RECT 1604.090 2593.080 1604.410 2593.140 ;
        RECT 1651.100 2593.080 1651.240 2593.220 ;
        RECT 1604.090 2592.940 1651.240 2593.080 ;
        RECT 1661.590 2593.080 1661.910 2593.140 ;
        RECT 1707.590 2593.080 1707.910 2593.140 ;
        RECT 1732.890 2593.080 1733.210 2593.140 ;
        RECT 2208.070 2593.080 2208.390 2593.140 ;
        RECT 1661.590 2592.940 1707.910 2593.080 ;
        RECT 1604.090 2592.880 1604.410 2592.940 ;
        RECT 1661.590 2592.880 1661.910 2592.940 ;
        RECT 1707.590 2592.880 1707.910 2592.940 ;
        RECT 1708.140 2592.940 2208.390 2593.080 ;
        RECT 1569.590 2592.740 1569.910 2592.800 ;
        RECT 1591.210 2592.740 1591.530 2592.800 ;
        RECT 1639.050 2592.740 1639.370 2592.800 ;
        RECT 1685.050 2592.740 1685.370 2592.800 ;
        RECT 1569.590 2592.600 1590.980 2592.740 ;
        RECT 1569.590 2592.540 1569.910 2592.600 ;
        RECT 1573.730 2592.400 1574.050 2592.460 ;
        RECT 1590.840 2592.400 1590.980 2592.600 ;
        RECT 1591.210 2592.600 1685.370 2592.740 ;
        RECT 1591.210 2592.540 1591.530 2592.600 ;
        RECT 1639.050 2592.540 1639.370 2592.600 ;
        RECT 1685.050 2592.540 1685.370 2592.600 ;
        RECT 1686.430 2592.740 1686.750 2592.800 ;
        RECT 1708.140 2592.740 1708.280 2592.940 ;
        RECT 1732.890 2592.880 1733.210 2592.940 ;
        RECT 2208.070 2592.880 2208.390 2592.940 ;
        RECT 2220.490 2593.080 2220.810 2593.140 ;
        RECT 2268.330 2593.080 2268.650 2593.140 ;
        RECT 2311.570 2593.080 2311.890 2593.140 ;
        RECT 2220.490 2592.940 2311.890 2593.080 ;
        RECT 2220.490 2592.880 2220.810 2592.940 ;
        RECT 2268.330 2592.880 2268.650 2592.940 ;
        RECT 2311.570 2592.880 2311.890 2592.940 ;
        RECT 1686.430 2592.600 1708.280 2592.740 ;
        RECT 1738.410 2592.740 1738.730 2592.800 ;
        RECT 2214.970 2592.740 2215.290 2592.800 ;
        RECT 1738.410 2592.600 2215.290 2592.740 ;
        RECT 1686.430 2592.540 1686.750 2592.600 ;
        RECT 1738.410 2592.540 1738.730 2592.600 ;
        RECT 2214.970 2592.540 2215.290 2592.600 ;
        RECT 2243.950 2592.740 2244.270 2592.800 ;
        RECT 2291.790 2592.740 2292.110 2592.800 ;
        RECT 2332.270 2592.740 2332.590 2592.800 ;
        RECT 2243.950 2592.600 2332.590 2592.740 ;
        RECT 2243.950 2592.540 2244.270 2592.600 ;
        RECT 2291.790 2592.540 2292.110 2592.600 ;
        RECT 2332.270 2592.540 2332.590 2592.600 ;
        RECT 1614.670 2592.400 1614.990 2592.460 ;
        RECT 1573.730 2592.260 1590.520 2592.400 ;
        RECT 1590.840 2592.260 1614.990 2592.400 ;
        RECT 1573.730 2592.200 1574.050 2592.260 ;
        RECT 1462.410 2592.060 1462.730 2592.120 ;
        RECT 1581.090 2592.060 1581.410 2592.120 ;
        RECT 1462.410 2591.920 1581.410 2592.060 ;
        RECT 1462.410 2591.860 1462.730 2591.920 ;
        RECT 1581.090 2591.860 1581.410 2591.920 ;
        RECT 1448.610 2591.720 1448.930 2591.780 ;
        RECT 1573.270 2591.720 1573.590 2591.780 ;
        RECT 1448.610 2591.580 1573.590 2591.720 ;
        RECT 1590.380 2591.720 1590.520 2592.260 ;
        RECT 1614.670 2592.200 1614.990 2592.260 ;
        RECT 1630.770 2592.400 1631.090 2592.460 ;
        RECT 1633.530 2592.400 1633.850 2592.460 ;
        RECT 1679.530 2592.400 1679.850 2592.460 ;
        RECT 1725.530 2592.400 1725.850 2592.460 ;
        RECT 1731.510 2592.400 1731.830 2592.460 ;
        RECT 1630.770 2592.260 1731.830 2592.400 ;
        RECT 1630.770 2592.200 1631.090 2592.260 ;
        RECT 1633.530 2592.200 1633.850 2592.260 ;
        RECT 1679.530 2592.200 1679.850 2592.260 ;
        RECT 1725.530 2592.200 1725.850 2592.260 ;
        RECT 1731.510 2592.200 1731.830 2592.260 ;
        RECT 1743.930 2592.400 1744.250 2592.460 ;
        RECT 2228.770 2592.400 2229.090 2592.460 ;
        RECT 1743.930 2592.260 2229.090 2592.400 ;
        RECT 1743.930 2592.200 1744.250 2592.260 ;
        RECT 2228.770 2592.200 2229.090 2592.260 ;
        RECT 2249.470 2592.400 2249.790 2592.460 ;
        RECT 2249.470 2592.260 2286.040 2592.400 ;
        RECT 2249.470 2592.200 2249.790 2592.260 ;
        RECT 1644.570 2592.060 1644.890 2592.120 ;
        RECT 1690.570 2592.060 1690.890 2592.120 ;
        RECT 1644.570 2591.920 1690.890 2592.060 ;
        RECT 1644.570 2591.860 1644.890 2591.920 ;
        RECT 1690.570 2591.860 1690.890 2591.920 ;
        RECT 1993.250 2592.060 1993.570 2592.120 ;
        RECT 2152.870 2592.060 2153.190 2592.120 ;
        RECT 1993.250 2591.920 2153.190 2592.060 ;
        RECT 1993.250 2591.860 1993.570 2591.920 ;
        RECT 2152.870 2591.860 2153.190 2591.920 ;
        RECT 2235.670 2592.060 2235.990 2592.120 ;
        RECT 2285.350 2592.060 2285.670 2592.120 ;
        RECT 2235.670 2591.920 2285.670 2592.060 ;
        RECT 2285.900 2592.060 2286.040 2592.260 ;
        RECT 2297.770 2592.060 2298.090 2592.120 ;
        RECT 2339.170 2592.060 2339.490 2592.120 ;
        RECT 2285.900 2591.920 2339.490 2592.060 ;
        RECT 2235.670 2591.860 2235.990 2591.920 ;
        RECT 2285.350 2591.860 2285.670 2591.920 ;
        RECT 2297.770 2591.860 2298.090 2591.920 ;
        RECT 2339.170 2591.860 2339.490 2591.920 ;
        RECT 1621.570 2591.720 1621.890 2591.780 ;
        RECT 1667.110 2591.720 1667.430 2591.780 ;
        RECT 1713.110 2591.720 1713.430 2591.780 ;
        RECT 1590.380 2591.580 1713.430 2591.720 ;
        RECT 1448.610 2591.520 1448.930 2591.580 ;
        RECT 1573.270 2591.520 1573.590 2591.580 ;
        RECT 1621.570 2591.520 1621.890 2591.580 ;
        RECT 1667.110 2591.520 1667.430 2591.580 ;
        RECT 1713.110 2591.520 1713.430 2591.580 ;
        RECT 1979.910 2591.720 1980.230 2591.780 ;
        RECT 2146.430 2591.720 2146.750 2591.780 ;
        RECT 1979.910 2591.580 2146.750 2591.720 ;
        RECT 1979.910 2591.520 1980.230 2591.580 ;
        RECT 2146.430 2591.520 2146.750 2591.580 ;
        RECT 2232.910 2591.720 2233.230 2591.780 ;
        RECT 2280.290 2591.720 2280.610 2591.780 ;
        RECT 2232.910 2591.580 2280.610 2591.720 ;
        RECT 2285.440 2591.720 2285.580 2591.860 ;
        RECT 2332.270 2591.720 2332.590 2591.780 ;
        RECT 2285.440 2591.580 2332.590 2591.720 ;
        RECT 2232.910 2591.520 2233.230 2591.580 ;
        RECT 2280.290 2591.520 2280.610 2591.580 ;
        RECT 2332.270 2591.520 2332.590 2591.580 ;
        RECT 1565.450 2591.380 1565.770 2591.440 ;
        RECT 1608.230 2591.380 1608.550 2591.440 ;
        RECT 1656.070 2591.380 1656.390 2591.440 ;
        RECT 1565.450 2591.240 1656.390 2591.380 ;
        RECT 1565.450 2591.180 1565.770 2591.240 ;
        RECT 1608.230 2591.180 1608.550 2591.240 ;
        RECT 1656.070 2591.180 1656.390 2591.240 ;
        RECT 1669.870 2591.380 1670.190 2591.440 ;
        RECT 1718.170 2591.380 1718.490 2591.440 ;
        RECT 1669.870 2591.240 1718.490 2591.380 ;
        RECT 1669.870 2591.180 1670.190 2591.240 ;
        RECT 1718.170 2591.180 1718.490 2591.240 ;
        RECT 1966.110 2591.380 1966.430 2591.440 ;
        RECT 2145.970 2591.380 2146.290 2591.440 ;
        RECT 1966.110 2591.240 2146.290 2591.380 ;
        RECT 1966.110 2591.180 1966.430 2591.240 ;
        RECT 2145.970 2591.180 2146.290 2591.240 ;
        RECT 2276.150 2591.380 2276.470 2591.440 ;
        RECT 2318.470 2591.380 2318.790 2591.440 ;
        RECT 2276.150 2591.240 2318.790 2591.380 ;
        RECT 2276.150 2591.180 2276.470 2591.240 ;
        RECT 2318.470 2591.180 2318.790 2591.240 ;
        RECT 2214.510 2591.040 2214.830 2591.100 ;
        RECT 2256.370 2591.040 2256.690 2591.100 ;
        RECT 2214.510 2590.900 2256.690 2591.040 ;
        RECT 2214.510 2590.840 2214.830 2590.900 ;
        RECT 2256.370 2590.840 2256.690 2590.900 ;
        RECT 2280.290 2591.040 2280.610 2591.100 ;
        RECT 2325.370 2591.040 2325.690 2591.100 ;
        RECT 2280.290 2590.900 2325.690 2591.040 ;
        RECT 2280.290 2590.840 2280.610 2590.900 ;
        RECT 2325.370 2590.840 2325.690 2590.900 ;
        RECT 1517.610 2590.700 1517.930 2590.760 ;
        RECT 1607.770 2590.700 1608.090 2590.760 ;
        RECT 1517.610 2590.560 1608.090 2590.700 ;
        RECT 1517.610 2590.500 1517.930 2590.560 ;
        RECT 1607.770 2590.500 1608.090 2590.560 ;
        RECT 1959.210 2590.700 1959.530 2590.760 ;
        RECT 2126.650 2590.700 2126.970 2590.760 ;
        RECT 1959.210 2590.560 2126.970 2590.700 ;
        RECT 1959.210 2590.500 1959.530 2590.560 ;
        RECT 2126.650 2590.500 2126.970 2590.560 ;
        RECT 1531.410 2590.360 1531.730 2590.420 ;
        RECT 1614.670 2590.360 1614.990 2590.420 ;
        RECT 1531.410 2590.220 1614.990 2590.360 ;
        RECT 1531.410 2590.160 1531.730 2590.220 ;
        RECT 1614.670 2590.160 1614.990 2590.220 ;
        RECT 1779.810 2590.360 1780.130 2590.420 ;
        RECT 2132.170 2590.360 2132.490 2590.420 ;
        RECT 1779.810 2590.220 2132.490 2590.360 ;
        RECT 1779.810 2590.160 1780.130 2590.220 ;
        RECT 2132.170 2590.160 2132.490 2590.220 ;
        RECT 2179.550 2590.360 2179.870 2590.420 ;
        RECT 2220.490 2590.360 2220.810 2590.420 ;
        RECT 2179.550 2590.220 2220.810 2590.360 ;
        RECT 2179.550 2590.160 2179.870 2590.220 ;
        RECT 2220.490 2590.160 2220.810 2590.220 ;
        RECT 1496.910 2590.020 1497.230 2590.080 ;
        RECT 1593.970 2590.020 1594.290 2590.080 ;
        RECT 1496.910 2589.880 1594.290 2590.020 ;
        RECT 1496.910 2589.820 1497.230 2589.880 ;
        RECT 1593.970 2589.820 1594.290 2589.880 ;
        RECT 1702.530 2590.020 1702.850 2590.080 ;
        RECT 2152.870 2590.020 2153.190 2590.080 ;
        RECT 1702.530 2589.880 2153.190 2590.020 ;
        RECT 1702.530 2589.820 1702.850 2589.880 ;
        RECT 2152.870 2589.820 2153.190 2589.880 ;
        RECT 2183.690 2590.020 2184.010 2590.080 ;
        RECT 2227.850 2590.020 2228.170 2590.080 ;
        RECT 2276.150 2590.020 2276.470 2590.080 ;
        RECT 2183.690 2589.880 2276.470 2590.020 ;
        RECT 2183.690 2589.820 2184.010 2589.880 ;
        RECT 2227.850 2589.820 2228.170 2589.880 ;
        RECT 2276.150 2589.820 2276.470 2589.880 ;
        RECT 1483.110 2589.680 1483.430 2589.740 ;
        RECT 1587.070 2589.680 1587.390 2589.740 ;
        RECT 1483.110 2589.540 1587.390 2589.680 ;
        RECT 1483.110 2589.480 1483.430 2589.540 ;
        RECT 1587.070 2589.480 1587.390 2589.540 ;
        RECT 1614.210 2589.680 1614.530 2589.740 ;
        RECT 1662.970 2589.680 1663.290 2589.740 ;
        RECT 1614.210 2589.540 1663.290 2589.680 ;
        RECT 1614.210 2589.480 1614.530 2589.540 ;
        RECT 1662.970 2589.480 1663.290 2589.540 ;
        RECT 1707.590 2589.680 1707.910 2589.740 ;
        RECT 2159.770 2589.680 2160.090 2589.740 ;
        RECT 1707.590 2589.540 2160.090 2589.680 ;
        RECT 1707.590 2589.480 1707.910 2589.540 ;
        RECT 2159.770 2589.480 2160.090 2589.540 ;
        RECT 2170.350 2589.680 2170.670 2589.740 ;
        RECT 2215.890 2589.680 2216.210 2589.740 ;
        RECT 2170.350 2589.540 2216.210 2589.680 ;
        RECT 2170.350 2589.480 2170.670 2589.540 ;
        RECT 2215.890 2589.480 2216.210 2589.540 ;
        RECT 1586.610 2589.340 1586.930 2589.400 ;
        RECT 1642.270 2589.340 1642.590 2589.400 ;
        RECT 1586.610 2589.200 1642.590 2589.340 ;
        RECT 1586.610 2589.140 1586.930 2589.200 ;
        RECT 1642.270 2589.140 1642.590 2589.200 ;
        RECT 1652.390 2589.340 1652.710 2589.400 ;
        RECT 1678.610 2589.340 1678.930 2589.400 ;
        RECT 1652.390 2589.200 1678.930 2589.340 ;
        RECT 1652.390 2589.140 1652.710 2589.200 ;
        RECT 1678.610 2589.140 1678.930 2589.200 ;
        RECT 1718.170 2589.340 1718.490 2589.400 ;
        RECT 2180.470 2589.340 2180.790 2589.400 ;
        RECT 1718.170 2589.200 2180.790 2589.340 ;
        RECT 1718.170 2589.140 1718.490 2589.200 ;
        RECT 2180.470 2589.140 2180.790 2589.200 ;
        RECT 2184.610 2589.340 2184.930 2589.400 ;
        RECT 2186.450 2589.340 2186.770 2589.400 ;
        RECT 2232.910 2589.340 2233.230 2589.400 ;
        RECT 2184.610 2589.200 2233.230 2589.340 ;
        RECT 2184.610 2589.140 2184.930 2589.200 ;
        RECT 2186.450 2589.140 2186.770 2589.200 ;
        RECT 2232.910 2589.140 2233.230 2589.200 ;
        RECT 1503.350 2589.000 1503.670 2589.060 ;
        RECT 1600.870 2589.000 1601.190 2589.060 ;
        RECT 1503.350 2588.860 1601.190 2589.000 ;
        RECT 1503.350 2588.800 1503.670 2588.860 ;
        RECT 1600.870 2588.800 1601.190 2588.860 ;
        RECT 1607.310 2589.000 1607.630 2589.060 ;
        RECT 1656.070 2589.000 1656.390 2589.060 ;
        RECT 1607.310 2588.860 1656.390 2589.000 ;
        RECT 1607.310 2588.800 1607.630 2588.860 ;
        RECT 1656.070 2588.800 1656.390 2588.860 ;
        RECT 2162.990 2589.000 2163.310 2589.060 ;
        RECT 2209.450 2589.000 2209.770 2589.060 ;
        RECT 2214.510 2589.000 2214.830 2589.060 ;
        RECT 2162.990 2588.860 2214.830 2589.000 ;
        RECT 2162.990 2588.800 2163.310 2588.860 ;
        RECT 2209.450 2588.800 2209.770 2588.860 ;
        RECT 2214.510 2588.800 2214.830 2588.860 ;
        RECT 1558.550 2588.660 1558.870 2588.720 ;
        RECT 1631.230 2588.660 1631.550 2588.720 ;
        RECT 1558.550 2588.520 1631.550 2588.660 ;
        RECT 1558.550 2588.460 1558.870 2588.520 ;
        RECT 1631.230 2588.460 1631.550 2588.520 ;
        RECT 1669.410 2588.660 1669.730 2588.720 ;
        RECT 1690.570 2588.660 1690.890 2588.720 ;
        RECT 1669.410 2588.520 1690.890 2588.660 ;
        RECT 1669.410 2588.460 1669.730 2588.520 ;
        RECT 1690.570 2588.460 1690.890 2588.520 ;
        RECT 2190.590 2588.660 2190.910 2588.720 ;
        RECT 2235.670 2588.660 2235.990 2588.720 ;
        RECT 2190.590 2588.520 2235.990 2588.660 ;
        RECT 2190.590 2588.460 2190.910 2588.520 ;
        RECT 2235.670 2588.460 2235.990 2588.520 ;
        RECT 1551.650 2588.320 1551.970 2588.380 ;
        RECT 1621.570 2588.320 1621.890 2588.380 ;
        RECT 1551.650 2588.180 1621.890 2588.320 ;
        RECT 1551.650 2588.120 1551.970 2588.180 ;
        RECT 1621.570 2588.120 1621.890 2588.180 ;
        RECT 1641.810 2588.320 1642.130 2588.380 ;
        RECT 1669.870 2588.320 1670.190 2588.380 ;
        RECT 1641.810 2588.180 1670.190 2588.320 ;
        RECT 1641.810 2588.120 1642.130 2588.180 ;
        RECT 1669.870 2588.120 1670.190 2588.180 ;
        RECT 1731.510 2588.320 1731.830 2588.380 ;
        RECT 2194.270 2588.320 2194.590 2588.380 ;
        RECT 1731.510 2588.180 2194.590 2588.320 ;
        RECT 1731.510 2588.120 1731.830 2588.180 ;
        RECT 2194.270 2588.120 2194.590 2588.180 ;
        RECT 2204.390 2588.320 2204.710 2588.380 ;
        RECT 2249.470 2588.320 2249.790 2588.380 ;
        RECT 2204.390 2588.180 2249.790 2588.320 ;
        RECT 2204.390 2588.120 2204.710 2588.180 ;
        RECT 2249.470 2588.120 2249.790 2588.180 ;
        RECT 1441.710 2587.980 1442.030 2588.040 ;
        RECT 1566.370 2587.980 1566.690 2588.040 ;
        RECT 1441.710 2587.840 1566.690 2587.980 ;
        RECT 1441.710 2587.780 1442.030 2587.840 ;
        RECT 1566.370 2587.780 1566.690 2587.840 ;
        RECT 1586.150 2587.980 1586.470 2588.040 ;
        RECT 1630.770 2587.980 1631.090 2588.040 ;
        RECT 1635.370 2587.980 1635.690 2588.040 ;
        RECT 1586.150 2587.840 1631.090 2587.980 ;
        RECT 1586.150 2587.780 1586.470 2587.840 ;
        RECT 1630.770 2587.780 1631.090 2587.840 ;
        RECT 1631.320 2587.840 1635.690 2587.980 ;
        RECT 1427.910 2587.640 1428.230 2587.700 ;
        RECT 1559.470 2587.640 1559.790 2587.700 ;
        RECT 1427.910 2587.500 1559.790 2587.640 ;
        RECT 1427.910 2587.440 1428.230 2587.500 ;
        RECT 1559.470 2587.440 1559.790 2587.500 ;
        RECT 1572.810 2587.640 1573.130 2587.700 ;
        RECT 1631.320 2587.640 1631.460 2587.840 ;
        RECT 1635.370 2587.780 1635.690 2587.840 ;
        RECT 1638.590 2587.980 1638.910 2588.040 ;
        RECT 1662.970 2587.980 1663.290 2588.040 ;
        RECT 1638.590 2587.840 1663.290 2587.980 ;
        RECT 1638.590 2587.780 1638.910 2587.840 ;
        RECT 1662.970 2587.780 1663.290 2587.840 ;
        RECT 1713.110 2587.980 1713.430 2588.040 ;
        RECT 2173.570 2587.980 2173.890 2588.040 ;
        RECT 1713.110 2587.840 2173.890 2587.980 ;
        RECT 1713.110 2587.780 1713.430 2587.840 ;
        RECT 2173.570 2587.780 2173.890 2587.840 ;
        RECT 2197.490 2587.980 2197.810 2588.040 ;
        RECT 2243.950 2587.980 2244.270 2588.040 ;
        RECT 2197.490 2587.840 2244.270 2587.980 ;
        RECT 2197.490 2587.780 2197.810 2587.840 ;
        RECT 2243.950 2587.780 2244.270 2587.840 ;
        RECT 1572.810 2587.500 1631.460 2587.640 ;
        RECT 1631.690 2587.640 1632.010 2587.700 ;
        RECT 1649.170 2587.640 1649.490 2587.700 ;
        RECT 1631.690 2587.500 1649.490 2587.640 ;
        RECT 1572.810 2587.440 1573.130 2587.500 ;
        RECT 1631.690 2587.440 1632.010 2587.500 ;
        RECT 1649.170 2587.440 1649.490 2587.500 ;
        RECT 1666.190 2587.640 1666.510 2587.700 ;
        RECT 1683.670 2587.640 1683.990 2587.700 ;
        RECT 1666.190 2587.500 1683.990 2587.640 ;
        RECT 1666.190 2587.440 1666.510 2587.500 ;
        RECT 1683.670 2587.440 1683.990 2587.500 ;
        RECT 1686.890 2587.640 1687.210 2587.700 ;
        RECT 1697.470 2587.640 1697.790 2587.700 ;
        RECT 1686.890 2587.500 1697.790 2587.640 ;
        RECT 1686.890 2587.440 1687.210 2587.500 ;
        RECT 1697.470 2587.440 1697.790 2587.500 ;
        RECT 1736.570 2587.640 1736.890 2587.700 ;
        RECT 1742.090 2587.640 1742.410 2587.700 ;
        RECT 1736.570 2587.500 1742.410 2587.640 ;
        RECT 1736.570 2587.440 1736.890 2587.500 ;
        RECT 1742.090 2587.440 1742.410 2587.500 ;
        RECT 2168.970 2511.820 2169.290 2511.880 ;
        RECT 2170.350 2511.820 2170.670 2511.880 ;
        RECT 2168.970 2511.680 2170.670 2511.820 ;
        RECT 2168.970 2511.620 2169.290 2511.680 ;
        RECT 2170.350 2511.620 2170.670 2511.680 ;
        RECT 2168.050 2463.200 2168.370 2463.260 ;
        RECT 2169.430 2463.200 2169.750 2463.260 ;
        RECT 2168.050 2463.060 2169.750 2463.200 ;
        RECT 2168.050 2463.000 2168.370 2463.060 ;
        RECT 2169.430 2463.000 2169.750 2463.060 ;
        RECT 1487.710 2414.920 1488.030 2414.980 ;
        RECT 1887.910 2414.920 1888.230 2414.980 ;
        RECT 1487.710 2414.780 1888.230 2414.920 ;
        RECT 1487.710 2414.720 1488.030 2414.780 ;
        RECT 1887.910 2414.720 1888.230 2414.780 ;
        RECT 2166.210 2414.920 2166.530 2414.980 ;
        RECT 2240.270 2414.920 2240.590 2414.980 ;
        RECT 2166.210 2414.780 2240.590 2414.920 ;
        RECT 2166.210 2414.720 2166.530 2414.780 ;
        RECT 2240.270 2414.720 2240.590 2414.780 ;
        RECT 2276.610 2414.920 2276.930 2414.980 ;
        RECT 2449.570 2414.920 2449.890 2414.980 ;
        RECT 2276.610 2414.780 2449.890 2414.920 ;
        RECT 2276.610 2414.720 2276.930 2414.780 ;
        RECT 2449.570 2414.720 2449.890 2414.780 ;
        RECT 1488.170 2414.580 1488.490 2414.640 ;
        RECT 1898.950 2414.580 1899.270 2414.640 ;
        RECT 1488.170 2414.440 1899.270 2414.580 ;
        RECT 1488.170 2414.380 1488.490 2414.440 ;
        RECT 1898.950 2414.380 1899.270 2414.440 ;
        RECT 2133.090 2414.580 2133.410 2414.640 ;
        RECT 2197.490 2414.580 2197.810 2414.640 ;
        RECT 2133.090 2414.440 2197.810 2414.580 ;
        RECT 2133.090 2414.380 2133.410 2414.440 ;
        RECT 2197.490 2414.380 2197.810 2414.440 ;
        RECT 2283.510 2414.580 2283.830 2414.640 ;
        RECT 2460.150 2414.580 2460.470 2414.640 ;
        RECT 2283.510 2414.440 2460.470 2414.580 ;
        RECT 2283.510 2414.380 2283.830 2414.440 ;
        RECT 2460.150 2414.380 2460.470 2414.440 ;
        RECT 1488.630 2414.240 1488.950 2414.300 ;
        RECT 1911.370 2414.240 1911.690 2414.300 ;
        RECT 1488.630 2414.100 1911.690 2414.240 ;
        RECT 1488.630 2414.040 1488.950 2414.100 ;
        RECT 1911.370 2414.040 1911.690 2414.100 ;
        RECT 2173.110 2414.240 2173.430 2414.300 ;
        RECT 2251.310 2414.240 2251.630 2414.300 ;
        RECT 2173.110 2414.100 2251.630 2414.240 ;
        RECT 2173.110 2414.040 2173.430 2414.100 ;
        RECT 2251.310 2414.040 2251.630 2414.100 ;
        RECT 2290.410 2414.240 2290.730 2414.300 ;
        RECT 2471.190 2414.240 2471.510 2414.300 ;
        RECT 2290.410 2414.100 2471.510 2414.240 ;
        RECT 2290.410 2414.040 2290.730 2414.100 ;
        RECT 2471.190 2414.040 2471.510 2414.100 ;
        RECT 1489.090 2413.900 1489.410 2413.960 ;
        RECT 1920.570 2413.900 1920.890 2413.960 ;
        RECT 1489.090 2413.760 1920.890 2413.900 ;
        RECT 1489.090 2413.700 1489.410 2413.760 ;
        RECT 1920.570 2413.700 1920.890 2413.760 ;
        RECT 2180.470 2413.900 2180.790 2413.960 ;
        RECT 2183.690 2413.900 2184.010 2413.960 ;
        RECT 2180.470 2413.760 2184.010 2413.900 ;
        RECT 2180.470 2413.700 2180.790 2413.760 ;
        RECT 2183.690 2413.700 2184.010 2413.760 ;
        RECT 2186.910 2413.900 2187.230 2413.960 ;
        RECT 2272.930 2413.900 2273.250 2413.960 ;
        RECT 2186.910 2413.760 2273.250 2413.900 ;
        RECT 2186.910 2413.700 2187.230 2413.760 ;
        RECT 2272.930 2413.700 2273.250 2413.760 ;
        RECT 2297.310 2413.900 2297.630 2413.960 ;
        RECT 2482.230 2413.900 2482.550 2413.960 ;
        RECT 2297.310 2413.760 2482.550 2413.900 ;
        RECT 2297.310 2413.700 2297.630 2413.760 ;
        RECT 2482.230 2413.700 2482.550 2413.760 ;
        RECT 1489.550 2413.560 1489.870 2413.620 ;
        RECT 1932.070 2413.560 1932.390 2413.620 ;
        RECT 1489.550 2413.420 1932.390 2413.560 ;
        RECT 1489.550 2413.360 1489.870 2413.420 ;
        RECT 1932.070 2413.360 1932.390 2413.420 ;
        RECT 1956.910 2413.560 1957.230 2413.620 ;
        RECT 1959.210 2413.560 1959.530 2413.620 ;
        RECT 1956.910 2413.420 1959.530 2413.560 ;
        RECT 1956.910 2413.360 1957.230 2413.420 ;
        RECT 1959.210 2413.360 1959.530 2413.420 ;
        RECT 1990.030 2413.560 1990.350 2413.620 ;
        RECT 1993.250 2413.560 1993.570 2413.620 ;
        RECT 1990.030 2413.420 1993.570 2413.560 ;
        RECT 1990.030 2413.360 1990.350 2413.420 ;
        RECT 1993.250 2413.360 1993.570 2413.420 ;
        RECT 2180.010 2413.560 2180.330 2413.620 ;
        RECT 2263.270 2413.560 2263.590 2413.620 ;
        RECT 2180.010 2413.420 2263.590 2413.560 ;
        RECT 2180.010 2413.360 2180.330 2413.420 ;
        RECT 2263.270 2413.360 2263.590 2413.420 ;
        RECT 2303.750 2413.560 2304.070 2413.620 ;
        RECT 2493.270 2413.560 2493.590 2413.620 ;
        RECT 2303.750 2413.420 2493.590 2413.560 ;
        RECT 2303.750 2413.360 2304.070 2413.420 ;
        RECT 2493.270 2413.360 2493.590 2413.420 ;
        RECT 1545.210 2413.220 1545.530 2413.280 ;
        RECT 1997.850 2413.220 1998.170 2413.280 ;
        RECT 1545.210 2413.080 1998.170 2413.220 ;
        RECT 1545.210 2413.020 1545.530 2413.080 ;
        RECT 1997.850 2413.020 1998.170 2413.080 ;
        RECT 2122.050 2413.220 2122.370 2413.280 ;
        RECT 2190.590 2413.220 2190.910 2413.280 ;
        RECT 2122.050 2413.080 2190.910 2413.220 ;
        RECT 2122.050 2413.020 2122.370 2413.080 ;
        RECT 2190.590 2413.020 2190.910 2413.080 ;
        RECT 2193.810 2413.220 2194.130 2413.280 ;
        RECT 2284.430 2413.220 2284.750 2413.280 ;
        RECT 2193.810 2413.080 2284.750 2413.220 ;
        RECT 2193.810 2413.020 2194.130 2413.080 ;
        RECT 2284.430 2413.020 2284.750 2413.080 ;
        RECT 2311.110 2413.220 2311.430 2413.280 ;
        RECT 2515.350 2413.220 2515.670 2413.280 ;
        RECT 2311.110 2413.080 2515.670 2413.220 ;
        RECT 2311.110 2413.020 2311.430 2413.080 ;
        RECT 2515.350 2413.020 2515.670 2413.080 ;
        RECT 1439.410 2412.880 1439.730 2412.940 ;
        RECT 1441.710 2412.880 1442.030 2412.940 ;
        RECT 1439.410 2412.740 1442.030 2412.880 ;
        RECT 1439.410 2412.680 1439.730 2412.740 ;
        RECT 1441.710 2412.680 1442.030 2412.740 ;
        RECT 1494.610 2412.880 1494.930 2412.940 ;
        RECT 1496.910 2412.880 1497.230 2412.940 ;
        RECT 1494.610 2412.740 1497.230 2412.880 ;
        RECT 1494.610 2412.680 1494.930 2412.740 ;
        RECT 1496.910 2412.680 1497.230 2412.740 ;
        RECT 1527.730 2412.880 1528.050 2412.940 ;
        RECT 1531.410 2412.880 1531.730 2412.940 ;
        RECT 1527.730 2412.740 1531.730 2412.880 ;
        RECT 1527.730 2412.680 1528.050 2412.740 ;
        RECT 1531.410 2412.680 1531.730 2412.740 ;
        RECT 1551.190 2412.880 1551.510 2412.940 ;
        RECT 2008.890 2412.880 2009.210 2412.940 ;
        RECT 1551.190 2412.740 2009.210 2412.880 ;
        RECT 1551.190 2412.680 1551.510 2412.740 ;
        RECT 2008.890 2412.680 2009.210 2412.740 ;
        RECT 2045.230 2412.880 2045.550 2412.940 ;
        RECT 2048.910 2412.880 2049.230 2412.940 ;
        RECT 2045.230 2412.740 2049.230 2412.880 ;
        RECT 2045.230 2412.680 2045.550 2412.740 ;
        RECT 2048.910 2412.680 2049.230 2412.740 ;
        RECT 2111.010 2412.880 2111.330 2412.940 ;
        RECT 2184.610 2412.880 2184.930 2412.940 ;
        RECT 2111.010 2412.740 2184.930 2412.880 ;
        RECT 2111.010 2412.680 2111.330 2412.740 ;
        RECT 2184.610 2412.680 2184.930 2412.740 ;
        RECT 2193.350 2412.880 2193.670 2412.940 ;
        RECT 2295.010 2412.880 2295.330 2412.940 ;
        RECT 2193.350 2412.740 2295.330 2412.880 ;
        RECT 2193.350 2412.680 2193.670 2412.740 ;
        RECT 2295.010 2412.680 2295.330 2412.740 ;
        RECT 2304.210 2412.880 2304.530 2412.940 ;
        RECT 2504.770 2412.880 2505.090 2412.940 ;
        RECT 2304.210 2412.740 2505.090 2412.880 ;
        RECT 2304.210 2412.680 2304.530 2412.740 ;
        RECT 2504.770 2412.680 2505.090 2412.740 ;
        RECT 1552.110 2412.540 1552.430 2412.600 ;
        RECT 2019.930 2412.540 2020.250 2412.600 ;
        RECT 1552.110 2412.400 2020.250 2412.540 ;
        RECT 1552.110 2412.340 1552.430 2412.400 ;
        RECT 2019.930 2412.340 2020.250 2412.400 ;
        RECT 2099.970 2412.540 2100.290 2412.600 ;
        RECT 2180.470 2412.540 2180.790 2412.600 ;
        RECT 2099.970 2412.400 2180.790 2412.540 ;
        RECT 2099.970 2412.340 2100.290 2412.400 ;
        RECT 2180.470 2412.340 2180.790 2412.400 ;
        RECT 2214.510 2412.540 2214.830 2412.600 ;
        RECT 2324.910 2412.540 2325.230 2412.600 ;
        RECT 2537.430 2412.540 2537.750 2412.600 ;
        RECT 2214.510 2412.400 2319.160 2412.540 ;
        RECT 2214.510 2412.340 2214.830 2412.400 ;
        RECT 1559.010 2412.200 1559.330 2412.260 ;
        RECT 2030.970 2412.200 2031.290 2412.260 ;
        RECT 1559.010 2412.060 2031.290 2412.200 ;
        RECT 1559.010 2412.000 1559.330 2412.060 ;
        RECT 2030.970 2412.000 2031.290 2412.060 ;
        RECT 2086.630 2412.200 2086.950 2412.260 ;
        RECT 2176.790 2412.200 2177.110 2412.260 ;
        RECT 2086.630 2412.060 2177.110 2412.200 ;
        RECT 2086.630 2412.000 2086.950 2412.060 ;
        RECT 2176.790 2412.000 2177.110 2412.060 ;
        RECT 2200.710 2412.200 2201.030 2412.260 ;
        RECT 2306.050 2412.200 2306.370 2412.260 ;
        RECT 2200.710 2412.060 2306.370 2412.200 ;
        RECT 2200.710 2412.000 2201.030 2412.060 ;
        RECT 2306.050 2412.000 2306.370 2412.060 ;
        RECT 1406.750 2411.860 1407.070 2411.920 ;
        RECT 1898.030 2411.860 1898.350 2411.920 ;
        RECT 1406.750 2411.720 1898.350 2411.860 ;
        RECT 1406.750 2411.660 1407.070 2411.720 ;
        RECT 1898.030 2411.660 1898.350 2411.720 ;
        RECT 2076.050 2411.860 2076.370 2411.920 ;
        RECT 2168.970 2411.860 2169.290 2411.920 ;
        RECT 2076.050 2411.720 2169.290 2411.860 ;
        RECT 2076.050 2411.660 2076.370 2411.720 ;
        RECT 2168.970 2411.660 2169.290 2411.720 ;
        RECT 2207.610 2411.860 2207.930 2411.920 ;
        RECT 2318.470 2411.860 2318.790 2411.920 ;
        RECT 2207.610 2411.720 2318.790 2411.860 ;
        RECT 2319.020 2411.860 2319.160 2412.400 ;
        RECT 2324.910 2412.400 2537.750 2412.540 ;
        RECT 2324.910 2412.340 2325.230 2412.400 ;
        RECT 2537.430 2412.340 2537.750 2412.400 ;
        RECT 2319.390 2412.200 2319.710 2412.260 ;
        RECT 2526.390 2412.200 2526.710 2412.260 ;
        RECT 2319.390 2412.060 2526.710 2412.200 ;
        RECT 2319.390 2412.000 2319.710 2412.060 ;
        RECT 2526.390 2412.000 2526.710 2412.060 ;
        RECT 2328.130 2411.860 2328.450 2411.920 ;
        RECT 2319.020 2411.720 2328.450 2411.860 ;
        RECT 2207.610 2411.660 2207.930 2411.720 ;
        RECT 2318.470 2411.660 2318.790 2411.720 ;
        RECT 2328.130 2411.660 2328.450 2411.720 ;
        RECT 2331.810 2411.860 2332.130 2411.920 ;
        RECT 2548.470 2411.860 2548.790 2411.920 ;
        RECT 2331.810 2411.720 2548.790 2411.860 ;
        RECT 2331.810 2411.660 2332.130 2411.720 ;
        RECT 2548.470 2411.660 2548.790 2411.720 ;
        RECT 1511.630 2411.520 1511.950 2411.580 ;
        RECT 1559.470 2411.520 1559.790 2411.580 ;
        RECT 1511.630 2411.380 1559.790 2411.520 ;
        RECT 1511.630 2411.320 1511.950 2411.380 ;
        RECT 1559.470 2411.320 1559.790 2411.380 ;
        RECT 1609.610 2411.520 1609.930 2411.580 ;
        RECT 1656.070 2411.520 1656.390 2411.580 ;
        RECT 1609.610 2411.380 1656.390 2411.520 ;
        RECT 1609.610 2411.320 1609.930 2411.380 ;
        RECT 1656.070 2411.320 1656.390 2411.380 ;
        RECT 1702.990 2411.520 1703.310 2411.580 ;
        RECT 1752.670 2411.520 1752.990 2411.580 ;
        RECT 1702.990 2411.380 1752.990 2411.520 ;
        RECT 1702.990 2411.320 1703.310 2411.380 ;
        RECT 1752.670 2411.320 1752.990 2411.380 ;
        RECT 1800.510 2411.520 1800.830 2411.580 ;
        RECT 1835.470 2411.520 1835.790 2411.580 ;
        RECT 1932.530 2411.520 1932.850 2411.580 ;
        RECT 1800.510 2411.380 1835.790 2411.520 ;
        RECT 1800.510 2411.320 1800.830 2411.380 ;
        RECT 1835.470 2411.320 1835.790 2411.380 ;
        RECT 1897.200 2411.380 1932.850 2411.520 ;
        RECT 1487.250 2411.180 1487.570 2411.240 ;
        RECT 1510.710 2411.180 1511.030 2411.240 ;
        RECT 1487.250 2411.040 1511.030 2411.180 ;
        RECT 1487.250 2410.980 1487.570 2411.040 ;
        RECT 1510.710 2410.980 1511.030 2411.040 ;
        RECT 1511.170 2411.180 1511.490 2411.240 ;
        RECT 1703.450 2411.180 1703.770 2411.240 ;
        RECT 1511.170 2411.040 1703.770 2411.180 ;
        RECT 1511.170 2410.980 1511.490 2411.040 ;
        RECT 1703.450 2410.980 1703.770 2411.040 ;
        RECT 1714.030 2411.180 1714.350 2411.240 ;
        RECT 1876.870 2411.180 1877.190 2411.240 ;
        RECT 1714.030 2411.040 1877.190 2411.180 ;
        RECT 1714.030 2410.980 1714.350 2411.040 ;
        RECT 1876.870 2410.980 1877.190 2411.040 ;
        RECT 1877.330 2411.180 1877.650 2411.240 ;
        RECT 1897.200 2411.180 1897.340 2411.380 ;
        RECT 1932.530 2411.320 1932.850 2411.380 ;
        RECT 1945.870 2411.520 1946.190 2411.580 ;
        RECT 2067.310 2411.520 2067.630 2411.580 ;
        RECT 2162.990 2411.520 2163.310 2411.580 ;
        RECT 1945.870 2411.380 1980.140 2411.520 ;
        RECT 1945.870 2411.320 1946.190 2411.380 ;
        RECT 1877.330 2411.040 1897.340 2411.180 ;
        RECT 1980.000 2411.180 1980.140 2411.380 ;
        RECT 2067.310 2411.380 2163.310 2411.520 ;
        RECT 2067.310 2411.320 2067.630 2411.380 ;
        RECT 2162.990 2411.320 2163.310 2411.380 ;
        RECT 2221.410 2411.520 2221.730 2411.580 ;
        RECT 2340.090 2411.520 2340.410 2411.580 ;
        RECT 2221.410 2411.380 2340.410 2411.520 ;
        RECT 2221.410 2411.320 2221.730 2411.380 ;
        RECT 2340.090 2411.320 2340.410 2411.380 ;
        RECT 2345.150 2411.520 2345.470 2411.580 ;
        RECT 2570.550 2411.520 2570.870 2411.580 ;
        RECT 2345.150 2411.380 2570.870 2411.520 ;
        RECT 2345.150 2411.320 2345.470 2411.380 ;
        RECT 2570.550 2411.320 2570.870 2411.380 ;
        RECT 2144.130 2411.180 2144.450 2411.240 ;
        RECT 2204.390 2411.180 2204.710 2411.240 ;
        RECT 1980.000 2411.040 1994.400 2411.180 ;
        RECT 1877.330 2410.980 1877.650 2411.040 ;
        RECT 1486.790 2410.840 1487.110 2410.900 ;
        RECT 1510.250 2410.840 1510.570 2410.900 ;
        RECT 1486.790 2410.700 1510.570 2410.840 ;
        RECT 1486.790 2410.640 1487.110 2410.700 ;
        RECT 1510.250 2410.640 1510.570 2410.700 ;
        RECT 1538.310 2410.840 1538.630 2410.900 ;
        RECT 1865.830 2410.840 1866.150 2410.900 ;
        RECT 1538.310 2410.700 1866.150 2410.840 ;
        RECT 1994.260 2410.840 1994.400 2411.040 ;
        RECT 2144.130 2411.040 2204.710 2411.180 ;
        RECT 2144.130 2410.980 2144.450 2411.040 ;
        RECT 2204.390 2410.980 2204.710 2411.040 ;
        RECT 2269.710 2411.180 2270.030 2411.240 ;
        RECT 2438.070 2411.180 2438.390 2411.240 ;
        RECT 2269.710 2411.040 2438.390 2411.180 ;
        RECT 2269.710 2410.980 2270.030 2411.040 ;
        RECT 2438.070 2410.980 2438.390 2411.040 ;
        RECT 2053.050 2410.840 2053.370 2410.900 ;
        RECT 1994.260 2410.700 2053.370 2410.840 ;
        RECT 1538.310 2410.640 1538.630 2410.700 ;
        RECT 1865.830 2410.640 1866.150 2410.700 ;
        RECT 2053.050 2410.640 2053.370 2410.700 ;
        RECT 2269.250 2410.840 2269.570 2410.900 ;
        RECT 2428.870 2410.840 2429.190 2410.900 ;
        RECT 2269.250 2410.700 2429.190 2410.840 ;
        RECT 2269.250 2410.640 2269.570 2410.700 ;
        RECT 2428.870 2410.640 2429.190 2410.700 ;
        RECT 1626.630 2410.500 1626.950 2410.560 ;
        RECT 1638.590 2410.500 1638.910 2410.560 ;
        RECT 1626.630 2410.360 1638.910 2410.500 ;
        RECT 1626.630 2410.300 1626.950 2410.360 ;
        RECT 1638.590 2410.300 1638.910 2410.360 ;
        RECT 1648.710 2410.500 1649.030 2410.560 ;
        RECT 1652.390 2410.500 1652.710 2410.560 ;
        RECT 1648.710 2410.360 1652.710 2410.500 ;
        RECT 1648.710 2410.300 1649.030 2410.360 ;
        RECT 1652.390 2410.300 1652.710 2410.360 ;
        RECT 1659.750 2410.500 1660.070 2410.560 ;
        RECT 1666.190 2410.500 1666.510 2410.560 ;
        RECT 1702.990 2410.500 1703.310 2410.560 ;
        RECT 1659.750 2410.360 1666.510 2410.500 ;
        RECT 1659.750 2410.300 1660.070 2410.360 ;
        RECT 1666.190 2410.300 1666.510 2410.360 ;
        RECT 1666.740 2410.360 1703.310 2410.500 ;
        RECT 1559.470 2410.160 1559.790 2410.220 ;
        RECT 1593.970 2410.160 1594.290 2410.220 ;
        RECT 1559.470 2410.020 1594.290 2410.160 ;
        RECT 1559.470 2409.960 1559.790 2410.020 ;
        RECT 1593.970 2409.960 1594.290 2410.020 ;
        RECT 1656.070 2410.160 1656.390 2410.220 ;
        RECT 1666.740 2410.160 1666.880 2410.360 ;
        RECT 1702.990 2410.300 1703.310 2410.360 ;
        RECT 1731.510 2410.500 1731.830 2410.560 ;
        RECT 1733.810 2410.500 1734.130 2410.560 ;
        RECT 1731.510 2410.360 1734.130 2410.500 ;
        RECT 1731.510 2410.300 1731.830 2410.360 ;
        RECT 1733.810 2410.300 1734.130 2410.360 ;
        RECT 1742.090 2410.500 1742.410 2410.560 ;
        RECT 1745.770 2410.500 1746.090 2410.560 ;
        RECT 1742.090 2410.360 1746.090 2410.500 ;
        RECT 1742.090 2410.300 1742.410 2410.360 ;
        RECT 1745.770 2410.300 1746.090 2410.360 ;
        RECT 1746.230 2410.500 1746.550 2410.560 ;
        RECT 1755.430 2410.500 1755.750 2410.560 ;
        RECT 1746.230 2410.360 1755.750 2410.500 ;
        RECT 1746.230 2410.300 1746.550 2410.360 ;
        RECT 1755.430 2410.300 1755.750 2410.360 ;
        RECT 1791.770 2410.500 1792.090 2410.560 ;
        RECT 2089.850 2410.500 2090.170 2410.560 ;
        RECT 1791.770 2410.360 2090.170 2410.500 ;
        RECT 1791.770 2410.300 1792.090 2410.360 ;
        RECT 2089.850 2410.300 2090.170 2410.360 ;
        RECT 2262.810 2410.500 2263.130 2410.560 ;
        RECT 2416.450 2410.500 2416.770 2410.560 ;
        RECT 2262.810 2410.360 2416.770 2410.500 ;
        RECT 2262.810 2410.300 2263.130 2410.360 ;
        RECT 2416.450 2410.300 2416.770 2410.360 ;
        RECT 1656.070 2410.020 1666.880 2410.160 ;
        RECT 1681.830 2410.160 1682.150 2410.220 ;
        RECT 1686.890 2410.160 1687.210 2410.220 ;
        RECT 1681.830 2410.020 1687.210 2410.160 ;
        RECT 1656.070 2409.960 1656.390 2410.020 ;
        RECT 1681.830 2409.960 1682.150 2410.020 ;
        RECT 1686.890 2409.960 1687.210 2410.020 ;
        RECT 1703.450 2410.160 1703.770 2410.220 ;
        RECT 1714.030 2410.160 1714.350 2410.220 ;
        RECT 1703.450 2410.020 1714.350 2410.160 ;
        RECT 1703.450 2409.960 1703.770 2410.020 ;
        RECT 1714.030 2409.960 1714.350 2410.020 ;
        RECT 1752.670 2410.160 1752.990 2410.220 ;
        RECT 1800.510 2410.160 1800.830 2410.220 ;
        RECT 1752.670 2410.020 1800.830 2410.160 ;
        RECT 1752.670 2409.960 1752.990 2410.020 ;
        RECT 1800.510 2409.960 1800.830 2410.020 ;
        RECT 1802.810 2410.160 1803.130 2410.220 ;
        RECT 2089.390 2410.160 2089.710 2410.220 ;
        RECT 1802.810 2410.020 2089.710 2410.160 ;
        RECT 1802.810 2409.960 1803.130 2410.020 ;
        RECT 2089.390 2409.960 2089.710 2410.020 ;
        RECT 2255.910 2410.160 2256.230 2410.220 ;
        RECT 2405.410 2410.160 2405.730 2410.220 ;
        RECT 2255.910 2410.020 2405.730 2410.160 ;
        RECT 2255.910 2409.960 2256.230 2410.020 ;
        RECT 2405.410 2409.960 2405.730 2410.020 ;
        RECT 1593.510 2409.820 1593.830 2409.880 ;
        RECT 1631.690 2409.820 1632.010 2409.880 ;
        RECT 1593.510 2409.680 1632.010 2409.820 ;
        RECT 1593.510 2409.620 1593.830 2409.680 ;
        RECT 1631.690 2409.620 1632.010 2409.680 ;
        RECT 1744.850 2409.820 1745.170 2409.880 ;
        RECT 1766.470 2409.820 1766.790 2409.880 ;
        RECT 1744.850 2409.680 1766.790 2409.820 ;
        RECT 1744.850 2409.620 1745.170 2409.680 ;
        RECT 1766.470 2409.620 1766.790 2409.680 ;
        RECT 1813.850 2409.820 1814.170 2409.880 ;
        RECT 2088.930 2409.820 2089.250 2409.880 ;
        RECT 1813.850 2409.680 2089.250 2409.820 ;
        RECT 1813.850 2409.620 1814.170 2409.680 ;
        RECT 2088.930 2409.620 2089.250 2409.680 ;
        RECT 2249.010 2409.820 2249.330 2409.880 ;
        RECT 2394.370 2409.820 2394.690 2409.880 ;
        RECT 2249.010 2409.680 2394.690 2409.820 ;
        RECT 2249.010 2409.620 2249.330 2409.680 ;
        RECT 2394.370 2409.620 2394.690 2409.680 ;
        RECT 1472.530 2409.480 1472.850 2409.540 ;
        RECT 1476.210 2409.480 1476.530 2409.540 ;
        RECT 1472.530 2409.340 1476.530 2409.480 ;
        RECT 1472.530 2409.280 1472.850 2409.340 ;
        RECT 1476.210 2409.280 1476.530 2409.340 ;
        RECT 1582.470 2409.480 1582.790 2409.540 ;
        RECT 1586.610 2409.480 1586.930 2409.540 ;
        RECT 1582.470 2409.340 1586.930 2409.480 ;
        RECT 1582.470 2409.280 1582.790 2409.340 ;
        RECT 1586.610 2409.280 1586.930 2409.340 ;
        RECT 1604.550 2409.480 1604.870 2409.540 ;
        RECT 1607.310 2409.480 1607.630 2409.540 ;
        RECT 1604.550 2409.340 1607.630 2409.480 ;
        RECT 1604.550 2409.280 1604.870 2409.340 ;
        RECT 1607.310 2409.280 1607.630 2409.340 ;
        RECT 1637.670 2409.480 1637.990 2409.540 ;
        RECT 1641.810 2409.480 1642.130 2409.540 ;
        RECT 1637.670 2409.340 1642.130 2409.480 ;
        RECT 1637.670 2409.280 1637.990 2409.340 ;
        RECT 1641.810 2409.280 1642.130 2409.340 ;
        RECT 1824.890 2409.480 1825.210 2409.540 ;
        RECT 2088.470 2409.480 2088.790 2409.540 ;
        RECT 1824.890 2409.340 2088.790 2409.480 ;
        RECT 1824.890 2409.280 1825.210 2409.340 ;
        RECT 2088.470 2409.280 2088.790 2409.340 ;
        RECT 2235.210 2409.480 2235.530 2409.540 ;
        RECT 2373.670 2409.480 2373.990 2409.540 ;
        RECT 2235.210 2409.340 2373.990 2409.480 ;
        RECT 2235.210 2409.280 2235.530 2409.340 ;
        RECT 2373.670 2409.280 2373.990 2409.340 ;
        RECT 1835.010 2409.140 1835.330 2409.200 ;
        RECT 2088.010 2409.140 2088.330 2409.200 ;
        RECT 1835.010 2409.000 2088.330 2409.140 ;
        RECT 1835.010 2408.940 1835.330 2409.000 ;
        RECT 2088.010 2408.940 2088.330 2409.000 ;
        RECT 2242.110 2409.140 2242.430 2409.200 ;
        RECT 2383.330 2409.140 2383.650 2409.200 ;
        RECT 2242.110 2409.000 2383.650 2409.140 ;
        RECT 2242.110 2408.940 2242.430 2409.000 ;
        RECT 2383.330 2408.940 2383.650 2409.000 ;
        RECT 1692.870 2408.800 1693.190 2408.860 ;
        RECT 1697.010 2408.800 1697.330 2408.860 ;
        RECT 1692.870 2408.660 1697.330 2408.800 ;
        RECT 1692.870 2408.600 1693.190 2408.660 ;
        RECT 1697.010 2408.600 1697.330 2408.660 ;
        RECT 1846.970 2408.800 1847.290 2408.860 ;
        RECT 2087.550 2408.800 2087.870 2408.860 ;
        RECT 1846.970 2408.660 2087.870 2408.800 ;
        RECT 1846.970 2408.600 1847.290 2408.660 ;
        RECT 2087.550 2408.600 2087.870 2408.660 ;
        RECT 2227.850 2408.800 2228.170 2408.860 ;
        RECT 2361.250 2408.800 2361.570 2408.860 ;
        RECT 2227.850 2408.660 2361.570 2408.800 ;
        RECT 2227.850 2408.600 2228.170 2408.660 ;
        RECT 2361.250 2408.600 2361.570 2408.660 ;
        RECT 1858.010 2408.460 1858.330 2408.520 ;
        RECT 2087.090 2408.460 2087.410 2408.520 ;
        RECT 1858.010 2408.320 2087.410 2408.460 ;
        RECT 1858.010 2408.260 1858.330 2408.320 ;
        RECT 2087.090 2408.260 2087.410 2408.320 ;
        RECT 2228.310 2408.460 2228.630 2408.520 ;
        RECT 2350.210 2408.460 2350.530 2408.520 ;
        RECT 2228.310 2408.320 2350.530 2408.460 ;
        RECT 2228.310 2408.260 2228.630 2408.320 ;
        RECT 2350.210 2408.260 2350.530 2408.320 ;
      LAYER met1 ;
        RECT 1404.670 1204.460 2595.010 2392.000 ;
      LAYER met1 ;
        RECT 2587.570 1197.040 2587.890 1197.100 ;
        RECT 2593.550 1197.040 2593.870 1197.100 ;
        RECT 2587.570 1196.900 2593.870 1197.040 ;
        RECT 2587.570 1196.840 2587.890 1196.900 ;
        RECT 2593.550 1196.840 2593.870 1196.900 ;
        RECT 1668.490 1193.640 1668.810 1193.700 ;
        RECT 1722.770 1193.640 1723.090 1193.700 ;
        RECT 1668.490 1193.500 1723.090 1193.640 ;
        RECT 1668.490 1193.440 1668.810 1193.500 ;
        RECT 1722.770 1193.440 1723.090 1193.500 ;
        RECT 2131.710 1193.640 2132.030 1193.700 ;
        RECT 2245.790 1193.640 2246.110 1193.700 ;
        RECT 2131.710 1193.500 2246.110 1193.640 ;
        RECT 2131.710 1193.440 2132.030 1193.500 ;
        RECT 2245.790 1193.440 2246.110 1193.500 ;
        RECT 2363.090 1193.640 2363.410 1193.700 ;
        RECT 2471.190 1193.640 2471.510 1193.700 ;
        RECT 2363.090 1193.500 2471.510 1193.640 ;
        RECT 2363.090 1193.440 2363.410 1193.500 ;
        RECT 2471.190 1193.440 2471.510 1193.500 ;
        RECT 1662.510 1193.300 1662.830 1193.360 ;
        RECT 1733.810 1193.300 1734.130 1193.360 ;
        RECT 1662.510 1193.160 1734.130 1193.300 ;
        RECT 1662.510 1193.100 1662.830 1193.160 ;
        RECT 1733.810 1193.100 1734.130 1193.160 ;
        RECT 2122.050 1193.300 2122.370 1193.360 ;
        RECT 2252.690 1193.300 2253.010 1193.360 ;
        RECT 2122.050 1193.160 2253.010 1193.300 ;
        RECT 2122.050 1193.100 2122.370 1193.160 ;
        RECT 2252.690 1193.100 2253.010 1193.160 ;
        RECT 2276.150 1193.300 2276.470 1193.360 ;
        RECT 2383.790 1193.300 2384.110 1193.360 ;
        RECT 2276.150 1193.160 2384.110 1193.300 ;
        RECT 2276.150 1193.100 2276.470 1193.160 ;
        RECT 2383.790 1193.100 2384.110 1193.160 ;
        RECT 1655.610 1192.960 1655.930 1193.020 ;
        RECT 1745.770 1192.960 1746.090 1193.020 ;
        RECT 1655.610 1192.820 1746.090 1192.960 ;
        RECT 1655.610 1192.760 1655.930 1192.820 ;
        RECT 1745.770 1192.760 1746.090 1192.820 ;
        RECT 1969.790 1192.960 1970.110 1193.020 ;
        RECT 2030.970 1192.960 2031.290 1193.020 ;
        RECT 1969.790 1192.820 2031.290 1192.960 ;
        RECT 1969.790 1192.760 1970.110 1192.820 ;
        RECT 2030.970 1192.760 2031.290 1192.820 ;
        RECT 2111.010 1192.960 2111.330 1193.020 ;
        RECT 2259.590 1192.960 2259.910 1193.020 ;
        RECT 2111.010 1192.820 2259.910 1192.960 ;
        RECT 2111.010 1192.760 2111.330 1192.820 ;
        RECT 2259.590 1192.760 2259.910 1192.820 ;
        RECT 2287.190 1192.960 2287.510 1193.020 ;
        RECT 2290.410 1192.960 2290.730 1193.020 ;
        RECT 2384.250 1192.960 2384.570 1193.020 ;
        RECT 2287.190 1192.820 2290.730 1192.960 ;
        RECT 2287.190 1192.760 2287.510 1192.820 ;
        RECT 2290.410 1192.760 2290.730 1192.820 ;
        RECT 2290.960 1192.820 2384.570 1192.960 ;
        RECT 1582.470 1192.620 1582.790 1192.680 ;
        RECT 1586.610 1192.620 1586.930 1192.680 ;
        RECT 1582.470 1192.480 1586.930 1192.620 ;
        RECT 1582.470 1192.420 1582.790 1192.480 ;
        RECT 1586.610 1192.420 1586.930 1192.480 ;
        RECT 1667.570 1192.620 1667.890 1192.680 ;
        RECT 1755.430 1192.620 1755.750 1192.680 ;
        RECT 1667.570 1192.480 1755.750 1192.620 ;
        RECT 1667.570 1192.420 1667.890 1192.480 ;
        RECT 1755.430 1192.420 1755.750 1192.480 ;
        RECT 1902.170 1192.620 1902.490 1192.680 ;
        RECT 1997.850 1192.620 1998.170 1192.680 ;
        RECT 1902.170 1192.480 1998.170 1192.620 ;
        RECT 1902.170 1192.420 1902.490 1192.480 ;
        RECT 1997.850 1192.420 1998.170 1192.480 ;
        RECT 2099.970 1192.620 2100.290 1192.680 ;
        RECT 2265.110 1192.620 2265.430 1192.680 ;
        RECT 2290.960 1192.620 2291.100 1192.820 ;
        RECT 2384.250 1192.760 2384.570 1192.820 ;
        RECT 2099.970 1192.480 2261.660 1192.620 ;
        RECT 2099.970 1192.420 2100.290 1192.480 ;
        RECT 1472.530 1192.280 1472.850 1192.340 ;
        RECT 1476.210 1192.280 1476.530 1192.340 ;
        RECT 1472.530 1192.140 1476.530 1192.280 ;
        RECT 1472.530 1192.080 1472.850 1192.140 ;
        RECT 1476.210 1192.080 1476.530 1192.140 ;
        RECT 1641.350 1192.280 1641.670 1192.340 ;
        RECT 1766.470 1192.280 1766.790 1192.340 ;
        RECT 1641.350 1192.140 1766.790 1192.280 ;
        RECT 1641.350 1192.080 1641.670 1192.140 ;
        RECT 1766.470 1192.080 1766.790 1192.140 ;
        RECT 1901.710 1192.280 1902.030 1192.340 ;
        RECT 2008.890 1192.280 2009.210 1192.340 ;
        RECT 1901.710 1192.140 2009.210 1192.280 ;
        RECT 1901.710 1192.080 1902.030 1192.140 ;
        RECT 2008.890 1192.080 2009.210 1192.140 ;
        RECT 2076.510 1192.280 2076.830 1192.340 ;
        RECT 2261.520 1192.280 2261.660 1192.480 ;
        RECT 2265.110 1192.480 2291.100 1192.620 ;
        RECT 2317.550 1192.620 2317.870 1192.680 ;
        RECT 2449.570 1192.620 2449.890 1192.680 ;
        RECT 2317.550 1192.480 2449.890 1192.620 ;
        RECT 2265.110 1192.420 2265.430 1192.480 ;
        RECT 2317.550 1192.420 2317.870 1192.480 ;
        RECT 2449.570 1192.420 2449.890 1192.480 ;
        RECT 2266.490 1192.280 2266.810 1192.340 ;
        RECT 2076.510 1192.140 2261.200 1192.280 ;
        RECT 2261.520 1192.140 2266.810 1192.280 ;
        RECT 2076.510 1192.080 2076.830 1192.140 ;
        RECT 1559.010 1191.940 1559.330 1192.000 ;
        RECT 1714.490 1191.940 1714.810 1192.000 ;
        RECT 1559.010 1191.800 1714.810 1191.940 ;
        RECT 1559.010 1191.740 1559.330 1191.800 ;
        RECT 1714.490 1191.740 1714.810 1191.800 ;
        RECT 1901.250 1191.940 1901.570 1192.000 ;
        RECT 2019.930 1191.940 2020.250 1192.000 ;
        RECT 1901.250 1191.800 2020.250 1191.940 ;
        RECT 1901.250 1191.740 1901.570 1191.800 ;
        RECT 2019.930 1191.740 2020.250 1191.800 ;
        RECT 2067.310 1191.940 2067.630 1192.000 ;
        RECT 2260.510 1191.940 2260.830 1192.000 ;
        RECT 2067.310 1191.800 2260.830 1191.940 ;
        RECT 2261.060 1191.940 2261.200 1192.140 ;
        RECT 2266.490 1192.080 2266.810 1192.140 ;
        RECT 2311.110 1192.280 2311.430 1192.340 ;
        RECT 2460.150 1192.280 2460.470 1192.340 ;
        RECT 2311.110 1192.140 2460.470 1192.280 ;
        RECT 2311.110 1192.080 2311.430 1192.140 ;
        RECT 2460.150 1192.080 2460.470 1192.140 ;
        RECT 2280.290 1191.940 2280.610 1192.000 ;
        RECT 2261.060 1191.800 2280.610 1191.940 ;
        RECT 2067.310 1191.740 2067.630 1191.800 ;
        RECT 2260.510 1191.740 2260.830 1191.800 ;
        RECT 2280.290 1191.740 2280.610 1191.800 ;
        RECT 2283.510 1191.940 2283.830 1192.000 ;
        RECT 2504.770 1191.940 2505.090 1192.000 ;
        RECT 2283.510 1191.800 2505.090 1191.940 ;
        RECT 2283.510 1191.740 2283.830 1191.800 ;
        RECT 2504.770 1191.740 2505.090 1191.800 ;
        RECT 1549.810 1191.600 1550.130 1191.660 ;
        RECT 1721.390 1191.600 1721.710 1191.660 ;
        RECT 1549.810 1191.460 1721.710 1191.600 ;
        RECT 1549.810 1191.400 1550.130 1191.460 ;
        RECT 1721.390 1191.400 1721.710 1191.460 ;
        RECT 1855.710 1191.600 1856.030 1191.660 ;
        RECT 1975.770 1191.600 1976.090 1191.660 ;
        RECT 1855.710 1191.460 1976.090 1191.600 ;
        RECT 1855.710 1191.400 1856.030 1191.460 ;
        RECT 1975.770 1191.400 1976.090 1191.460 ;
        RECT 1997.390 1191.600 1997.710 1191.660 ;
        RECT 2042.470 1191.600 2042.790 1191.660 ;
        RECT 1997.390 1191.460 2042.790 1191.600 ;
        RECT 1997.390 1191.400 1997.710 1191.460 ;
        RECT 2042.470 1191.400 2042.790 1191.460 ;
        RECT 2089.390 1191.600 2089.710 1191.660 ;
        RECT 2273.390 1191.600 2273.710 1191.660 ;
        RECT 2089.390 1191.460 2273.710 1191.600 ;
        RECT 2089.390 1191.400 2089.710 1191.460 ;
        RECT 2273.390 1191.400 2273.710 1191.460 ;
        RECT 2276.610 1191.600 2276.930 1191.660 ;
        RECT 2526.390 1191.600 2526.710 1191.660 ;
        RECT 2276.610 1191.460 2526.710 1191.600 ;
        RECT 2276.610 1191.400 2276.930 1191.460 ;
        RECT 2526.390 1191.400 2526.710 1191.460 ;
        RECT 1527.730 1191.260 1528.050 1191.320 ;
        RECT 1714.950 1191.260 1715.270 1191.320 ;
        RECT 1527.730 1191.120 1715.270 1191.260 ;
        RECT 1527.730 1191.060 1528.050 1191.120 ;
        RECT 1714.950 1191.060 1715.270 1191.120 ;
        RECT 1965.650 1191.260 1965.970 1191.320 ;
        RECT 2260.050 1191.260 2260.370 1191.320 ;
        RECT 1965.650 1191.120 2260.370 1191.260 ;
        RECT 1965.650 1191.060 1965.970 1191.120 ;
        RECT 2260.050 1191.060 2260.370 1191.120 ;
        RECT 2260.510 1191.260 2260.830 1191.320 ;
        RECT 2281.210 1191.260 2281.530 1191.320 ;
        RECT 2260.510 1191.120 2281.530 1191.260 ;
        RECT 2260.510 1191.060 2260.830 1191.120 ;
        RECT 2281.210 1191.060 2281.530 1191.120 ;
        RECT 2296.850 1191.260 2297.170 1191.320 ;
        RECT 2482.230 1191.260 2482.550 1191.320 ;
        RECT 2296.850 1191.120 2482.550 1191.260 ;
        RECT 2296.850 1191.060 2297.170 1191.120 ;
        RECT 2482.230 1191.060 2482.550 1191.120 ;
        RECT 1417.330 1190.920 1417.650 1190.980 ;
        RECT 1490.010 1190.920 1490.330 1190.980 ;
        RECT 1417.330 1190.780 1490.330 1190.920 ;
        RECT 1417.330 1190.720 1417.650 1190.780 ;
        RECT 1490.010 1190.720 1490.330 1190.780 ;
        RECT 1516.690 1190.920 1517.010 1190.980 ;
        RECT 1707.590 1190.920 1707.910 1190.980 ;
        RECT 1516.690 1190.780 1707.910 1190.920 ;
        RECT 1516.690 1190.720 1517.010 1190.780 ;
        RECT 1707.590 1190.720 1707.910 1190.780 ;
        RECT 1900.790 1190.920 1901.110 1190.980 ;
        RECT 2053.050 1190.920 2053.370 1190.980 ;
        RECT 1900.790 1190.780 2053.370 1190.920 ;
        RECT 1900.790 1190.720 1901.110 1190.780 ;
        RECT 2053.050 1190.720 2053.370 1190.780 ;
        RECT 2144.130 1190.920 2144.450 1190.980 ;
        RECT 2238.890 1190.920 2239.210 1190.980 ;
        RECT 2144.130 1190.780 2239.210 1190.920 ;
        RECT 2144.130 1190.720 2144.450 1190.780 ;
        RECT 2238.890 1190.720 2239.210 1190.780 ;
        RECT 2242.110 1190.920 2242.430 1190.980 ;
        RECT 2581.590 1190.920 2581.910 1190.980 ;
        RECT 2242.110 1190.780 2581.910 1190.920 ;
        RECT 2242.110 1190.720 2242.430 1190.780 ;
        RECT 2581.590 1190.720 2581.910 1190.780 ;
        RECT 1538.310 1190.580 1538.630 1190.640 ;
        RECT 1735.190 1190.580 1735.510 1190.640 ;
        RECT 1538.310 1190.440 1735.510 1190.580 ;
        RECT 1538.310 1190.380 1538.630 1190.440 ;
        RECT 1735.190 1190.380 1735.510 1190.440 ;
        RECT 1802.810 1190.580 1803.130 1190.640 ;
        RECT 2369.990 1190.580 2370.310 1190.640 ;
        RECT 1802.810 1190.440 2370.310 1190.580 ;
        RECT 1802.810 1190.380 1803.130 1190.440 ;
        RECT 2369.990 1190.380 2370.310 1190.440 ;
        RECT 1427.910 1190.240 1428.230 1190.300 ;
        RECT 1728.290 1190.240 1728.610 1190.300 ;
        RECT 1427.910 1190.100 1728.610 1190.240 ;
        RECT 1427.910 1190.040 1428.230 1190.100 ;
        RECT 1728.290 1190.040 1728.610 1190.100 ;
        RECT 1869.050 1190.240 1869.370 1190.300 ;
        RECT 2481.770 1190.240 2482.090 1190.300 ;
        RECT 1869.050 1190.100 2482.090 1190.240 ;
        RECT 1869.050 1190.040 1869.370 1190.100 ;
        RECT 2481.770 1190.040 2482.090 1190.100 ;
        RECT 2260.050 1189.900 2260.370 1189.960 ;
        RECT 2287.190 1189.900 2287.510 1189.960 ;
        RECT 2260.050 1189.760 2287.510 1189.900 ;
        RECT 2260.050 1189.700 2260.370 1189.760 ;
        RECT 2287.190 1189.700 2287.510 1189.760 ;
        RECT 2324.450 1189.900 2324.770 1189.960 ;
        RECT 2428.870 1189.900 2429.190 1189.960 ;
        RECT 2324.450 1189.760 2429.190 1189.900 ;
        RECT 2324.450 1189.700 2324.770 1189.760 ;
        RECT 2428.870 1189.700 2429.190 1189.760 ;
        RECT 2364.010 1189.560 2364.330 1189.620 ;
        RECT 2438.070 1189.560 2438.390 1189.620 ;
        RECT 2364.010 1189.420 2438.390 1189.560 ;
        RECT 2364.010 1189.360 2364.330 1189.420 ;
        RECT 2438.070 1189.360 2438.390 1189.420 ;
        RECT 1675.850 1189.220 1676.170 1189.280 ;
        RECT 1711.730 1189.220 1712.050 1189.280 ;
        RECT 1675.850 1189.080 1712.050 1189.220 ;
        RECT 1675.850 1189.020 1676.170 1189.080 ;
        RECT 1711.730 1189.020 1712.050 1189.080 ;
        RECT 2338.710 1189.220 2339.030 1189.280 ;
        RECT 2405.410 1189.220 2405.730 1189.280 ;
        RECT 2338.710 1189.080 2405.730 1189.220 ;
        RECT 2338.710 1189.020 2339.030 1189.080 ;
        RECT 2405.410 1189.020 2405.730 1189.080 ;
        RECT 2309.270 1188.880 2309.590 1188.940 ;
        RECT 2364.470 1188.880 2364.790 1188.940 ;
        RECT 2309.270 1188.740 2364.790 1188.880 ;
        RECT 2309.270 1188.680 2309.590 1188.740 ;
        RECT 2364.470 1188.680 2364.790 1188.740 ;
        RECT 1659.750 1188.540 1660.070 1188.600 ;
        RECT 1697.930 1188.540 1698.250 1188.600 ;
        RECT 1659.750 1188.400 1698.250 1188.540 ;
        RECT 1659.750 1188.340 1660.070 1188.400 ;
        RECT 1697.930 1188.340 1698.250 1188.400 ;
        RECT 1880.090 1188.540 1880.410 1188.600 ;
        RECT 1884.230 1188.540 1884.550 1188.600 ;
        RECT 1880.090 1188.400 1884.550 1188.540 ;
        RECT 1880.090 1188.340 1880.410 1188.400 ;
        RECT 1884.230 1188.340 1884.550 1188.400 ;
        RECT 2351.590 1188.540 2351.910 1188.600 ;
        RECT 2383.330 1188.540 2383.650 1188.600 ;
        RECT 2351.590 1188.400 2383.650 1188.540 ;
        RECT 2351.590 1188.340 2351.910 1188.400 ;
        RECT 2383.330 1188.340 2383.650 1188.400 ;
        RECT 1676.310 1188.200 1676.630 1188.260 ;
        RECT 1700.690 1188.200 1701.010 1188.260 ;
        RECT 1676.310 1188.060 1701.010 1188.200 ;
        RECT 1676.310 1188.000 1676.630 1188.060 ;
        RECT 1700.690 1188.000 1701.010 1188.060 ;
        RECT 1669.410 1187.860 1669.730 1187.920 ;
        RECT 1691.030 1187.860 1691.350 1187.920 ;
        RECT 1669.410 1187.720 1691.350 1187.860 ;
        RECT 1669.410 1187.660 1669.730 1187.720 ;
        RECT 1691.030 1187.660 1691.350 1187.720 ;
        RECT 1686.890 1187.520 1687.210 1187.580 ;
        RECT 1657.080 1187.380 1687.210 1187.520 ;
        RECT 1439.410 1187.180 1439.730 1187.240 ;
        RECT 1441.710 1187.180 1442.030 1187.240 ;
        RECT 1439.410 1187.040 1442.030 1187.180 ;
        RECT 1439.410 1186.980 1439.730 1187.040 ;
        RECT 1441.710 1186.980 1442.030 1187.040 ;
        RECT 1494.610 1187.180 1494.930 1187.240 ;
        RECT 1496.910 1187.180 1497.230 1187.240 ;
        RECT 1494.610 1187.040 1497.230 1187.180 ;
        RECT 1494.610 1186.980 1494.930 1187.040 ;
        RECT 1496.910 1186.980 1497.230 1187.040 ;
        RECT 1604.550 1187.180 1604.870 1187.240 ;
        RECT 1607.310 1187.180 1607.630 1187.240 ;
        RECT 1604.550 1187.040 1607.630 1187.180 ;
        RECT 1604.550 1186.980 1604.870 1187.040 ;
        RECT 1607.310 1186.980 1607.630 1187.040 ;
        RECT 1637.670 1187.180 1637.990 1187.240 ;
        RECT 1641.810 1187.180 1642.130 1187.240 ;
        RECT 1637.670 1187.040 1642.130 1187.180 ;
        RECT 1637.670 1186.980 1637.990 1187.040 ;
        RECT 1641.810 1186.980 1642.130 1187.040 ;
        RECT 1648.710 1187.180 1649.030 1187.240 ;
        RECT 1657.080 1187.180 1657.220 1187.380 ;
        RECT 1686.890 1187.320 1687.210 1187.380 ;
        RECT 1834.090 1187.520 1834.410 1187.580 ;
        RECT 1843.750 1187.520 1844.070 1187.580 ;
        RECT 1834.090 1187.380 1844.070 1187.520 ;
        RECT 1834.090 1187.320 1834.410 1187.380 ;
        RECT 1843.750 1187.320 1844.070 1187.380 ;
        RECT 2331.350 1187.520 2331.670 1187.580 ;
        RECT 2363.550 1187.520 2363.870 1187.580 ;
        RECT 2331.350 1187.380 2363.870 1187.520 ;
        RECT 2331.350 1187.320 2331.670 1187.380 ;
        RECT 2363.550 1187.320 2363.870 1187.380 ;
        RECT 1648.710 1187.040 1657.220 1187.180 ;
        RECT 1668.490 1187.180 1668.810 1187.240 ;
        RECT 1669.410 1187.180 1669.730 1187.240 ;
        RECT 1668.490 1187.040 1669.730 1187.180 ;
        RECT 1648.710 1186.980 1649.030 1187.040 ;
        RECT 1668.490 1186.980 1668.810 1187.040 ;
        RECT 1669.410 1186.980 1669.730 1187.040 ;
        RECT 1684.130 1187.180 1684.450 1187.240 ;
        RECT 1690.570 1187.180 1690.890 1187.240 ;
        RECT 1684.130 1187.040 1690.890 1187.180 ;
        RECT 1684.130 1186.980 1684.450 1187.040 ;
        RECT 1690.570 1186.980 1690.890 1187.040 ;
        RECT 1824.890 1187.180 1825.210 1187.240 ;
        RECT 1831.790 1187.180 1832.110 1187.240 ;
        RECT 1824.890 1187.040 1832.110 1187.180 ;
        RECT 1824.890 1186.980 1825.210 1187.040 ;
        RECT 1831.790 1186.980 1832.110 1187.040 ;
        RECT 1835.010 1187.180 1835.330 1187.240 ;
        RECT 1856.170 1187.180 1856.490 1187.240 ;
        RECT 1835.010 1187.040 1856.490 1187.180 ;
        RECT 1835.010 1186.980 1835.330 1187.040 ;
        RECT 1856.170 1186.980 1856.490 1187.040 ;
        RECT 1913.210 1187.180 1913.530 1187.240 ;
        RECT 1917.810 1187.180 1918.130 1187.240 ;
        RECT 1913.210 1187.040 1918.130 1187.180 ;
        RECT 1913.210 1186.980 1913.530 1187.040 ;
        RECT 1917.810 1186.980 1918.130 1187.040 ;
        RECT 1934.830 1187.180 1935.150 1187.240 ;
        RECT 1938.510 1187.180 1938.830 1187.240 ;
        RECT 1934.830 1187.040 1938.830 1187.180 ;
        RECT 1934.830 1186.980 1935.150 1187.040 ;
        RECT 1938.510 1186.980 1938.830 1187.040 ;
        RECT 1956.910 1187.180 1957.230 1187.240 ;
        RECT 1959.210 1187.180 1959.530 1187.240 ;
        RECT 1956.910 1187.040 1959.530 1187.180 ;
        RECT 1956.910 1186.980 1957.230 1187.040 ;
        RECT 1959.210 1186.980 1959.530 1187.040 ;
        RECT 1976.690 1187.180 1977.010 1187.240 ;
        RECT 1987.270 1187.180 1987.590 1187.240 ;
        RECT 1976.690 1187.040 1987.590 1187.180 ;
        RECT 1976.690 1186.980 1977.010 1187.040 ;
        RECT 1987.270 1186.980 1987.590 1187.040 ;
        RECT 2320.310 1187.180 2320.630 1187.240 ;
        RECT 2324.910 1187.180 2325.230 1187.240 ;
        RECT 2320.310 1187.040 2325.230 1187.180 ;
        RECT 2320.310 1186.980 2320.630 1187.040 ;
        RECT 2324.910 1186.980 2325.230 1187.040 ;
        RECT 2342.390 1187.180 2342.710 1187.240 ;
        RECT 2345.610 1187.180 2345.930 1187.240 ;
        RECT 2342.390 1187.040 2345.930 1187.180 ;
        RECT 2342.390 1186.980 2342.710 1187.040 ;
        RECT 2345.610 1186.980 2345.930 1187.040 ;
        RECT 1648.710 1159.300 1649.030 1159.360 ;
        RECT 1667.570 1159.300 1667.890 1159.360 ;
        RECT 1648.710 1159.160 1667.890 1159.300 ;
        RECT 1648.710 1159.100 1649.030 1159.160 ;
        RECT 1667.570 1159.100 1667.890 1159.160 ;
        RECT 1682.290 1159.300 1682.610 1159.360 ;
        RECT 1684.130 1159.300 1684.450 1159.360 ;
        RECT 1682.290 1159.160 1684.450 1159.300 ;
        RECT 1682.290 1159.100 1682.610 1159.160 ;
        RECT 1684.130 1159.100 1684.450 1159.160 ;
        RECT 1682.750 1104.220 1683.070 1104.280 ;
        RECT 1683.210 1104.220 1683.530 1104.280 ;
        RECT 1682.750 1104.080 1683.530 1104.220 ;
        RECT 1682.750 1104.020 1683.070 1104.080 ;
        RECT 1683.210 1104.020 1683.530 1104.080 ;
        RECT 1683.210 1076.820 1683.530 1077.080 ;
        RECT 1683.300 1076.400 1683.440 1076.820 ;
        RECT 1683.210 1076.140 1683.530 1076.400 ;
        RECT 1462.410 1051.860 1462.730 1051.920 ;
        RECT 1496.450 1051.860 1496.770 1051.920 ;
        RECT 1462.410 1051.720 1496.770 1051.860 ;
        RECT 1462.410 1051.660 1462.730 1051.720 ;
        RECT 1496.450 1051.660 1496.770 1051.720 ;
        RECT 2287.190 1028.400 2287.510 1028.460 ;
        RECT 2288.110 1028.400 2288.430 1028.460 ;
        RECT 2287.190 1028.260 2288.430 1028.400 ;
        RECT 2287.190 1028.200 2287.510 1028.260 ;
        RECT 2288.110 1028.200 2288.430 1028.260 ;
        RECT 2352.050 1028.060 2352.370 1028.120 ;
        RECT 2359.870 1028.060 2360.190 1028.120 ;
        RECT 2352.050 1027.920 2360.190 1028.060 ;
        RECT 2352.050 1027.860 2352.370 1027.920 ;
        RECT 2359.870 1027.860 2360.190 1027.920 ;
        RECT 2352.510 1026.360 2352.830 1026.420 ;
        RECT 2373.670 1026.360 2373.990 1026.420 ;
        RECT 2352.510 1026.220 2373.990 1026.360 ;
        RECT 2352.510 1026.160 2352.830 1026.220 ;
        RECT 2373.670 1026.160 2373.990 1026.220 ;
        RECT 2330.890 1026.020 2331.210 1026.080 ;
        RECT 2415.070 1026.020 2415.390 1026.080 ;
        RECT 2330.890 1025.880 2415.390 1026.020 ;
        RECT 2330.890 1025.820 2331.210 1025.880 ;
        RECT 2415.070 1025.820 2415.390 1025.880 ;
        RECT 2345.150 1025.680 2345.470 1025.740 ;
        RECT 2394.370 1025.680 2394.690 1025.740 ;
        RECT 2345.150 1025.540 2394.690 1025.680 ;
        RECT 2345.150 1025.480 2345.470 1025.540 ;
        RECT 2394.370 1025.480 2394.690 1025.540 ;
        RECT 2255.910 1025.340 2256.230 1025.400 ;
        RECT 2415.070 1025.340 2415.390 1025.400 ;
        RECT 2255.910 1025.200 2415.390 1025.340 ;
        RECT 2255.910 1025.140 2256.230 1025.200 ;
        RECT 2415.070 1025.140 2415.390 1025.200 ;
        RECT 2241.650 1025.000 2241.970 1025.060 ;
        RECT 2421.970 1025.000 2422.290 1025.060 ;
        RECT 2241.650 1024.860 2422.290 1025.000 ;
        RECT 2241.650 1024.800 2241.970 1024.860 ;
        RECT 2421.970 1024.800 2422.290 1024.860 ;
        RECT 1890.210 1024.660 1890.530 1024.720 ;
        RECT 2450.950 1024.660 2451.270 1024.720 ;
        RECT 1890.210 1024.520 2451.270 1024.660 ;
        RECT 1890.210 1024.460 1890.530 1024.520 ;
        RECT 2450.950 1024.460 2451.270 1024.520 ;
        RECT 2363.550 1021.940 2363.870 1022.000 ;
        RECT 2363.550 1021.800 2365.160 1021.940 ;
        RECT 2363.550 1021.740 2363.870 1021.800 ;
        RECT 2363.180 1021.460 2364.700 1021.600 ;
        RECT 1686.890 1021.260 1687.210 1021.320 ;
        RECT 1704.370 1021.260 1704.690 1021.320 ;
        RECT 1686.890 1021.120 1704.690 1021.260 ;
        RECT 1686.890 1021.060 1687.210 1021.120 ;
        RECT 1704.370 1021.060 1704.690 1021.120 ;
        RECT 1706.210 1021.260 1706.530 1021.320 ;
        RECT 1731.970 1021.260 1732.290 1021.320 ;
        RECT 1706.210 1021.120 1732.290 1021.260 ;
        RECT 1706.210 1021.060 1706.530 1021.120 ;
        RECT 1731.970 1021.060 1732.290 1021.120 ;
        RECT 1735.190 1021.260 1735.510 1021.320 ;
        RECT 1759.570 1021.260 1759.890 1021.320 ;
        RECT 1735.190 1021.120 1759.890 1021.260 ;
        RECT 1735.190 1021.060 1735.510 1021.120 ;
        RECT 1759.570 1021.060 1759.890 1021.120 ;
        RECT 1831.790 1021.260 1832.110 1021.320 ;
        RECT 1842.370 1021.260 1842.690 1021.320 ;
        RECT 1831.790 1021.120 1842.690 1021.260 ;
        RECT 1831.790 1021.060 1832.110 1021.120 ;
        RECT 1842.370 1021.060 1842.690 1021.120 ;
        RECT 1918.270 1021.260 1918.590 1021.320 ;
        RECT 1966.110 1021.260 1966.430 1021.320 ;
        RECT 1918.270 1021.120 1966.430 1021.260 ;
        RECT 1918.270 1021.060 1918.590 1021.120 ;
        RECT 1966.110 1021.060 1966.430 1021.120 ;
        RECT 2014.870 1021.260 2015.190 1021.320 ;
        RECT 2062.710 1021.260 2063.030 1021.320 ;
        RECT 2014.870 1021.120 2063.030 1021.260 ;
        RECT 2014.870 1021.060 2015.190 1021.120 ;
        RECT 2062.710 1021.060 2063.030 1021.120 ;
        RECT 2111.470 1021.260 2111.790 1021.320 ;
        RECT 2159.310 1021.260 2159.630 1021.320 ;
        RECT 2111.470 1021.120 2159.630 1021.260 ;
        RECT 2111.470 1021.060 2111.790 1021.120 ;
        RECT 2159.310 1021.060 2159.630 1021.120 ;
        RECT 2252.690 1021.260 2253.010 1021.320 ;
        RECT 2254.530 1021.260 2254.850 1021.320 ;
        RECT 2303.290 1021.260 2303.610 1021.320 ;
        RECT 2252.690 1021.120 2303.610 1021.260 ;
        RECT 2252.690 1021.060 2253.010 1021.120 ;
        RECT 2254.530 1021.060 2254.850 1021.120 ;
        RECT 2303.290 1021.060 2303.610 1021.120 ;
        RECT 2324.910 1021.260 2325.230 1021.320 ;
        RECT 2363.180 1021.260 2363.320 1021.460 ;
        RECT 2324.910 1021.120 2363.320 1021.260 ;
        RECT 2324.910 1021.060 2325.230 1021.120 ;
        RECT 1496.910 1020.720 1497.230 1020.980 ;
        RECT 1641.810 1020.920 1642.130 1020.980 ;
        RECT 1711.270 1020.920 1711.590 1020.980 ;
        RECT 1641.810 1020.780 1711.590 1020.920 ;
        RECT 1641.810 1020.720 1642.130 1020.780 ;
        RECT 1711.270 1020.720 1711.590 1020.780 ;
        RECT 1717.250 1020.920 1717.570 1020.980 ;
        RECT 1741.630 1020.920 1741.950 1020.980 ;
        RECT 1748.070 1020.920 1748.390 1020.980 ;
        RECT 1717.250 1020.780 1748.390 1020.920 ;
        RECT 1717.250 1020.720 1717.570 1020.780 ;
        RECT 1741.630 1020.720 1741.950 1020.780 ;
        RECT 1748.070 1020.720 1748.390 1020.780 ;
        RECT 1752.210 1020.920 1752.530 1020.980 ;
        RECT 1786.710 1020.920 1787.030 1020.980 ;
        RECT 1752.210 1020.780 1787.030 1020.920 ;
        RECT 1752.210 1020.720 1752.530 1020.780 ;
        RECT 1786.710 1020.720 1787.030 1020.780 ;
        RECT 1787.630 1020.920 1787.950 1020.980 ;
        RECT 2214.970 1020.920 2215.290 1020.980 ;
        RECT 1787.630 1020.780 2215.290 1020.920 ;
        RECT 1787.630 1020.720 1787.950 1020.780 ;
        RECT 2214.970 1020.720 2215.290 1020.780 ;
        RECT 2266.490 1020.920 2266.810 1020.980 ;
        RECT 2312.030 1020.920 2312.350 1020.980 ;
        RECT 2266.490 1020.780 2312.350 1020.920 ;
        RECT 2266.490 1020.720 2266.810 1020.780 ;
        RECT 2312.030 1020.720 2312.350 1020.780 ;
        RECT 2318.010 1020.920 2318.330 1020.980 ;
        RECT 2364.010 1020.920 2364.330 1020.980 ;
        RECT 2318.010 1020.780 2364.330 1020.920 ;
        RECT 2364.560 1020.920 2364.700 1021.460 ;
        RECT 2365.020 1021.260 2365.160 1021.800 ;
        RECT 2373.670 1021.260 2373.990 1021.320 ;
        RECT 2365.020 1021.120 2373.990 1021.260 ;
        RECT 2373.670 1021.060 2373.990 1021.120 ;
        RECT 2383.790 1021.260 2384.110 1021.320 ;
        RECT 2403.110 1021.260 2403.430 1021.320 ;
        RECT 2383.790 1021.120 2403.430 1021.260 ;
        RECT 2383.790 1021.060 2384.110 1021.120 ;
        RECT 2403.110 1021.060 2403.430 1021.120 ;
        RECT 2380.570 1020.920 2380.890 1020.980 ;
        RECT 2364.560 1020.780 2380.890 1020.920 ;
        RECT 2318.010 1020.720 2318.330 1020.780 ;
        RECT 2364.010 1020.720 2364.330 1020.780 ;
        RECT 2380.570 1020.720 2380.890 1020.780 ;
        RECT 2384.250 1020.920 2384.570 1020.980 ;
        RECT 2408.170 1020.920 2408.490 1020.980 ;
        RECT 2384.250 1020.780 2408.490 1020.920 ;
        RECT 2384.250 1020.720 2384.570 1020.780 ;
        RECT 2408.170 1020.720 2408.490 1020.780 ;
        RECT 1497.000 1020.580 1497.140 1020.720 ;
        RECT 1787.170 1020.580 1787.490 1020.640 ;
        RECT 1497.000 1020.440 1787.490 1020.580 ;
        RECT 1787.170 1020.380 1787.490 1020.440 ;
        RECT 1790.390 1020.580 1790.710 1020.640 ;
        RECT 2208.070 1020.580 2208.390 1020.640 ;
        RECT 1790.390 1020.440 2208.390 1020.580 ;
        RECT 1790.390 1020.380 1790.710 1020.440 ;
        RECT 2208.070 1020.380 2208.390 1020.440 ;
        RECT 2245.790 1020.580 2246.110 1020.640 ;
        RECT 2293.630 1020.580 2293.950 1020.640 ;
        RECT 2245.790 1020.440 2293.950 1020.580 ;
        RECT 2245.790 1020.380 2246.110 1020.440 ;
        RECT 2293.630 1020.380 2293.950 1020.440 ;
        RECT 2353.890 1020.580 2354.210 1020.640 ;
        RECT 2363.550 1020.580 2363.870 1020.640 ;
        RECT 2353.890 1020.440 2363.870 1020.580 ;
        RECT 2353.890 1020.380 2354.210 1020.440 ;
        RECT 2363.550 1020.380 2363.870 1020.440 ;
        RECT 2364.470 1020.580 2364.790 1020.640 ;
        RECT 2387.470 1020.580 2387.790 1020.640 ;
        RECT 2364.470 1020.440 2387.790 1020.580 ;
        RECT 2364.470 1020.380 2364.790 1020.440 ;
        RECT 2387.470 1020.380 2387.790 1020.440 ;
        RECT 1503.810 1020.240 1504.130 1020.300 ;
        RECT 1780.270 1020.240 1780.590 1020.300 ;
        RECT 1503.810 1020.100 1780.590 1020.240 ;
        RECT 1503.810 1020.040 1504.130 1020.100 ;
        RECT 1780.270 1020.040 1780.590 1020.100 ;
        RECT 1800.050 1020.240 1800.370 1020.300 ;
        RECT 1821.670 1020.240 1821.990 1020.300 ;
        RECT 1800.050 1020.100 1821.990 1020.240 ;
        RECT 1800.050 1020.040 1800.370 1020.100 ;
        RECT 1821.670 1020.040 1821.990 1020.100 ;
        RECT 1869.510 1020.240 1869.830 1020.300 ;
        RECT 1918.270 1020.240 1918.590 1020.300 ;
        RECT 1869.510 1020.100 1918.590 1020.240 ;
        RECT 1869.510 1020.040 1869.830 1020.100 ;
        RECT 1918.270 1020.040 1918.590 1020.100 ;
        RECT 1966.110 1020.240 1966.430 1020.300 ;
        RECT 2014.870 1020.240 2015.190 1020.300 ;
        RECT 1966.110 1020.100 2015.190 1020.240 ;
        RECT 1966.110 1020.040 1966.430 1020.100 ;
        RECT 2014.870 1020.040 2015.190 1020.100 ;
        RECT 2062.710 1020.240 2063.030 1020.300 ;
        RECT 2111.470 1020.240 2111.790 1020.300 ;
        RECT 2062.710 1020.100 2111.790 1020.240 ;
        RECT 2062.710 1020.040 2063.030 1020.100 ;
        RECT 2111.470 1020.040 2111.790 1020.100 ;
        RECT 2159.310 1020.240 2159.630 1020.300 ;
        RECT 2194.270 1020.240 2194.590 1020.300 ;
        RECT 2159.310 1020.100 2194.590 1020.240 ;
        RECT 2159.310 1020.040 2159.630 1020.100 ;
        RECT 2194.270 1020.040 2194.590 1020.100 ;
        RECT 2269.710 1020.240 2270.030 1020.300 ;
        RECT 2532.370 1020.240 2532.690 1020.300 ;
        RECT 2269.710 1020.100 2532.690 1020.240 ;
        RECT 2269.710 1020.040 2270.030 1020.100 ;
        RECT 2532.370 1020.040 2532.690 1020.100 ;
        RECT 1572.810 1019.900 1573.130 1019.960 ;
        RECT 1745.770 1019.900 1746.090 1019.960 ;
        RECT 1572.810 1019.760 1746.090 1019.900 ;
        RECT 1572.810 1019.700 1573.130 1019.760 ;
        RECT 1745.770 1019.700 1746.090 1019.760 ;
        RECT 1759.110 1019.900 1759.430 1019.960 ;
        RECT 1806.030 1019.900 1806.350 1019.960 ;
        RECT 2180.470 1019.900 2180.790 1019.960 ;
        RECT 1759.110 1019.760 2180.790 1019.900 ;
        RECT 1759.110 1019.700 1759.430 1019.760 ;
        RECT 1806.030 1019.700 1806.350 1019.760 ;
        RECT 2180.470 1019.700 2180.790 1019.760 ;
        RECT 2276.610 1019.900 2276.930 1019.960 ;
        RECT 2511.670 1019.900 2511.990 1019.960 ;
        RECT 2276.610 1019.760 2511.990 1019.900 ;
        RECT 2276.610 1019.700 2276.930 1019.760 ;
        RECT 2511.670 1019.700 2511.990 1019.760 ;
        RECT 1586.610 1019.560 1586.930 1019.620 ;
        RECT 1738.870 1019.560 1739.190 1019.620 ;
        RECT 1586.610 1019.420 1739.190 1019.560 ;
        RECT 1586.610 1019.360 1586.930 1019.420 ;
        RECT 1738.870 1019.360 1739.190 1019.420 ;
        RECT 1807.870 1019.560 1808.190 1019.620 ;
        RECT 1812.930 1019.560 1813.250 1019.620 ;
        RECT 2173.570 1019.560 2173.890 1019.620 ;
        RECT 1807.870 1019.420 2173.890 1019.560 ;
        RECT 1807.870 1019.360 1808.190 1019.420 ;
        RECT 1812.930 1019.360 1813.250 1019.420 ;
        RECT 2173.570 1019.360 2173.890 1019.420 ;
        RECT 2238.890 1019.560 2239.210 1019.620 ;
        RECT 2242.110 1019.560 2242.430 1019.620 ;
        RECT 2287.190 1019.560 2287.510 1019.620 ;
        RECT 2238.890 1019.420 2287.510 1019.560 ;
        RECT 2238.890 1019.360 2239.210 1019.420 ;
        RECT 2242.110 1019.360 2242.430 1019.420 ;
        RECT 2287.190 1019.360 2287.510 1019.420 ;
        RECT 2289.950 1019.560 2290.270 1019.620 ;
        RECT 2490.970 1019.560 2491.290 1019.620 ;
        RECT 2289.950 1019.420 2491.290 1019.560 ;
        RECT 2289.950 1019.360 2290.270 1019.420 ;
        RECT 2490.970 1019.360 2491.290 1019.420 ;
        RECT 1593.510 1019.220 1593.830 1019.280 ;
        RECT 1679.990 1019.220 1680.310 1019.280 ;
        RECT 1714.950 1019.220 1715.270 1019.280 ;
        RECT 1766.470 1019.220 1766.790 1019.280 ;
        RECT 1593.510 1019.080 1680.310 1019.220 ;
        RECT 1593.510 1019.020 1593.830 1019.080 ;
        RECT 1679.990 1019.020 1680.310 1019.080 ;
        RECT 1680.540 1019.080 1714.720 1019.220 ;
        RECT 1607.310 1018.880 1607.630 1018.940 ;
        RECT 1680.540 1018.880 1680.680 1019.080 ;
        RECT 1607.310 1018.740 1680.680 1018.880 ;
        RECT 1714.580 1018.880 1714.720 1019.080 ;
        RECT 1714.950 1019.080 1766.790 1019.220 ;
        RECT 1714.950 1019.020 1715.270 1019.080 ;
        RECT 1766.470 1019.020 1766.790 1019.080 ;
        RECT 1772.910 1019.220 1773.230 1019.280 ;
        RECT 1817.530 1019.220 1817.850 1019.280 ;
        RECT 2159.770 1019.220 2160.090 1019.280 ;
        RECT 1772.910 1019.080 2160.090 1019.220 ;
        RECT 1772.910 1019.020 1773.230 1019.080 ;
        RECT 1817.530 1019.020 1817.850 1019.080 ;
        RECT 2159.770 1019.020 2160.090 1019.080 ;
        RECT 2290.410 1019.220 2290.730 1019.280 ;
        RECT 2394.370 1019.220 2394.690 1019.280 ;
        RECT 2290.410 1019.080 2394.690 1019.220 ;
        RECT 2290.410 1019.020 2290.730 1019.080 ;
        RECT 2394.370 1019.020 2394.690 1019.080 ;
        RECT 1725.070 1018.880 1725.390 1018.940 ;
        RECT 1714.580 1018.740 1725.390 1018.880 ;
        RECT 1607.310 1018.680 1607.630 1018.740 ;
        RECT 1725.070 1018.680 1725.390 1018.740 ;
        RECT 1728.290 1018.880 1728.610 1018.940 ;
        RECT 1821.670 1018.880 1821.990 1018.940 ;
        RECT 1823.970 1018.880 1824.290 1018.940 ;
        RECT 2152.870 1018.880 2153.190 1018.940 ;
        RECT 1728.290 1018.740 1821.990 1018.880 ;
        RECT 1728.290 1018.680 1728.610 1018.740 ;
        RECT 1821.670 1018.680 1821.990 1018.740 ;
        RECT 1822.220 1018.740 2153.190 1018.880 ;
        RECT 1614.210 1018.540 1614.530 1018.600 ;
        RECT 1718.170 1018.540 1718.490 1018.600 ;
        RECT 1773.370 1018.540 1773.690 1018.600 ;
        RECT 1807.870 1018.540 1808.190 1018.600 ;
        RECT 1614.210 1018.400 1718.490 1018.540 ;
        RECT 1614.210 1018.340 1614.530 1018.400 ;
        RECT 1718.170 1018.340 1718.490 1018.400 ;
        RECT 1718.720 1018.400 1773.690 1018.540 ;
        RECT 1628.010 1018.200 1628.330 1018.260 ;
        RECT 1707.590 1018.200 1707.910 1018.260 ;
        RECT 1718.720 1018.200 1718.860 1018.400 ;
        RECT 1773.370 1018.340 1773.690 1018.400 ;
        RECT 1773.920 1018.400 1808.190 1018.540 ;
        RECT 1628.010 1018.060 1707.360 1018.200 ;
        RECT 1628.010 1018.000 1628.330 1018.060 ;
        RECT 1679.990 1017.860 1680.310 1017.920 ;
        RECT 1707.220 1017.860 1707.360 1018.060 ;
        RECT 1707.590 1018.060 1718.860 1018.200 ;
        RECT 1731.970 1018.200 1732.290 1018.260 ;
        RECT 1735.650 1018.200 1735.970 1018.260 ;
        RECT 1766.010 1018.200 1766.330 1018.260 ;
        RECT 1773.920 1018.200 1774.060 1018.400 ;
        RECT 1807.870 1018.340 1808.190 1018.400 ;
        RECT 1731.970 1018.060 1747.840 1018.200 ;
        RECT 1707.590 1018.000 1707.910 1018.060 ;
        RECT 1731.970 1018.000 1732.290 1018.060 ;
        RECT 1735.650 1018.000 1735.970 1018.060 ;
        RECT 1711.270 1017.860 1711.590 1017.920 ;
        RECT 1679.990 1017.720 1706.900 1017.860 ;
        RECT 1707.220 1017.720 1711.590 1017.860 ;
        RECT 1679.990 1017.660 1680.310 1017.720 ;
        RECT 1641.810 1017.520 1642.130 1017.580 ;
        RECT 1689.650 1017.520 1689.970 1017.580 ;
        RECT 1706.210 1017.520 1706.530 1017.580 ;
        RECT 1641.810 1017.380 1706.530 1017.520 ;
        RECT 1706.760 1017.520 1706.900 1017.720 ;
        RECT 1711.270 1017.660 1711.590 1017.720 ;
        RECT 1713.200 1017.720 1747.380 1017.860 ;
        RECT 1712.190 1017.520 1712.510 1017.580 ;
        RECT 1706.760 1017.380 1712.510 1017.520 ;
        RECT 1641.810 1017.320 1642.130 1017.380 ;
        RECT 1689.650 1017.320 1689.970 1017.380 ;
        RECT 1706.210 1017.320 1706.530 1017.380 ;
        RECT 1712.190 1017.320 1712.510 1017.380 ;
        RECT 1654.690 1017.180 1655.010 1017.240 ;
        RECT 1700.690 1017.180 1701.010 1017.240 ;
        RECT 1713.200 1017.180 1713.340 1017.720 ;
        RECT 1713.570 1017.520 1713.890 1017.580 ;
        RECT 1731.970 1017.520 1732.290 1017.580 ;
        RECT 1713.570 1017.380 1732.290 1017.520 ;
        RECT 1713.570 1017.320 1713.890 1017.380 ;
        RECT 1731.970 1017.320 1732.290 1017.380 ;
        RECT 1718.170 1017.180 1718.490 1017.240 ;
        RECT 1747.240 1017.180 1747.380 1017.720 ;
        RECT 1747.700 1017.520 1747.840 1018.060 ;
        RECT 1766.010 1018.060 1774.060 1018.200 ;
        RECT 1777.970 1018.200 1778.290 1018.260 ;
        RECT 1822.220 1018.200 1822.360 1018.740 ;
        RECT 1823.970 1018.680 1824.290 1018.740 ;
        RECT 2152.870 1018.680 2153.190 1018.740 ;
        RECT 2297.310 1018.880 2297.630 1018.940 ;
        RECT 2388.390 1018.880 2388.710 1018.940 ;
        RECT 2297.310 1018.740 2388.710 1018.880 ;
        RECT 2297.310 1018.680 2297.630 1018.740 ;
        RECT 2388.390 1018.680 2388.710 1018.740 ;
        RECT 2304.210 1018.540 2304.530 1018.600 ;
        RECT 2363.090 1018.540 2363.410 1018.600 ;
        RECT 2304.210 1018.400 2363.410 1018.540 ;
        RECT 2304.210 1018.340 2304.530 1018.400 ;
        RECT 2363.090 1018.340 2363.410 1018.400 ;
        RECT 2369.990 1018.540 2370.310 1018.600 ;
        RECT 2428.870 1018.540 2429.190 1018.600 ;
        RECT 2369.990 1018.400 2429.190 1018.540 ;
        RECT 2369.990 1018.340 2370.310 1018.400 ;
        RECT 2428.870 1018.340 2429.190 1018.400 ;
        RECT 1777.970 1018.060 1822.360 1018.200 ;
        RECT 2259.590 1018.200 2259.910 1018.260 ;
        RECT 2307.890 1018.200 2308.210 1018.260 ;
        RECT 2355.730 1018.200 2356.050 1018.260 ;
        RECT 2259.590 1018.060 2356.050 1018.200 ;
        RECT 1766.010 1018.000 1766.330 1018.060 ;
        RECT 1777.970 1018.000 1778.290 1018.060 ;
        RECT 2259.590 1018.000 2259.910 1018.060 ;
        RECT 2307.890 1018.000 2308.210 1018.060 ;
        RECT 2355.730 1018.000 2356.050 1018.060 ;
        RECT 1748.070 1017.860 1748.390 1017.920 ;
        RECT 1787.630 1017.860 1787.950 1017.920 ;
        RECT 1748.070 1017.720 1787.950 1017.860 ;
        RECT 1748.070 1017.660 1748.390 1017.720 ;
        RECT 1787.630 1017.660 1787.950 1017.720 ;
        RECT 1822.130 1017.860 1822.450 1017.920 ;
        RECT 1869.510 1017.860 1869.830 1017.920 ;
        RECT 1822.130 1017.720 1869.830 1017.860 ;
        RECT 1822.130 1017.660 1822.450 1017.720 ;
        RECT 1869.510 1017.660 1869.830 1017.720 ;
        RECT 2273.390 1017.860 2273.710 1017.920 ;
        RECT 2317.090 1017.860 2317.410 1017.920 ;
        RECT 2353.890 1017.860 2354.210 1017.920 ;
        RECT 2373.210 1017.860 2373.530 1017.920 ;
        RECT 2273.390 1017.720 2354.210 1017.860 ;
        RECT 2273.390 1017.660 2273.710 1017.720 ;
        RECT 2317.090 1017.660 2317.410 1017.720 ;
        RECT 2353.890 1017.660 2354.210 1017.720 ;
        RECT 2354.440 1017.720 2373.530 1017.860 ;
        RECT 1782.110 1017.520 1782.430 1017.580 ;
        RECT 2228.770 1017.520 2229.090 1017.580 ;
        RECT 1747.700 1017.380 2229.090 1017.520 ;
        RECT 1782.110 1017.320 1782.430 1017.380 ;
        RECT 2228.770 1017.320 2229.090 1017.380 ;
        RECT 2283.510 1017.520 2283.830 1017.580 ;
        RECT 2323.530 1017.520 2323.850 1017.580 ;
        RECT 2354.440 1017.520 2354.580 1017.720 ;
        RECT 2373.210 1017.660 2373.530 1017.720 ;
        RECT 2373.670 1017.860 2373.990 1017.920 ;
        RECT 2408.170 1017.860 2408.490 1017.920 ;
        RECT 2373.670 1017.720 2408.490 1017.860 ;
        RECT 2373.670 1017.660 2373.990 1017.720 ;
        RECT 2408.170 1017.660 2408.490 1017.720 ;
        RECT 2283.510 1017.380 2354.580 1017.520 ;
        RECT 2358.030 1017.520 2358.350 1017.580 ;
        RECT 2377.810 1017.520 2378.130 1017.580 ;
        RECT 2421.970 1017.520 2422.290 1017.580 ;
        RECT 2358.030 1017.380 2422.290 1017.520 ;
        RECT 2283.510 1017.320 2283.830 1017.380 ;
        RECT 2323.530 1017.320 2323.850 1017.380 ;
        RECT 2358.030 1017.320 2358.350 1017.380 ;
        RECT 2377.810 1017.320 2378.130 1017.380 ;
        RECT 2421.970 1017.320 2422.290 1017.380 ;
        RECT 1748.070 1017.180 1748.390 1017.240 ;
        RECT 1790.390 1017.180 1790.710 1017.240 ;
        RECT 1654.690 1017.040 1713.340 1017.180 ;
        RECT 1713.660 1017.040 1746.920 1017.180 ;
        RECT 1747.240 1017.040 1790.710 1017.180 ;
        RECT 1654.690 1016.980 1655.010 1017.040 ;
        RECT 1700.690 1016.980 1701.010 1017.040 ;
        RECT 1675.390 1016.840 1675.710 1016.900 ;
        RECT 1713.660 1016.840 1713.800 1017.040 ;
        RECT 1718.170 1016.980 1718.490 1017.040 ;
        RECT 1746.780 1016.840 1746.920 1017.040 ;
        RECT 1748.070 1016.980 1748.390 1017.040 ;
        RECT 1790.390 1016.980 1790.710 1017.040 ;
        RECT 2303.290 1017.180 2303.610 1017.240 ;
        RECT 2346.990 1017.180 2347.310 1017.240 ;
        RECT 2387.930 1017.180 2388.250 1017.240 ;
        RECT 2303.290 1017.040 2388.250 1017.180 ;
        RECT 2303.290 1016.980 2303.610 1017.040 ;
        RECT 2346.990 1016.980 2347.310 1017.040 ;
        RECT 2387.930 1016.980 2388.250 1017.040 ;
        RECT 1766.010 1016.840 1766.330 1016.900 ;
        RECT 1675.390 1016.700 1713.800 1016.840 ;
        RECT 1714.120 1016.700 1746.460 1016.840 ;
        RECT 1746.780 1016.700 1766.330 1016.840 ;
        RECT 1675.390 1016.640 1675.710 1016.700 ;
        RECT 1662.050 1016.500 1662.370 1016.560 ;
        RECT 1707.130 1016.500 1707.450 1016.560 ;
        RECT 1714.120 1016.500 1714.260 1016.700 ;
        RECT 1662.050 1016.360 1714.260 1016.500 ;
        RECT 1714.490 1016.500 1714.810 1016.560 ;
        RECT 1745.770 1016.500 1746.090 1016.560 ;
        RECT 1714.490 1016.360 1746.090 1016.500 ;
        RECT 1746.320 1016.500 1746.460 1016.700 ;
        RECT 1766.010 1016.640 1766.330 1016.700 ;
        RECT 2293.630 1016.840 2293.950 1016.900 ;
        RECT 2342.390 1016.840 2342.710 1016.900 ;
        RECT 2387.470 1016.840 2387.790 1016.900 ;
        RECT 2293.630 1016.700 2387.790 1016.840 ;
        RECT 2293.630 1016.640 2293.950 1016.700 ;
        RECT 2342.390 1016.640 2342.710 1016.700 ;
        RECT 2387.470 1016.640 2387.790 1016.700 ;
        RECT 2281.210 1016.500 2281.530 1016.560 ;
        RECT 2329.510 1016.500 2329.830 1016.560 ;
        RECT 2358.030 1016.500 2358.350 1016.560 ;
        RECT 1746.320 1016.360 1756.120 1016.500 ;
        RECT 1662.050 1016.300 1662.370 1016.360 ;
        RECT 1707.130 1016.300 1707.450 1016.360 ;
        RECT 1714.490 1016.300 1714.810 1016.360 ;
        RECT 1745.770 1016.300 1746.090 1016.360 ;
        RECT 1755.980 1016.220 1756.120 1016.360 ;
        RECT 2281.210 1016.360 2358.350 1016.500 ;
        RECT 2281.210 1016.300 2281.530 1016.360 ;
        RECT 2329.510 1016.300 2329.830 1016.360 ;
        RECT 2358.030 1016.300 2358.350 1016.360 ;
        RECT 2363.550 1016.500 2363.870 1016.560 ;
        RECT 2373.670 1016.500 2373.990 1016.560 ;
        RECT 2363.550 1016.360 2373.990 1016.500 ;
        RECT 2363.550 1016.300 2363.870 1016.360 ;
        RECT 2373.670 1016.300 2373.990 1016.360 ;
        RECT 1668.950 1016.160 1669.270 1016.220 ;
        RECT 1713.570 1016.160 1713.890 1016.220 ;
        RECT 1717.710 1016.160 1718.030 1016.220 ;
        RECT 1668.950 1016.020 1718.030 1016.160 ;
        RECT 1668.950 1015.960 1669.270 1016.020 ;
        RECT 1713.570 1015.960 1713.890 1016.020 ;
        RECT 1717.710 1015.960 1718.030 1016.020 ;
        RECT 1721.390 1016.160 1721.710 1016.220 ;
        RECT 1755.430 1016.160 1755.750 1016.220 ;
        RECT 1721.390 1016.020 1755.750 1016.160 ;
        RECT 1721.390 1015.960 1721.710 1016.020 ;
        RECT 1755.430 1015.960 1755.750 1016.020 ;
        RECT 1755.890 1016.160 1756.210 1016.220 ;
        RECT 1800.050 1016.160 1800.370 1016.220 ;
        RECT 1755.890 1016.020 1800.370 1016.160 ;
        RECT 1755.890 1015.960 1756.210 1016.020 ;
        RECT 1800.050 1015.960 1800.370 1016.020 ;
        RECT 2287.190 1016.160 2287.510 1016.220 ;
        RECT 2335.490 1016.160 2335.810 1016.220 ;
        RECT 2380.570 1016.160 2380.890 1016.220 ;
        RECT 2287.190 1016.020 2380.890 1016.160 ;
        RECT 2287.190 1015.960 2287.510 1016.020 ;
        RECT 2335.490 1015.960 2335.810 1016.020 ;
        RECT 2380.570 1015.960 2380.890 1016.020 ;
        RECT 2381.030 1016.160 2381.350 1016.220 ;
        RECT 2381.030 1016.020 2395.060 1016.160 ;
        RECT 2381.030 1015.960 2381.350 1016.020 ;
        RECT 1683.210 1015.820 1683.530 1015.880 ;
        RECT 1729.670 1015.820 1729.990 1015.880 ;
        RECT 1777.970 1015.820 1778.290 1015.880 ;
        RECT 1683.210 1015.680 1778.290 1015.820 ;
        RECT 1683.210 1015.620 1683.530 1015.680 ;
        RECT 1729.670 1015.620 1729.990 1015.680 ;
        RECT 1777.970 1015.620 1778.290 1015.680 ;
        RECT 2312.030 1015.820 2312.350 1015.880 ;
        RECT 2355.270 1015.820 2355.590 1015.880 ;
        RECT 2312.030 1015.680 2355.590 1015.820 ;
        RECT 2312.030 1015.620 2312.350 1015.680 ;
        RECT 2355.270 1015.620 2355.590 1015.680 ;
        RECT 2355.730 1015.820 2356.050 1015.880 ;
        RECT 2394.370 1015.820 2394.690 1015.880 ;
        RECT 2355.730 1015.680 2394.690 1015.820 ;
        RECT 2394.920 1015.820 2395.060 1016.020 ;
        RECT 2402.190 1015.820 2402.510 1015.880 ;
        RECT 2394.920 1015.680 2402.510 1015.820 ;
        RECT 2355.730 1015.620 2356.050 1015.680 ;
        RECT 2394.370 1015.620 2394.690 1015.680 ;
        RECT 2402.190 1015.620 2402.510 1015.680 ;
        RECT 1648.710 1015.480 1649.030 1015.540 ;
        RECT 1696.090 1015.480 1696.410 1015.540 ;
        RECT 1717.250 1015.480 1717.570 1015.540 ;
        RECT 1648.710 1015.340 1717.570 1015.480 ;
        RECT 1648.710 1015.280 1649.030 1015.340 ;
        RECT 1696.090 1015.280 1696.410 1015.340 ;
        RECT 1717.250 1015.280 1717.570 1015.340 ;
        RECT 1717.710 1015.480 1718.030 1015.540 ;
        RECT 1759.110 1015.480 1759.430 1015.540 ;
        RECT 1717.710 1015.340 1759.430 1015.480 ;
        RECT 1717.710 1015.280 1718.030 1015.340 ;
        RECT 1759.110 1015.280 1759.430 1015.340 ;
        RECT 2254.990 1015.480 2255.310 1015.540 ;
        RECT 2559.970 1015.480 2560.290 1015.540 ;
        RECT 2254.990 1015.340 2560.290 1015.480 ;
        RECT 2254.990 1015.280 2255.310 1015.340 ;
        RECT 2559.970 1015.280 2560.290 1015.340 ;
        RECT 1683.210 1015.140 1683.530 1015.200 ;
        RECT 1724.610 1015.140 1724.930 1015.200 ;
        RECT 1772.910 1015.140 1773.230 1015.200 ;
        RECT 1683.210 1015.000 1773.230 1015.140 ;
        RECT 1683.210 1014.940 1683.530 1015.000 ;
        RECT 1724.610 1014.940 1724.930 1015.000 ;
        RECT 1772.910 1014.940 1773.230 1015.000 ;
        RECT 2249.010 1015.140 2249.330 1015.200 ;
        RECT 2566.870 1015.140 2567.190 1015.200 ;
        RECT 2249.010 1015.000 2567.190 1015.140 ;
        RECT 2249.010 1014.940 2249.330 1015.000 ;
        RECT 2566.870 1014.940 2567.190 1015.000 ;
        RECT 1483.110 1014.800 1483.430 1014.860 ;
        RECT 1787.170 1014.800 1787.490 1014.860 ;
        RECT 1483.110 1014.660 1787.490 1014.800 ;
        RECT 1483.110 1014.600 1483.430 1014.660 ;
        RECT 1787.170 1014.600 1787.490 1014.660 ;
        RECT 2345.610 1014.800 2345.930 1014.860 ;
        RECT 2366.770 1014.800 2367.090 1014.860 ;
        RECT 2345.610 1014.660 2367.090 1014.800 ;
        RECT 2345.610 1014.600 2345.930 1014.660 ;
        RECT 2366.770 1014.600 2367.090 1014.660 ;
        RECT 2373.210 1014.800 2373.530 1014.860 ;
        RECT 2415.070 1014.800 2415.390 1014.860 ;
        RECT 2373.210 1014.660 2415.390 1014.800 ;
        RECT 2373.210 1014.600 2373.530 1014.660 ;
        RECT 2415.070 1014.600 2415.390 1014.660 ;
        RECT 1476.210 1014.460 1476.530 1014.520 ;
        RECT 1794.070 1014.460 1794.390 1014.520 ;
        RECT 1476.210 1014.320 1794.390 1014.460 ;
        RECT 1476.210 1014.260 1476.530 1014.320 ;
        RECT 1794.070 1014.260 1794.390 1014.320 ;
        RECT 2262.810 1014.460 2263.130 1014.520 ;
        RECT 2546.170 1014.460 2546.490 1014.520 ;
        RECT 2262.810 1014.320 2546.490 1014.460 ;
        RECT 2262.810 1014.260 2263.130 1014.320 ;
        RECT 2546.170 1014.260 2546.490 1014.320 ;
        RECT 1945.410 1007.320 1945.730 1007.380 ;
        RECT 2498.790 1007.320 2499.110 1007.380 ;
        RECT 1945.410 1007.180 2499.110 1007.320 ;
        RECT 1945.410 1007.120 1945.730 1007.180 ;
        RECT 2498.790 1007.120 2499.110 1007.180 ;
        RECT 1938.510 1006.980 1938.830 1007.040 ;
        RECT 2499.250 1006.980 2499.570 1007.040 ;
        RECT 1938.510 1006.840 2499.570 1006.980 ;
        RECT 1938.510 1006.780 1938.830 1006.840 ;
        RECT 2499.250 1006.780 2499.570 1006.840 ;
        RECT 1924.710 1006.640 1925.030 1006.700 ;
        RECT 2499.710 1006.640 2500.030 1006.700 ;
        RECT 1924.710 1006.500 2500.030 1006.640 ;
        RECT 1924.710 1006.440 1925.030 1006.500 ;
        RECT 2499.710 1006.440 2500.030 1006.500 ;
        RECT 1917.810 1006.300 1918.130 1006.360 ;
        RECT 2500.170 1006.300 2500.490 1006.360 ;
        RECT 1917.810 1006.160 2500.490 1006.300 ;
        RECT 1917.810 1006.100 1918.130 1006.160 ;
        RECT 2500.170 1006.100 2500.490 1006.160 ;
        RECT 1904.010 1005.960 1904.330 1006.020 ;
        RECT 2500.630 1005.960 2500.950 1006.020 ;
        RECT 1904.010 1005.820 2500.950 1005.960 ;
        RECT 1904.010 1005.760 1904.330 1005.820 ;
        RECT 2500.630 1005.760 2500.950 1005.820 ;
        RECT 1959.210 1003.580 1959.530 1003.640 ;
        RECT 2498.330 1003.580 2498.650 1003.640 ;
        RECT 1959.210 1003.440 2498.650 1003.580 ;
        RECT 1959.210 1003.380 1959.530 1003.440 ;
        RECT 2498.330 1003.380 2498.650 1003.440 ;
        RECT 2287.650 1003.240 2287.970 1003.300 ;
        RECT 2497.870 1003.240 2498.190 1003.300 ;
        RECT 2287.650 1003.100 2498.190 1003.240 ;
        RECT 2287.650 1003.040 2287.970 1003.100 ;
        RECT 2497.870 1003.040 2498.190 1003.100 ;
        RECT 2093.990 1001.540 2094.310 1001.600 ;
        RECT 2587.570 1001.540 2587.890 1001.600 ;
        RECT 2093.990 1001.400 2587.890 1001.540 ;
        RECT 2093.990 1001.340 2094.310 1001.400 ;
        RECT 2587.570 1001.340 2587.890 1001.400 ;
      LAYER met1 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
      LAYER met1 ;
        RECT 1898.950 917.560 1899.270 917.620 ;
        RECT 2093.990 917.560 2094.310 917.620 ;
        RECT 1898.950 917.420 2094.310 917.560 ;
        RECT 1898.950 917.360 1899.270 917.420 ;
        RECT 2093.990 917.360 2094.310 917.420 ;
        RECT 1899.870 620.740 1900.190 620.800 ;
        RECT 1976.690 620.740 1977.010 620.800 ;
        RECT 1899.870 620.600 1977.010 620.740 ;
        RECT 1899.870 620.540 1900.190 620.600 ;
        RECT 1976.690 620.540 1977.010 620.600 ;
        RECT 1900.330 593.200 1900.650 593.260 ;
        RECT 1969.790 593.200 1970.110 593.260 ;
        RECT 1900.330 593.060 1970.110 593.200 ;
        RECT 1900.330 593.000 1900.650 593.060 ;
        RECT 1969.790 593.000 1970.110 593.060 ;
        RECT 1900.330 579.600 1900.650 579.660 ;
        RECT 1997.390 579.600 1997.710 579.660 ;
        RECT 1900.330 579.460 1997.710 579.600 ;
        RECT 1900.330 579.400 1900.650 579.460 ;
        RECT 1997.390 579.400 1997.710 579.460 ;
      LAYER met1 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met1 ;
        RECT 2504.310 917.560 2504.630 917.620 ;
        RECT 2587.570 917.560 2587.890 917.620 ;
        RECT 2504.310 917.420 2587.890 917.560 ;
        RECT 2504.310 917.360 2504.630 917.420 ;
        RECT 2587.570 917.360 2587.890 917.420 ;
        RECT 1503.810 554.780 1504.130 554.840 ;
        RECT 2083.870 554.780 2084.190 554.840 ;
        RECT 1503.810 554.640 2084.190 554.780 ;
        RECT 1503.810 554.580 1504.130 554.640 ;
        RECT 2083.870 554.580 2084.190 554.640 ;
      LAYER via ;
        RECT 2442.700 3066.840 2442.960 3067.100 ;
        RECT 2469.840 3066.840 2470.100 3067.100 ;
        RECT 1868.160 3063.780 1868.420 3064.040 ;
        RECT 1898.060 3063.780 1898.320 3064.040 ;
        RECT 2442.700 3063.780 2442.960 3064.040 ;
        RECT 2469.840 3063.780 2470.100 3064.040 ;
        RECT 2497.900 3063.780 2498.160 3064.040 ;
        RECT 1899.900 3051.880 1900.160 3052.140 ;
        RECT 2482.260 3051.880 2482.520 3052.140 ;
        RECT 2048.940 2697.940 2049.200 2698.200 ;
        RECT 2083.900 2697.940 2084.160 2698.200 ;
        RECT 1486.360 2604.440 1486.620 2604.700 ;
        RECT 2090.340 2604.440 2090.600 2604.700 ;
        RECT 1614.700 2594.240 1614.960 2594.500 ;
        RECT 1661.620 2594.240 1661.880 2594.500 ;
        RECT 1537.880 2593.900 1538.140 2594.160 ;
        RECT 1621.600 2593.900 1621.860 2594.160 ;
        RECT 1656.100 2593.900 1656.360 2594.160 ;
        RECT 1702.560 2593.900 1702.820 2594.160 ;
        RECT 1586.640 2593.560 1586.900 2593.820 ;
        RECT 1626.660 2593.560 1626.920 2593.820 ;
        RECT 1669.900 2593.560 1670.160 2593.820 ;
        RECT 1690.600 2593.560 1690.860 2593.820 ;
        RECT 1738.440 2593.560 1738.700 2593.820 ;
        RECT 2256.400 2593.560 2256.660 2593.820 ;
        RECT 2297.800 2593.560 2298.060 2593.820 ;
        RECT 1598.600 2593.220 1598.860 2593.480 ;
        RECT 1644.600 2593.220 1644.860 2593.480 ;
        RECT 1651.040 2593.220 1651.300 2593.480 ;
        RECT 1697.960 2593.220 1698.220 2593.480 ;
        RECT 1743.960 2593.220 1744.220 2593.480 ;
        RECT 2215.920 2593.220 2216.180 2593.480 ;
        RECT 2262.840 2593.220 2263.100 2593.480 ;
        RECT 2305.160 2593.220 2305.420 2593.480 ;
        RECT 1476.240 2592.880 1476.500 2593.140 ;
        RECT 1587.100 2592.880 1587.360 2593.140 ;
        RECT 1604.120 2592.880 1604.380 2593.140 ;
        RECT 1661.620 2592.880 1661.880 2593.140 ;
        RECT 1707.620 2592.880 1707.880 2593.140 ;
        RECT 1569.620 2592.540 1569.880 2592.800 ;
        RECT 1573.760 2592.200 1574.020 2592.460 ;
        RECT 1591.240 2592.540 1591.500 2592.800 ;
        RECT 1639.080 2592.540 1639.340 2592.800 ;
        RECT 1685.080 2592.540 1685.340 2592.800 ;
        RECT 1686.460 2592.540 1686.720 2592.800 ;
        RECT 1732.920 2592.880 1733.180 2593.140 ;
        RECT 2208.100 2592.880 2208.360 2593.140 ;
        RECT 2220.520 2592.880 2220.780 2593.140 ;
        RECT 2268.360 2592.880 2268.620 2593.140 ;
        RECT 2311.600 2592.880 2311.860 2593.140 ;
        RECT 1738.440 2592.540 1738.700 2592.800 ;
        RECT 2215.000 2592.540 2215.260 2592.800 ;
        RECT 2243.980 2592.540 2244.240 2592.800 ;
        RECT 2291.820 2592.540 2292.080 2592.800 ;
        RECT 2332.300 2592.540 2332.560 2592.800 ;
        RECT 1462.440 2591.860 1462.700 2592.120 ;
        RECT 1581.120 2591.860 1581.380 2592.120 ;
        RECT 1448.640 2591.520 1448.900 2591.780 ;
        RECT 1573.300 2591.520 1573.560 2591.780 ;
        RECT 1614.700 2592.200 1614.960 2592.460 ;
        RECT 1630.800 2592.200 1631.060 2592.460 ;
        RECT 1633.560 2592.200 1633.820 2592.460 ;
        RECT 1679.560 2592.200 1679.820 2592.460 ;
        RECT 1725.560 2592.200 1725.820 2592.460 ;
        RECT 1731.540 2592.200 1731.800 2592.460 ;
        RECT 1743.960 2592.200 1744.220 2592.460 ;
        RECT 2228.800 2592.200 2229.060 2592.460 ;
        RECT 2249.500 2592.200 2249.760 2592.460 ;
        RECT 1644.600 2591.860 1644.860 2592.120 ;
        RECT 1690.600 2591.860 1690.860 2592.120 ;
        RECT 1993.280 2591.860 1993.540 2592.120 ;
        RECT 2152.900 2591.860 2153.160 2592.120 ;
        RECT 2235.700 2591.860 2235.960 2592.120 ;
        RECT 2285.380 2591.860 2285.640 2592.120 ;
        RECT 2297.800 2591.860 2298.060 2592.120 ;
        RECT 2339.200 2591.860 2339.460 2592.120 ;
        RECT 1621.600 2591.520 1621.860 2591.780 ;
        RECT 1667.140 2591.520 1667.400 2591.780 ;
        RECT 1713.140 2591.520 1713.400 2591.780 ;
        RECT 1979.940 2591.520 1980.200 2591.780 ;
        RECT 2146.460 2591.520 2146.720 2591.780 ;
        RECT 2232.940 2591.520 2233.200 2591.780 ;
        RECT 2280.320 2591.520 2280.580 2591.780 ;
        RECT 2332.300 2591.520 2332.560 2591.780 ;
        RECT 1565.480 2591.180 1565.740 2591.440 ;
        RECT 1608.260 2591.180 1608.520 2591.440 ;
        RECT 1656.100 2591.180 1656.360 2591.440 ;
        RECT 1669.900 2591.180 1670.160 2591.440 ;
        RECT 1718.200 2591.180 1718.460 2591.440 ;
        RECT 1966.140 2591.180 1966.400 2591.440 ;
        RECT 2146.000 2591.180 2146.260 2591.440 ;
        RECT 2276.180 2591.180 2276.440 2591.440 ;
        RECT 2318.500 2591.180 2318.760 2591.440 ;
        RECT 2214.540 2590.840 2214.800 2591.100 ;
        RECT 2256.400 2590.840 2256.660 2591.100 ;
        RECT 2280.320 2590.840 2280.580 2591.100 ;
        RECT 2325.400 2590.840 2325.660 2591.100 ;
        RECT 1517.640 2590.500 1517.900 2590.760 ;
        RECT 1607.800 2590.500 1608.060 2590.760 ;
        RECT 1959.240 2590.500 1959.500 2590.760 ;
        RECT 2126.680 2590.500 2126.940 2590.760 ;
        RECT 1531.440 2590.160 1531.700 2590.420 ;
        RECT 1614.700 2590.160 1614.960 2590.420 ;
        RECT 1779.840 2590.160 1780.100 2590.420 ;
        RECT 2132.200 2590.160 2132.460 2590.420 ;
        RECT 2179.580 2590.160 2179.840 2590.420 ;
        RECT 2220.520 2590.160 2220.780 2590.420 ;
        RECT 1496.940 2589.820 1497.200 2590.080 ;
        RECT 1594.000 2589.820 1594.260 2590.080 ;
        RECT 1702.560 2589.820 1702.820 2590.080 ;
        RECT 2152.900 2589.820 2153.160 2590.080 ;
        RECT 2183.720 2589.820 2183.980 2590.080 ;
        RECT 2227.880 2589.820 2228.140 2590.080 ;
        RECT 2276.180 2589.820 2276.440 2590.080 ;
        RECT 1483.140 2589.480 1483.400 2589.740 ;
        RECT 1587.100 2589.480 1587.360 2589.740 ;
        RECT 1614.240 2589.480 1614.500 2589.740 ;
        RECT 1663.000 2589.480 1663.260 2589.740 ;
        RECT 1707.620 2589.480 1707.880 2589.740 ;
        RECT 2159.800 2589.480 2160.060 2589.740 ;
        RECT 2170.380 2589.480 2170.640 2589.740 ;
        RECT 2215.920 2589.480 2216.180 2589.740 ;
        RECT 1586.640 2589.140 1586.900 2589.400 ;
        RECT 1642.300 2589.140 1642.560 2589.400 ;
        RECT 1652.420 2589.140 1652.680 2589.400 ;
        RECT 1678.640 2589.140 1678.900 2589.400 ;
        RECT 1718.200 2589.140 1718.460 2589.400 ;
        RECT 2180.500 2589.140 2180.760 2589.400 ;
        RECT 2184.640 2589.140 2184.900 2589.400 ;
        RECT 2186.480 2589.140 2186.740 2589.400 ;
        RECT 2232.940 2589.140 2233.200 2589.400 ;
        RECT 1503.380 2588.800 1503.640 2589.060 ;
        RECT 1600.900 2588.800 1601.160 2589.060 ;
        RECT 1607.340 2588.800 1607.600 2589.060 ;
        RECT 1656.100 2588.800 1656.360 2589.060 ;
        RECT 2163.020 2588.800 2163.280 2589.060 ;
        RECT 2209.480 2588.800 2209.740 2589.060 ;
        RECT 2214.540 2588.800 2214.800 2589.060 ;
        RECT 1558.580 2588.460 1558.840 2588.720 ;
        RECT 1631.260 2588.460 1631.520 2588.720 ;
        RECT 1669.440 2588.460 1669.700 2588.720 ;
        RECT 1690.600 2588.460 1690.860 2588.720 ;
        RECT 2190.620 2588.460 2190.880 2588.720 ;
        RECT 2235.700 2588.460 2235.960 2588.720 ;
        RECT 1551.680 2588.120 1551.940 2588.380 ;
        RECT 1621.600 2588.120 1621.860 2588.380 ;
        RECT 1641.840 2588.120 1642.100 2588.380 ;
        RECT 1669.900 2588.120 1670.160 2588.380 ;
        RECT 1731.540 2588.120 1731.800 2588.380 ;
        RECT 2194.300 2588.120 2194.560 2588.380 ;
        RECT 2204.420 2588.120 2204.680 2588.380 ;
        RECT 2249.500 2588.120 2249.760 2588.380 ;
        RECT 1441.740 2587.780 1442.000 2588.040 ;
        RECT 1566.400 2587.780 1566.660 2588.040 ;
        RECT 1586.180 2587.780 1586.440 2588.040 ;
        RECT 1630.800 2587.780 1631.060 2588.040 ;
        RECT 1427.940 2587.440 1428.200 2587.700 ;
        RECT 1559.500 2587.440 1559.760 2587.700 ;
        RECT 1572.840 2587.440 1573.100 2587.700 ;
        RECT 1635.400 2587.780 1635.660 2588.040 ;
        RECT 1638.620 2587.780 1638.880 2588.040 ;
        RECT 1663.000 2587.780 1663.260 2588.040 ;
        RECT 1713.140 2587.780 1713.400 2588.040 ;
        RECT 2173.600 2587.780 2173.860 2588.040 ;
        RECT 2197.520 2587.780 2197.780 2588.040 ;
        RECT 2243.980 2587.780 2244.240 2588.040 ;
        RECT 1631.720 2587.440 1631.980 2587.700 ;
        RECT 1649.200 2587.440 1649.460 2587.700 ;
        RECT 1666.220 2587.440 1666.480 2587.700 ;
        RECT 1683.700 2587.440 1683.960 2587.700 ;
        RECT 1686.920 2587.440 1687.180 2587.700 ;
        RECT 1697.500 2587.440 1697.760 2587.700 ;
        RECT 1736.600 2587.440 1736.860 2587.700 ;
        RECT 1742.120 2587.440 1742.380 2587.700 ;
        RECT 2169.000 2511.620 2169.260 2511.880 ;
        RECT 2170.380 2511.620 2170.640 2511.880 ;
        RECT 2168.080 2463.000 2168.340 2463.260 ;
        RECT 2169.460 2463.000 2169.720 2463.260 ;
        RECT 1487.740 2414.720 1488.000 2414.980 ;
        RECT 1887.940 2414.720 1888.200 2414.980 ;
        RECT 2166.240 2414.720 2166.500 2414.980 ;
        RECT 2240.300 2414.720 2240.560 2414.980 ;
        RECT 2276.640 2414.720 2276.900 2414.980 ;
        RECT 2449.600 2414.720 2449.860 2414.980 ;
        RECT 1488.200 2414.380 1488.460 2414.640 ;
        RECT 1898.980 2414.380 1899.240 2414.640 ;
        RECT 2133.120 2414.380 2133.380 2414.640 ;
        RECT 2197.520 2414.380 2197.780 2414.640 ;
        RECT 2283.540 2414.380 2283.800 2414.640 ;
        RECT 2460.180 2414.380 2460.440 2414.640 ;
        RECT 1488.660 2414.040 1488.920 2414.300 ;
        RECT 1911.400 2414.040 1911.660 2414.300 ;
        RECT 2173.140 2414.040 2173.400 2414.300 ;
        RECT 2251.340 2414.040 2251.600 2414.300 ;
        RECT 2290.440 2414.040 2290.700 2414.300 ;
        RECT 2471.220 2414.040 2471.480 2414.300 ;
        RECT 1489.120 2413.700 1489.380 2413.960 ;
        RECT 1920.600 2413.700 1920.860 2413.960 ;
        RECT 2180.500 2413.700 2180.760 2413.960 ;
        RECT 2183.720 2413.700 2183.980 2413.960 ;
        RECT 2186.940 2413.700 2187.200 2413.960 ;
        RECT 2272.960 2413.700 2273.220 2413.960 ;
        RECT 2297.340 2413.700 2297.600 2413.960 ;
        RECT 2482.260 2413.700 2482.520 2413.960 ;
        RECT 1489.580 2413.360 1489.840 2413.620 ;
        RECT 1932.100 2413.360 1932.360 2413.620 ;
        RECT 1956.940 2413.360 1957.200 2413.620 ;
        RECT 1959.240 2413.360 1959.500 2413.620 ;
        RECT 1990.060 2413.360 1990.320 2413.620 ;
        RECT 1993.280 2413.360 1993.540 2413.620 ;
        RECT 2180.040 2413.360 2180.300 2413.620 ;
        RECT 2263.300 2413.360 2263.560 2413.620 ;
        RECT 2303.780 2413.360 2304.040 2413.620 ;
        RECT 2493.300 2413.360 2493.560 2413.620 ;
        RECT 1545.240 2413.020 1545.500 2413.280 ;
        RECT 1997.880 2413.020 1998.140 2413.280 ;
        RECT 2122.080 2413.020 2122.340 2413.280 ;
        RECT 2190.620 2413.020 2190.880 2413.280 ;
        RECT 2193.840 2413.020 2194.100 2413.280 ;
        RECT 2284.460 2413.020 2284.720 2413.280 ;
        RECT 2311.140 2413.020 2311.400 2413.280 ;
        RECT 2515.380 2413.020 2515.640 2413.280 ;
        RECT 1439.440 2412.680 1439.700 2412.940 ;
        RECT 1441.740 2412.680 1442.000 2412.940 ;
        RECT 1494.640 2412.680 1494.900 2412.940 ;
        RECT 1496.940 2412.680 1497.200 2412.940 ;
        RECT 1527.760 2412.680 1528.020 2412.940 ;
        RECT 1531.440 2412.680 1531.700 2412.940 ;
        RECT 1551.220 2412.680 1551.480 2412.940 ;
        RECT 2008.920 2412.680 2009.180 2412.940 ;
        RECT 2045.260 2412.680 2045.520 2412.940 ;
        RECT 2048.940 2412.680 2049.200 2412.940 ;
        RECT 2111.040 2412.680 2111.300 2412.940 ;
        RECT 2184.640 2412.680 2184.900 2412.940 ;
        RECT 2193.380 2412.680 2193.640 2412.940 ;
        RECT 2295.040 2412.680 2295.300 2412.940 ;
        RECT 2304.240 2412.680 2304.500 2412.940 ;
        RECT 2504.800 2412.680 2505.060 2412.940 ;
        RECT 1552.140 2412.340 1552.400 2412.600 ;
        RECT 2019.960 2412.340 2020.220 2412.600 ;
        RECT 2100.000 2412.340 2100.260 2412.600 ;
        RECT 2180.500 2412.340 2180.760 2412.600 ;
        RECT 2214.540 2412.340 2214.800 2412.600 ;
        RECT 1559.040 2412.000 1559.300 2412.260 ;
        RECT 2031.000 2412.000 2031.260 2412.260 ;
        RECT 2086.660 2412.000 2086.920 2412.260 ;
        RECT 2176.820 2412.000 2177.080 2412.260 ;
        RECT 2200.740 2412.000 2201.000 2412.260 ;
        RECT 2306.080 2412.000 2306.340 2412.260 ;
        RECT 1406.780 2411.660 1407.040 2411.920 ;
        RECT 1898.060 2411.660 1898.320 2411.920 ;
        RECT 2076.080 2411.660 2076.340 2411.920 ;
        RECT 2169.000 2411.660 2169.260 2411.920 ;
        RECT 2207.640 2411.660 2207.900 2411.920 ;
        RECT 2318.500 2411.660 2318.760 2411.920 ;
        RECT 2324.940 2412.340 2325.200 2412.600 ;
        RECT 2537.460 2412.340 2537.720 2412.600 ;
        RECT 2319.420 2412.000 2319.680 2412.260 ;
        RECT 2526.420 2412.000 2526.680 2412.260 ;
        RECT 2328.160 2411.660 2328.420 2411.920 ;
        RECT 2331.840 2411.660 2332.100 2411.920 ;
        RECT 2548.500 2411.660 2548.760 2411.920 ;
        RECT 1511.660 2411.320 1511.920 2411.580 ;
        RECT 1559.500 2411.320 1559.760 2411.580 ;
        RECT 1609.640 2411.320 1609.900 2411.580 ;
        RECT 1656.100 2411.320 1656.360 2411.580 ;
        RECT 1703.020 2411.320 1703.280 2411.580 ;
        RECT 1752.700 2411.320 1752.960 2411.580 ;
        RECT 1800.540 2411.320 1800.800 2411.580 ;
        RECT 1835.500 2411.320 1835.760 2411.580 ;
        RECT 1487.280 2410.980 1487.540 2411.240 ;
        RECT 1510.740 2410.980 1511.000 2411.240 ;
        RECT 1511.200 2410.980 1511.460 2411.240 ;
        RECT 1703.480 2410.980 1703.740 2411.240 ;
        RECT 1714.060 2410.980 1714.320 2411.240 ;
        RECT 1876.900 2410.980 1877.160 2411.240 ;
        RECT 1877.360 2410.980 1877.620 2411.240 ;
        RECT 1932.560 2411.320 1932.820 2411.580 ;
        RECT 1945.900 2411.320 1946.160 2411.580 ;
        RECT 2067.340 2411.320 2067.600 2411.580 ;
        RECT 2163.020 2411.320 2163.280 2411.580 ;
        RECT 2221.440 2411.320 2221.700 2411.580 ;
        RECT 2340.120 2411.320 2340.380 2411.580 ;
        RECT 2345.180 2411.320 2345.440 2411.580 ;
        RECT 2570.580 2411.320 2570.840 2411.580 ;
        RECT 1486.820 2410.640 1487.080 2410.900 ;
        RECT 1510.280 2410.640 1510.540 2410.900 ;
        RECT 1538.340 2410.640 1538.600 2410.900 ;
        RECT 1865.860 2410.640 1866.120 2410.900 ;
        RECT 2144.160 2410.980 2144.420 2411.240 ;
        RECT 2204.420 2410.980 2204.680 2411.240 ;
        RECT 2269.740 2410.980 2270.000 2411.240 ;
        RECT 2438.100 2410.980 2438.360 2411.240 ;
        RECT 2053.080 2410.640 2053.340 2410.900 ;
        RECT 2269.280 2410.640 2269.540 2410.900 ;
        RECT 2428.900 2410.640 2429.160 2410.900 ;
        RECT 1626.660 2410.300 1626.920 2410.560 ;
        RECT 1638.620 2410.300 1638.880 2410.560 ;
        RECT 1648.740 2410.300 1649.000 2410.560 ;
        RECT 1652.420 2410.300 1652.680 2410.560 ;
        RECT 1659.780 2410.300 1660.040 2410.560 ;
        RECT 1666.220 2410.300 1666.480 2410.560 ;
        RECT 1559.500 2409.960 1559.760 2410.220 ;
        RECT 1594.000 2409.960 1594.260 2410.220 ;
        RECT 1656.100 2409.960 1656.360 2410.220 ;
        RECT 1703.020 2410.300 1703.280 2410.560 ;
        RECT 1731.540 2410.300 1731.800 2410.560 ;
        RECT 1733.840 2410.300 1734.100 2410.560 ;
        RECT 1742.120 2410.300 1742.380 2410.560 ;
        RECT 1745.800 2410.300 1746.060 2410.560 ;
        RECT 1746.260 2410.300 1746.520 2410.560 ;
        RECT 1755.460 2410.300 1755.720 2410.560 ;
        RECT 1791.800 2410.300 1792.060 2410.560 ;
        RECT 2089.880 2410.300 2090.140 2410.560 ;
        RECT 2262.840 2410.300 2263.100 2410.560 ;
        RECT 2416.480 2410.300 2416.740 2410.560 ;
        RECT 1681.860 2409.960 1682.120 2410.220 ;
        RECT 1686.920 2409.960 1687.180 2410.220 ;
        RECT 1703.480 2409.960 1703.740 2410.220 ;
        RECT 1714.060 2409.960 1714.320 2410.220 ;
        RECT 1752.700 2409.960 1752.960 2410.220 ;
        RECT 1800.540 2409.960 1800.800 2410.220 ;
        RECT 1802.840 2409.960 1803.100 2410.220 ;
        RECT 2089.420 2409.960 2089.680 2410.220 ;
        RECT 2255.940 2409.960 2256.200 2410.220 ;
        RECT 2405.440 2409.960 2405.700 2410.220 ;
        RECT 1593.540 2409.620 1593.800 2409.880 ;
        RECT 1631.720 2409.620 1631.980 2409.880 ;
        RECT 1744.880 2409.620 1745.140 2409.880 ;
        RECT 1766.500 2409.620 1766.760 2409.880 ;
        RECT 1813.880 2409.620 1814.140 2409.880 ;
        RECT 2088.960 2409.620 2089.220 2409.880 ;
        RECT 2249.040 2409.620 2249.300 2409.880 ;
        RECT 2394.400 2409.620 2394.660 2409.880 ;
        RECT 1472.560 2409.280 1472.820 2409.540 ;
        RECT 1476.240 2409.280 1476.500 2409.540 ;
        RECT 1582.500 2409.280 1582.760 2409.540 ;
        RECT 1586.640 2409.280 1586.900 2409.540 ;
        RECT 1604.580 2409.280 1604.840 2409.540 ;
        RECT 1607.340 2409.280 1607.600 2409.540 ;
        RECT 1637.700 2409.280 1637.960 2409.540 ;
        RECT 1641.840 2409.280 1642.100 2409.540 ;
        RECT 1824.920 2409.280 1825.180 2409.540 ;
        RECT 2088.500 2409.280 2088.760 2409.540 ;
        RECT 2235.240 2409.280 2235.500 2409.540 ;
        RECT 2373.700 2409.280 2373.960 2409.540 ;
        RECT 1835.040 2408.940 1835.300 2409.200 ;
        RECT 2088.040 2408.940 2088.300 2409.200 ;
        RECT 2242.140 2408.940 2242.400 2409.200 ;
        RECT 2383.360 2408.940 2383.620 2409.200 ;
        RECT 1692.900 2408.600 1693.160 2408.860 ;
        RECT 1697.040 2408.600 1697.300 2408.860 ;
        RECT 1847.000 2408.600 1847.260 2408.860 ;
        RECT 2087.580 2408.600 2087.840 2408.860 ;
        RECT 2227.880 2408.600 2228.140 2408.860 ;
        RECT 2361.280 2408.600 2361.540 2408.860 ;
        RECT 1858.040 2408.260 1858.300 2408.520 ;
        RECT 2087.120 2408.260 2087.380 2408.520 ;
        RECT 2228.340 2408.260 2228.600 2408.520 ;
        RECT 2350.240 2408.260 2350.500 2408.520 ;
        RECT 2587.600 1196.840 2587.860 1197.100 ;
        RECT 2593.580 1196.840 2593.840 1197.100 ;
        RECT 1668.520 1193.440 1668.780 1193.700 ;
        RECT 1722.800 1193.440 1723.060 1193.700 ;
        RECT 2131.740 1193.440 2132.000 1193.700 ;
        RECT 2245.820 1193.440 2246.080 1193.700 ;
        RECT 2363.120 1193.440 2363.380 1193.700 ;
        RECT 2471.220 1193.440 2471.480 1193.700 ;
        RECT 1662.540 1193.100 1662.800 1193.360 ;
        RECT 1733.840 1193.100 1734.100 1193.360 ;
        RECT 2122.080 1193.100 2122.340 1193.360 ;
        RECT 2252.720 1193.100 2252.980 1193.360 ;
        RECT 2276.180 1193.100 2276.440 1193.360 ;
        RECT 2383.820 1193.100 2384.080 1193.360 ;
        RECT 1655.640 1192.760 1655.900 1193.020 ;
        RECT 1745.800 1192.760 1746.060 1193.020 ;
        RECT 1969.820 1192.760 1970.080 1193.020 ;
        RECT 2031.000 1192.760 2031.260 1193.020 ;
        RECT 2111.040 1192.760 2111.300 1193.020 ;
        RECT 2259.620 1192.760 2259.880 1193.020 ;
        RECT 2287.220 1192.760 2287.480 1193.020 ;
        RECT 2290.440 1192.760 2290.700 1193.020 ;
        RECT 1582.500 1192.420 1582.760 1192.680 ;
        RECT 1586.640 1192.420 1586.900 1192.680 ;
        RECT 1667.600 1192.420 1667.860 1192.680 ;
        RECT 1755.460 1192.420 1755.720 1192.680 ;
        RECT 1902.200 1192.420 1902.460 1192.680 ;
        RECT 1997.880 1192.420 1998.140 1192.680 ;
        RECT 2100.000 1192.420 2100.260 1192.680 ;
        RECT 1472.560 1192.080 1472.820 1192.340 ;
        RECT 1476.240 1192.080 1476.500 1192.340 ;
        RECT 1641.380 1192.080 1641.640 1192.340 ;
        RECT 1766.500 1192.080 1766.760 1192.340 ;
        RECT 1901.740 1192.080 1902.000 1192.340 ;
        RECT 2008.920 1192.080 2009.180 1192.340 ;
        RECT 2076.540 1192.080 2076.800 1192.340 ;
        RECT 2265.140 1192.420 2265.400 1192.680 ;
        RECT 2384.280 1192.760 2384.540 1193.020 ;
        RECT 2317.580 1192.420 2317.840 1192.680 ;
        RECT 2449.600 1192.420 2449.860 1192.680 ;
        RECT 1559.040 1191.740 1559.300 1192.000 ;
        RECT 1714.520 1191.740 1714.780 1192.000 ;
        RECT 1901.280 1191.740 1901.540 1192.000 ;
        RECT 2019.960 1191.740 2020.220 1192.000 ;
        RECT 2067.340 1191.740 2067.600 1192.000 ;
        RECT 2260.540 1191.740 2260.800 1192.000 ;
        RECT 2266.520 1192.080 2266.780 1192.340 ;
        RECT 2311.140 1192.080 2311.400 1192.340 ;
        RECT 2460.180 1192.080 2460.440 1192.340 ;
        RECT 2280.320 1191.740 2280.580 1192.000 ;
        RECT 2283.540 1191.740 2283.800 1192.000 ;
        RECT 2504.800 1191.740 2505.060 1192.000 ;
        RECT 1549.840 1191.400 1550.100 1191.660 ;
        RECT 1721.420 1191.400 1721.680 1191.660 ;
        RECT 1855.740 1191.400 1856.000 1191.660 ;
        RECT 1975.800 1191.400 1976.060 1191.660 ;
        RECT 1997.420 1191.400 1997.680 1191.660 ;
        RECT 2042.500 1191.400 2042.760 1191.660 ;
        RECT 2089.420 1191.400 2089.680 1191.660 ;
        RECT 2273.420 1191.400 2273.680 1191.660 ;
        RECT 2276.640 1191.400 2276.900 1191.660 ;
        RECT 2526.420 1191.400 2526.680 1191.660 ;
        RECT 1527.760 1191.060 1528.020 1191.320 ;
        RECT 1714.980 1191.060 1715.240 1191.320 ;
        RECT 1965.680 1191.060 1965.940 1191.320 ;
        RECT 2260.080 1191.060 2260.340 1191.320 ;
        RECT 2260.540 1191.060 2260.800 1191.320 ;
        RECT 2281.240 1191.060 2281.500 1191.320 ;
        RECT 2296.880 1191.060 2297.140 1191.320 ;
        RECT 2482.260 1191.060 2482.520 1191.320 ;
        RECT 1417.360 1190.720 1417.620 1190.980 ;
        RECT 1490.040 1190.720 1490.300 1190.980 ;
        RECT 1516.720 1190.720 1516.980 1190.980 ;
        RECT 1707.620 1190.720 1707.880 1190.980 ;
        RECT 1900.820 1190.720 1901.080 1190.980 ;
        RECT 2053.080 1190.720 2053.340 1190.980 ;
        RECT 2144.160 1190.720 2144.420 1190.980 ;
        RECT 2238.920 1190.720 2239.180 1190.980 ;
        RECT 2242.140 1190.720 2242.400 1190.980 ;
        RECT 2581.620 1190.720 2581.880 1190.980 ;
        RECT 1538.340 1190.380 1538.600 1190.640 ;
        RECT 1735.220 1190.380 1735.480 1190.640 ;
        RECT 1802.840 1190.380 1803.100 1190.640 ;
        RECT 2370.020 1190.380 2370.280 1190.640 ;
        RECT 1427.940 1190.040 1428.200 1190.300 ;
        RECT 1728.320 1190.040 1728.580 1190.300 ;
        RECT 1869.080 1190.040 1869.340 1190.300 ;
        RECT 2481.800 1190.040 2482.060 1190.300 ;
        RECT 2260.080 1189.700 2260.340 1189.960 ;
        RECT 2287.220 1189.700 2287.480 1189.960 ;
        RECT 2324.480 1189.700 2324.740 1189.960 ;
        RECT 2428.900 1189.700 2429.160 1189.960 ;
        RECT 2364.040 1189.360 2364.300 1189.620 ;
        RECT 2438.100 1189.360 2438.360 1189.620 ;
        RECT 1675.880 1189.020 1676.140 1189.280 ;
        RECT 1711.760 1189.020 1712.020 1189.280 ;
        RECT 2338.740 1189.020 2339.000 1189.280 ;
        RECT 2405.440 1189.020 2405.700 1189.280 ;
        RECT 2309.300 1188.680 2309.560 1188.940 ;
        RECT 2364.500 1188.680 2364.760 1188.940 ;
        RECT 1659.780 1188.340 1660.040 1188.600 ;
        RECT 1697.960 1188.340 1698.220 1188.600 ;
        RECT 1880.120 1188.340 1880.380 1188.600 ;
        RECT 1884.260 1188.340 1884.520 1188.600 ;
        RECT 2351.620 1188.340 2351.880 1188.600 ;
        RECT 2383.360 1188.340 2383.620 1188.600 ;
        RECT 1676.340 1188.000 1676.600 1188.260 ;
        RECT 1700.720 1188.000 1700.980 1188.260 ;
        RECT 1669.440 1187.660 1669.700 1187.920 ;
        RECT 1691.060 1187.660 1691.320 1187.920 ;
        RECT 1439.440 1186.980 1439.700 1187.240 ;
        RECT 1441.740 1186.980 1442.000 1187.240 ;
        RECT 1494.640 1186.980 1494.900 1187.240 ;
        RECT 1496.940 1186.980 1497.200 1187.240 ;
        RECT 1604.580 1186.980 1604.840 1187.240 ;
        RECT 1607.340 1186.980 1607.600 1187.240 ;
        RECT 1637.700 1186.980 1637.960 1187.240 ;
        RECT 1641.840 1186.980 1642.100 1187.240 ;
        RECT 1648.740 1186.980 1649.000 1187.240 ;
        RECT 1686.920 1187.320 1687.180 1187.580 ;
        RECT 1834.120 1187.320 1834.380 1187.580 ;
        RECT 1843.780 1187.320 1844.040 1187.580 ;
        RECT 2331.380 1187.320 2331.640 1187.580 ;
        RECT 2363.580 1187.320 2363.840 1187.580 ;
        RECT 1668.520 1186.980 1668.780 1187.240 ;
        RECT 1669.440 1186.980 1669.700 1187.240 ;
        RECT 1684.160 1186.980 1684.420 1187.240 ;
        RECT 1690.600 1186.980 1690.860 1187.240 ;
        RECT 1824.920 1186.980 1825.180 1187.240 ;
        RECT 1831.820 1186.980 1832.080 1187.240 ;
        RECT 1835.040 1186.980 1835.300 1187.240 ;
        RECT 1856.200 1186.980 1856.460 1187.240 ;
        RECT 1913.240 1186.980 1913.500 1187.240 ;
        RECT 1917.840 1186.980 1918.100 1187.240 ;
        RECT 1934.860 1186.980 1935.120 1187.240 ;
        RECT 1938.540 1186.980 1938.800 1187.240 ;
        RECT 1956.940 1186.980 1957.200 1187.240 ;
        RECT 1959.240 1186.980 1959.500 1187.240 ;
        RECT 1976.720 1186.980 1976.980 1187.240 ;
        RECT 1987.300 1186.980 1987.560 1187.240 ;
        RECT 2320.340 1186.980 2320.600 1187.240 ;
        RECT 2324.940 1186.980 2325.200 1187.240 ;
        RECT 2342.420 1186.980 2342.680 1187.240 ;
        RECT 2345.640 1186.980 2345.900 1187.240 ;
        RECT 1648.740 1159.100 1649.000 1159.360 ;
        RECT 1667.600 1159.100 1667.860 1159.360 ;
        RECT 1682.320 1159.100 1682.580 1159.360 ;
        RECT 1684.160 1159.100 1684.420 1159.360 ;
        RECT 1682.780 1104.020 1683.040 1104.280 ;
        RECT 1683.240 1104.020 1683.500 1104.280 ;
        RECT 1683.240 1076.820 1683.500 1077.080 ;
        RECT 1683.240 1076.140 1683.500 1076.400 ;
        RECT 1462.440 1051.660 1462.700 1051.920 ;
        RECT 1496.480 1051.660 1496.740 1051.920 ;
        RECT 2287.220 1028.200 2287.480 1028.460 ;
        RECT 2288.140 1028.200 2288.400 1028.460 ;
        RECT 2352.080 1027.860 2352.340 1028.120 ;
        RECT 2359.900 1027.860 2360.160 1028.120 ;
        RECT 2352.540 1026.160 2352.800 1026.420 ;
        RECT 2373.700 1026.160 2373.960 1026.420 ;
        RECT 2330.920 1025.820 2331.180 1026.080 ;
        RECT 2415.100 1025.820 2415.360 1026.080 ;
        RECT 2345.180 1025.480 2345.440 1025.740 ;
        RECT 2394.400 1025.480 2394.660 1025.740 ;
        RECT 2255.940 1025.140 2256.200 1025.400 ;
        RECT 2415.100 1025.140 2415.360 1025.400 ;
        RECT 2241.680 1024.800 2241.940 1025.060 ;
        RECT 2422.000 1024.800 2422.260 1025.060 ;
        RECT 1890.240 1024.460 1890.500 1024.720 ;
        RECT 2450.980 1024.460 2451.240 1024.720 ;
        RECT 2363.580 1021.740 2363.840 1022.000 ;
        RECT 1686.920 1021.060 1687.180 1021.320 ;
        RECT 1704.400 1021.060 1704.660 1021.320 ;
        RECT 1706.240 1021.060 1706.500 1021.320 ;
        RECT 1732.000 1021.060 1732.260 1021.320 ;
        RECT 1735.220 1021.060 1735.480 1021.320 ;
        RECT 1759.600 1021.060 1759.860 1021.320 ;
        RECT 1831.820 1021.060 1832.080 1021.320 ;
        RECT 1842.400 1021.060 1842.660 1021.320 ;
        RECT 1918.300 1021.060 1918.560 1021.320 ;
        RECT 1966.140 1021.060 1966.400 1021.320 ;
        RECT 2014.900 1021.060 2015.160 1021.320 ;
        RECT 2062.740 1021.060 2063.000 1021.320 ;
        RECT 2111.500 1021.060 2111.760 1021.320 ;
        RECT 2159.340 1021.060 2159.600 1021.320 ;
        RECT 2252.720 1021.060 2252.980 1021.320 ;
        RECT 2254.560 1021.060 2254.820 1021.320 ;
        RECT 2303.320 1021.060 2303.580 1021.320 ;
        RECT 2324.940 1021.060 2325.200 1021.320 ;
        RECT 1496.940 1020.720 1497.200 1020.980 ;
        RECT 1641.840 1020.720 1642.100 1020.980 ;
        RECT 1711.300 1020.720 1711.560 1020.980 ;
        RECT 1717.280 1020.720 1717.540 1020.980 ;
        RECT 1741.660 1020.720 1741.920 1020.980 ;
        RECT 1748.100 1020.720 1748.360 1020.980 ;
        RECT 1752.240 1020.720 1752.500 1020.980 ;
        RECT 1786.740 1020.720 1787.000 1020.980 ;
        RECT 1787.660 1020.720 1787.920 1020.980 ;
        RECT 2215.000 1020.720 2215.260 1020.980 ;
        RECT 2266.520 1020.720 2266.780 1020.980 ;
        RECT 2312.060 1020.720 2312.320 1020.980 ;
        RECT 2318.040 1020.720 2318.300 1020.980 ;
        RECT 2364.040 1020.720 2364.300 1020.980 ;
        RECT 2373.700 1021.060 2373.960 1021.320 ;
        RECT 2383.820 1021.060 2384.080 1021.320 ;
        RECT 2403.140 1021.060 2403.400 1021.320 ;
        RECT 2380.600 1020.720 2380.860 1020.980 ;
        RECT 2384.280 1020.720 2384.540 1020.980 ;
        RECT 2408.200 1020.720 2408.460 1020.980 ;
        RECT 1787.200 1020.380 1787.460 1020.640 ;
        RECT 1790.420 1020.380 1790.680 1020.640 ;
        RECT 2208.100 1020.380 2208.360 1020.640 ;
        RECT 2245.820 1020.380 2246.080 1020.640 ;
        RECT 2293.660 1020.380 2293.920 1020.640 ;
        RECT 2353.920 1020.380 2354.180 1020.640 ;
        RECT 2363.580 1020.380 2363.840 1020.640 ;
        RECT 2364.500 1020.380 2364.760 1020.640 ;
        RECT 2387.500 1020.380 2387.760 1020.640 ;
        RECT 1503.840 1020.040 1504.100 1020.300 ;
        RECT 1780.300 1020.040 1780.560 1020.300 ;
        RECT 1800.080 1020.040 1800.340 1020.300 ;
        RECT 1821.700 1020.040 1821.960 1020.300 ;
        RECT 1869.540 1020.040 1869.800 1020.300 ;
        RECT 1918.300 1020.040 1918.560 1020.300 ;
        RECT 1966.140 1020.040 1966.400 1020.300 ;
        RECT 2014.900 1020.040 2015.160 1020.300 ;
        RECT 2062.740 1020.040 2063.000 1020.300 ;
        RECT 2111.500 1020.040 2111.760 1020.300 ;
        RECT 2159.340 1020.040 2159.600 1020.300 ;
        RECT 2194.300 1020.040 2194.560 1020.300 ;
        RECT 2269.740 1020.040 2270.000 1020.300 ;
        RECT 2532.400 1020.040 2532.660 1020.300 ;
        RECT 1572.840 1019.700 1573.100 1019.960 ;
        RECT 1745.800 1019.700 1746.060 1019.960 ;
        RECT 1759.140 1019.700 1759.400 1019.960 ;
        RECT 1806.060 1019.700 1806.320 1019.960 ;
        RECT 2180.500 1019.700 2180.760 1019.960 ;
        RECT 2276.640 1019.700 2276.900 1019.960 ;
        RECT 2511.700 1019.700 2511.960 1019.960 ;
        RECT 1586.640 1019.360 1586.900 1019.620 ;
        RECT 1738.900 1019.360 1739.160 1019.620 ;
        RECT 1807.900 1019.360 1808.160 1019.620 ;
        RECT 1812.960 1019.360 1813.220 1019.620 ;
        RECT 2173.600 1019.360 2173.860 1019.620 ;
        RECT 2238.920 1019.360 2239.180 1019.620 ;
        RECT 2242.140 1019.360 2242.400 1019.620 ;
        RECT 2287.220 1019.360 2287.480 1019.620 ;
        RECT 2289.980 1019.360 2290.240 1019.620 ;
        RECT 2491.000 1019.360 2491.260 1019.620 ;
        RECT 1593.540 1019.020 1593.800 1019.280 ;
        RECT 1680.020 1019.020 1680.280 1019.280 ;
        RECT 1607.340 1018.680 1607.600 1018.940 ;
        RECT 1714.980 1019.020 1715.240 1019.280 ;
        RECT 1766.500 1019.020 1766.760 1019.280 ;
        RECT 1772.940 1019.020 1773.200 1019.280 ;
        RECT 1817.560 1019.020 1817.820 1019.280 ;
        RECT 2159.800 1019.020 2160.060 1019.280 ;
        RECT 2290.440 1019.020 2290.700 1019.280 ;
        RECT 2394.400 1019.020 2394.660 1019.280 ;
        RECT 1725.100 1018.680 1725.360 1018.940 ;
        RECT 1728.320 1018.680 1728.580 1018.940 ;
        RECT 1821.700 1018.680 1821.960 1018.940 ;
        RECT 1614.240 1018.340 1614.500 1018.600 ;
        RECT 1718.200 1018.340 1718.460 1018.600 ;
        RECT 1628.040 1018.000 1628.300 1018.260 ;
        RECT 1680.020 1017.660 1680.280 1017.920 ;
        RECT 1707.620 1018.000 1707.880 1018.260 ;
        RECT 1773.400 1018.340 1773.660 1018.600 ;
        RECT 1732.000 1018.000 1732.260 1018.260 ;
        RECT 1735.680 1018.000 1735.940 1018.260 ;
        RECT 1641.840 1017.320 1642.100 1017.580 ;
        RECT 1689.680 1017.320 1689.940 1017.580 ;
        RECT 1706.240 1017.320 1706.500 1017.580 ;
        RECT 1711.300 1017.660 1711.560 1017.920 ;
        RECT 1712.220 1017.320 1712.480 1017.580 ;
        RECT 1654.720 1016.980 1654.980 1017.240 ;
        RECT 1700.720 1016.980 1700.980 1017.240 ;
        RECT 1713.600 1017.320 1713.860 1017.580 ;
        RECT 1732.000 1017.320 1732.260 1017.580 ;
        RECT 1675.420 1016.640 1675.680 1016.900 ;
        RECT 1718.200 1016.980 1718.460 1017.240 ;
        RECT 1766.040 1018.000 1766.300 1018.260 ;
        RECT 1807.900 1018.340 1808.160 1018.600 ;
        RECT 1778.000 1018.000 1778.260 1018.260 ;
        RECT 1824.000 1018.680 1824.260 1018.940 ;
        RECT 2152.900 1018.680 2153.160 1018.940 ;
        RECT 2297.340 1018.680 2297.600 1018.940 ;
        RECT 2388.420 1018.680 2388.680 1018.940 ;
        RECT 2304.240 1018.340 2304.500 1018.600 ;
        RECT 2363.120 1018.340 2363.380 1018.600 ;
        RECT 2370.020 1018.340 2370.280 1018.600 ;
        RECT 2428.900 1018.340 2429.160 1018.600 ;
        RECT 2259.620 1018.000 2259.880 1018.260 ;
        RECT 2307.920 1018.000 2308.180 1018.260 ;
        RECT 2355.760 1018.000 2356.020 1018.260 ;
        RECT 1748.100 1017.660 1748.360 1017.920 ;
        RECT 1787.660 1017.660 1787.920 1017.920 ;
        RECT 1822.160 1017.660 1822.420 1017.920 ;
        RECT 1869.540 1017.660 1869.800 1017.920 ;
        RECT 2273.420 1017.660 2273.680 1017.920 ;
        RECT 2317.120 1017.660 2317.380 1017.920 ;
        RECT 2353.920 1017.660 2354.180 1017.920 ;
        RECT 1782.140 1017.320 1782.400 1017.580 ;
        RECT 2228.800 1017.320 2229.060 1017.580 ;
        RECT 2283.540 1017.320 2283.800 1017.580 ;
        RECT 2323.560 1017.320 2323.820 1017.580 ;
        RECT 2373.240 1017.660 2373.500 1017.920 ;
        RECT 2373.700 1017.660 2373.960 1017.920 ;
        RECT 2408.200 1017.660 2408.460 1017.920 ;
        RECT 2358.060 1017.320 2358.320 1017.580 ;
        RECT 2377.840 1017.320 2378.100 1017.580 ;
        RECT 2422.000 1017.320 2422.260 1017.580 ;
        RECT 1748.100 1016.980 1748.360 1017.240 ;
        RECT 1790.420 1016.980 1790.680 1017.240 ;
        RECT 2303.320 1016.980 2303.580 1017.240 ;
        RECT 2347.020 1016.980 2347.280 1017.240 ;
        RECT 2387.960 1016.980 2388.220 1017.240 ;
        RECT 1662.080 1016.300 1662.340 1016.560 ;
        RECT 1707.160 1016.300 1707.420 1016.560 ;
        RECT 1714.520 1016.300 1714.780 1016.560 ;
        RECT 1745.800 1016.300 1746.060 1016.560 ;
        RECT 1766.040 1016.640 1766.300 1016.900 ;
        RECT 2293.660 1016.640 2293.920 1016.900 ;
        RECT 2342.420 1016.640 2342.680 1016.900 ;
        RECT 2387.500 1016.640 2387.760 1016.900 ;
        RECT 2281.240 1016.300 2281.500 1016.560 ;
        RECT 2329.540 1016.300 2329.800 1016.560 ;
        RECT 2358.060 1016.300 2358.320 1016.560 ;
        RECT 2363.580 1016.300 2363.840 1016.560 ;
        RECT 2373.700 1016.300 2373.960 1016.560 ;
        RECT 1668.980 1015.960 1669.240 1016.220 ;
        RECT 1713.600 1015.960 1713.860 1016.220 ;
        RECT 1717.740 1015.960 1718.000 1016.220 ;
        RECT 1721.420 1015.960 1721.680 1016.220 ;
        RECT 1755.460 1015.960 1755.720 1016.220 ;
        RECT 1755.920 1015.960 1756.180 1016.220 ;
        RECT 1800.080 1015.960 1800.340 1016.220 ;
        RECT 2287.220 1015.960 2287.480 1016.220 ;
        RECT 2335.520 1015.960 2335.780 1016.220 ;
        RECT 2380.600 1015.960 2380.860 1016.220 ;
        RECT 2381.060 1015.960 2381.320 1016.220 ;
        RECT 1683.240 1015.620 1683.500 1015.880 ;
        RECT 1729.700 1015.620 1729.960 1015.880 ;
        RECT 1778.000 1015.620 1778.260 1015.880 ;
        RECT 2312.060 1015.620 2312.320 1015.880 ;
        RECT 2355.300 1015.620 2355.560 1015.880 ;
        RECT 2355.760 1015.620 2356.020 1015.880 ;
        RECT 2394.400 1015.620 2394.660 1015.880 ;
        RECT 2402.220 1015.620 2402.480 1015.880 ;
        RECT 1648.740 1015.280 1649.000 1015.540 ;
        RECT 1696.120 1015.280 1696.380 1015.540 ;
        RECT 1717.280 1015.280 1717.540 1015.540 ;
        RECT 1717.740 1015.280 1718.000 1015.540 ;
        RECT 1759.140 1015.280 1759.400 1015.540 ;
        RECT 2255.020 1015.280 2255.280 1015.540 ;
        RECT 2560.000 1015.280 2560.260 1015.540 ;
        RECT 1683.240 1014.940 1683.500 1015.200 ;
        RECT 1724.640 1014.940 1724.900 1015.200 ;
        RECT 1772.940 1014.940 1773.200 1015.200 ;
        RECT 2249.040 1014.940 2249.300 1015.200 ;
        RECT 2566.900 1014.940 2567.160 1015.200 ;
        RECT 1483.140 1014.600 1483.400 1014.860 ;
        RECT 1787.200 1014.600 1787.460 1014.860 ;
        RECT 2345.640 1014.600 2345.900 1014.860 ;
        RECT 2366.800 1014.600 2367.060 1014.860 ;
        RECT 2373.240 1014.600 2373.500 1014.860 ;
        RECT 2415.100 1014.600 2415.360 1014.860 ;
        RECT 1476.240 1014.260 1476.500 1014.520 ;
        RECT 1794.100 1014.260 1794.360 1014.520 ;
        RECT 2262.840 1014.260 2263.100 1014.520 ;
        RECT 2546.200 1014.260 2546.460 1014.520 ;
        RECT 1945.440 1007.120 1945.700 1007.380 ;
        RECT 2498.820 1007.120 2499.080 1007.380 ;
        RECT 1938.540 1006.780 1938.800 1007.040 ;
        RECT 2499.280 1006.780 2499.540 1007.040 ;
        RECT 1924.740 1006.440 1925.000 1006.700 ;
        RECT 2499.740 1006.440 2500.000 1006.700 ;
        RECT 1917.840 1006.100 1918.100 1006.360 ;
        RECT 2500.200 1006.100 2500.460 1006.360 ;
        RECT 1904.040 1005.760 1904.300 1006.020 ;
        RECT 2500.660 1005.760 2500.920 1006.020 ;
        RECT 1959.240 1003.380 1959.500 1003.640 ;
        RECT 2498.360 1003.380 2498.620 1003.640 ;
        RECT 2287.680 1003.040 2287.940 1003.300 ;
        RECT 2497.900 1003.040 2498.160 1003.300 ;
        RECT 2094.020 1001.340 2094.280 1001.600 ;
        RECT 2587.600 1001.340 2587.860 1001.600 ;
        RECT 1898.980 917.360 1899.240 917.620 ;
        RECT 2094.020 917.360 2094.280 917.620 ;
        RECT 1899.900 620.540 1900.160 620.800 ;
        RECT 1976.720 620.540 1976.980 620.800 ;
        RECT 1900.360 593.000 1900.620 593.260 ;
        RECT 1969.820 593.000 1970.080 593.260 ;
        RECT 1900.360 579.400 1900.620 579.660 ;
        RECT 1997.420 579.400 1997.680 579.660 ;
        RECT 2504.340 917.360 2504.600 917.620 ;
        RECT 2587.600 917.360 2587.860 917.620 ;
        RECT 1503.840 554.580 1504.100 554.840 ;
        RECT 2083.900 554.580 2084.160 554.840 ;
      LAYER met2 ;
        RECT 2442.700 3066.810 2442.960 3067.130 ;
        RECT 2469.840 3066.810 2470.100 3067.130 ;
        RECT 2442.760 3064.070 2442.900 3066.810 ;
        RECT 2469.900 3064.070 2470.040 3066.810 ;
        RECT 1868.160 3063.925 1868.420 3064.070 ;
        RECT 1868.150 3063.555 1868.430 3063.925 ;
        RECT 1898.060 3063.750 1898.320 3064.070 ;
        RECT 2442.700 3063.925 2442.960 3064.070 ;
        RECT 2469.840 3063.925 2470.100 3064.070 ;
        RECT 1490.030 3032.955 1490.310 3033.325 ;
        RECT 1489.570 3026.835 1489.850 3027.205 ;
        RECT 1489.110 3018.675 1489.390 3019.045 ;
        RECT 1488.650 3012.555 1488.930 3012.925 ;
        RECT 1488.190 3004.395 1488.470 3004.765 ;
        RECT 1487.730 2998.955 1488.010 2999.325 ;
        RECT 1487.270 2990.115 1487.550 2990.485 ;
        RECT 1486.810 2701.115 1487.090 2701.485 ;
        RECT 1486.350 2692.275 1486.630 2692.645 ;
        RECT 1486.420 2604.730 1486.560 2692.275 ;
        RECT 1486.360 2604.410 1486.620 2604.730 ;
        RECT 1476.240 2592.850 1476.500 2593.170 ;
        RECT 1462.440 2591.830 1462.700 2592.150 ;
        RECT 1448.640 2591.490 1448.900 2591.810 ;
        RECT 1441.740 2587.750 1442.000 2588.070 ;
        RECT 1427.940 2587.410 1428.200 2587.730 ;
        RECT 1406.780 2411.630 1407.040 2411.950 ;
        RECT 1405.150 2399.450 1405.430 2400.000 ;
        RECT 1406.840 2399.450 1406.980 2411.630 ;
        RECT 1417.350 2410.755 1417.630 2411.125 ;
        RECT 1405.150 2399.310 1406.980 2399.450 ;
        RECT 1415.730 2399.450 1416.010 2400.000 ;
        RECT 1417.420 2399.450 1417.560 2410.755 ;
        RECT 1415.730 2399.310 1417.560 2399.450 ;
        RECT 1426.770 2399.450 1427.050 2400.000 ;
        RECT 1428.000 2399.450 1428.140 2587.410 ;
        RECT 1441.800 2412.970 1441.940 2587.750 ;
        RECT 1439.440 2412.650 1439.700 2412.970 ;
        RECT 1441.740 2412.650 1442.000 2412.970 ;
        RECT 1426.770 2399.310 1428.140 2399.450 ;
        RECT 1437.810 2399.450 1438.090 2400.000 ;
        RECT 1439.500 2399.450 1439.640 2412.650 ;
        RECT 1448.700 2400.130 1448.840 2591.490 ;
        RECT 1448.700 2400.000 1449.070 2400.130 ;
        RECT 1448.700 2399.990 1449.130 2400.000 ;
        RECT 1437.810 2399.310 1439.640 2399.450 ;
        RECT 1405.150 2396.000 1405.430 2399.310 ;
        RECT 1415.730 2396.000 1416.010 2399.310 ;
        RECT 1426.770 2396.000 1427.050 2399.310 ;
        RECT 1437.810 2396.000 1438.090 2399.310 ;
        RECT 1448.850 2396.000 1449.130 2399.990 ;
        RECT 1459.890 2398.770 1460.170 2400.000 ;
        RECT 1462.500 2398.770 1462.640 2591.830 ;
        RECT 1476.300 2409.570 1476.440 2592.850 ;
        RECT 1483.140 2589.450 1483.400 2589.770 ;
        RECT 1472.560 2409.250 1472.820 2409.570 ;
        RECT 1476.240 2409.250 1476.500 2409.570 ;
        RECT 1459.890 2398.630 1462.640 2398.770 ;
        RECT 1470.930 2399.450 1471.210 2400.000 ;
        RECT 1472.620 2399.450 1472.760 2409.250 ;
        RECT 1470.930 2399.310 1472.760 2399.450 ;
        RECT 1481.970 2399.450 1482.250 2400.000 ;
        RECT 1483.200 2399.450 1483.340 2589.450 ;
        RECT 1486.880 2410.930 1487.020 2701.115 ;
        RECT 1487.340 2411.270 1487.480 2990.115 ;
        RECT 1487.800 2415.010 1487.940 2998.955 ;
        RECT 1487.740 2414.690 1488.000 2415.010 ;
        RECT 1488.260 2414.670 1488.400 3004.395 ;
        RECT 1488.200 2414.350 1488.460 2414.670 ;
        RECT 1488.720 2414.330 1488.860 3012.555 ;
        RECT 1488.660 2414.010 1488.920 2414.330 ;
        RECT 1489.180 2413.990 1489.320 3018.675 ;
        RECT 1489.120 2413.670 1489.380 2413.990 ;
        RECT 1489.640 2413.650 1489.780 3026.835 ;
        RECT 1489.580 2413.330 1489.840 2413.650 ;
        RECT 1490.100 2411.805 1490.240 3032.955 ;
      LAYER met2 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
      LAYER met2 ;
        RECT 1898.120 2747.045 1898.260 3063.750 ;
        RECT 2442.690 3063.555 2442.970 3063.925 ;
        RECT 2469.830 3063.555 2470.110 3063.925 ;
        RECT 2497.900 3063.750 2498.160 3064.070 ;
        RECT 1899.900 3051.850 1900.160 3052.170 ;
        RECT 2482.260 3051.850 2482.520 3052.170 ;
        RECT 1899.960 3048.285 1900.100 3051.850 ;
        RECT 1898.510 3047.915 1898.790 3048.285 ;
        RECT 1899.890 3047.915 1900.170 3048.285 ;
        RECT 1898.050 2746.675 1898.330 2747.045 ;
        RECT 1898.050 2704.515 1898.330 2704.885 ;
        RECT 1614.700 2594.210 1614.960 2594.530 ;
        RECT 1661.620 2594.210 1661.880 2594.530 ;
        RECT 1537.880 2593.870 1538.140 2594.190 ;
        RECT 1614.760 2594.045 1614.900 2594.210 ;
        RECT 1621.600 2594.045 1621.860 2594.190 ;
        RECT 1517.640 2590.470 1517.900 2590.790 ;
        RECT 1496.940 2589.790 1497.200 2590.110 ;
        RECT 1497.000 2412.970 1497.140 2589.790 ;
        RECT 1503.380 2588.770 1503.640 2589.090 ;
        RECT 1494.640 2412.650 1494.900 2412.970 ;
        RECT 1496.940 2412.650 1497.200 2412.970 ;
        RECT 1490.030 2411.435 1490.310 2411.805 ;
        RECT 1487.280 2410.950 1487.540 2411.270 ;
        RECT 1486.820 2410.610 1487.080 2410.930 ;
        RECT 1481.970 2399.310 1483.340 2399.450 ;
        RECT 1493.010 2399.450 1493.290 2400.000 ;
        RECT 1494.700 2399.450 1494.840 2412.650 ;
        RECT 1493.010 2399.310 1494.840 2399.450 ;
        RECT 1503.440 2399.450 1503.580 2588.770 ;
        RECT 1510.340 2411.610 1511.860 2411.690 ;
        RECT 1510.340 2411.550 1511.920 2411.610 ;
        RECT 1510.340 2410.930 1510.480 2411.550 ;
        RECT 1511.660 2411.290 1511.920 2411.550 ;
        RECT 1510.740 2411.010 1511.000 2411.270 ;
        RECT 1511.200 2411.010 1511.460 2411.270 ;
        RECT 1510.740 2410.950 1511.460 2411.010 ;
        RECT 1510.280 2410.610 1510.540 2410.930 ;
        RECT 1510.800 2410.870 1511.400 2410.950 ;
        RECT 1517.700 2400.130 1517.840 2590.470 ;
        RECT 1531.440 2590.130 1531.700 2590.450 ;
        RECT 1531.500 2412.970 1531.640 2590.130 ;
        RECT 1527.760 2412.650 1528.020 2412.970 ;
        RECT 1531.440 2412.650 1531.700 2412.970 ;
        RECT 1504.050 2399.450 1504.330 2400.000 ;
        RECT 1503.440 2399.310 1504.330 2399.450 ;
        RECT 1459.890 2396.000 1460.170 2398.630 ;
        RECT 1470.930 2396.000 1471.210 2399.310 ;
        RECT 1481.970 2396.000 1482.250 2399.310 ;
        RECT 1493.010 2396.000 1493.290 2399.310 ;
        RECT 1504.050 2396.000 1504.330 2399.310 ;
        RECT 1515.090 2399.450 1515.370 2400.000 ;
        RECT 1516.780 2399.990 1517.840 2400.130 ;
        RECT 1516.780 2399.450 1516.920 2399.990 ;
        RECT 1515.090 2399.310 1516.920 2399.450 ;
        RECT 1526.130 2399.450 1526.410 2400.000 ;
        RECT 1527.820 2399.450 1527.960 2412.650 ;
        RECT 1526.130 2399.310 1527.960 2399.450 ;
        RECT 1537.170 2399.450 1537.450 2400.000 ;
        RECT 1537.940 2399.450 1538.080 2593.870 ;
        RECT 1569.610 2593.675 1569.890 2594.045 ;
        RECT 1573.750 2593.675 1574.030 2594.045 ;
        RECT 1586.630 2593.675 1586.910 2594.045 ;
        RECT 1591.230 2593.675 1591.510 2594.045 ;
        RECT 1598.590 2593.675 1598.870 2594.045 ;
        RECT 1604.110 2593.675 1604.390 2594.045 ;
        RECT 1614.690 2593.675 1614.970 2594.045 ;
        RECT 1621.590 2593.675 1621.870 2594.045 ;
        RECT 1626.650 2593.675 1626.930 2594.045 ;
        RECT 1651.030 2593.675 1651.310 2594.045 ;
        RECT 1656.100 2593.870 1656.360 2594.190 ;
        RECT 1661.680 2594.045 1661.820 2594.210 ;
        RECT 1569.680 2592.830 1569.820 2593.675 ;
        RECT 1565.470 2592.315 1565.750 2592.685 ;
        RECT 1569.620 2592.510 1569.880 2592.830 ;
        RECT 1573.290 2592.315 1573.570 2592.685 ;
        RECT 1573.820 2592.490 1573.960 2593.675 ;
        RECT 1586.640 2593.530 1586.900 2593.675 ;
        RECT 1581.110 2592.995 1581.390 2593.365 ;
        RECT 1587.090 2592.995 1587.370 2593.365 ;
        RECT 1565.540 2591.470 1565.680 2592.315 ;
        RECT 1573.360 2591.810 1573.500 2592.315 ;
        RECT 1573.760 2592.170 1574.020 2592.490 ;
        RECT 1581.180 2592.150 1581.320 2592.995 ;
        RECT 1587.100 2592.850 1587.360 2592.995 ;
        RECT 1591.300 2592.830 1591.440 2593.675 ;
        RECT 1598.660 2593.510 1598.800 2593.675 ;
        RECT 1598.600 2593.190 1598.860 2593.510 ;
        RECT 1604.180 2593.170 1604.320 2593.675 ;
        RECT 1604.120 2592.850 1604.380 2593.170 ;
        RECT 1591.240 2592.510 1591.500 2592.830 ;
        RECT 1608.250 2592.315 1608.530 2592.685 ;
        RECT 1614.760 2592.490 1614.900 2593.675 ;
        RECT 1626.660 2593.530 1626.920 2593.675 ;
        RECT 1644.660 2593.510 1644.800 2593.665 ;
        RECT 1651.100 2593.510 1651.240 2593.675 ;
        RECT 1644.600 2593.365 1644.860 2593.510 ;
        RECT 1639.070 2592.995 1639.350 2593.365 ;
        RECT 1644.590 2592.995 1644.870 2593.365 ;
        RECT 1651.040 2593.190 1651.300 2593.510 ;
        RECT 1656.160 2593.365 1656.300 2593.870 ;
        RECT 1661.610 2593.675 1661.890 2594.045 ;
        RECT 1669.890 2593.675 1670.170 2594.045 ;
        RECT 1690.590 2593.675 1690.870 2594.045 ;
        RECT 1697.950 2593.675 1698.230 2594.045 ;
        RECT 1702.560 2593.870 1702.820 2594.190 ;
        RECT 1656.090 2592.995 1656.370 2593.365 ;
        RECT 1661.680 2593.170 1661.820 2593.675 ;
        RECT 1669.900 2593.530 1670.160 2593.675 ;
        RECT 1690.600 2593.530 1690.860 2593.675 ;
        RECT 1639.140 2592.830 1639.280 2592.995 ;
        RECT 1581.120 2591.830 1581.380 2592.150 ;
        RECT 1573.300 2591.490 1573.560 2591.810 ;
        RECT 1607.790 2591.635 1608.070 2592.005 ;
        RECT 1565.480 2591.150 1565.740 2591.470 ;
        RECT 1586.170 2590.955 1586.450 2591.325 ;
        RECT 1566.390 2589.595 1566.670 2589.965 ;
        RECT 1551.680 2588.090 1551.940 2588.410 ;
        RECT 1552.130 2588.235 1552.410 2588.605 ;
        RECT 1558.580 2588.430 1558.840 2588.750 ;
        RECT 1538.330 2587.555 1538.610 2587.925 ;
        RECT 1545.230 2587.555 1545.510 2587.925 ;
        RECT 1551.210 2587.555 1551.490 2587.925 ;
        RECT 1538.400 2410.930 1538.540 2587.555 ;
        RECT 1545.300 2413.310 1545.440 2587.555 ;
        RECT 1545.240 2412.990 1545.500 2413.310 ;
        RECT 1551.280 2412.970 1551.420 2587.555 ;
        RECT 1551.220 2412.650 1551.480 2412.970 ;
        RECT 1538.340 2410.610 1538.600 2410.930 ;
        RECT 1551.740 2405.570 1551.880 2588.090 ;
        RECT 1552.200 2412.630 1552.340 2588.235 ;
        RECT 1552.140 2412.310 1552.400 2412.630 ;
        RECT 1550.360 2405.430 1551.880 2405.570 ;
        RECT 1537.170 2399.310 1538.080 2399.450 ;
        RECT 1548.210 2399.450 1548.490 2400.000 ;
        RECT 1550.360 2399.450 1550.500 2405.430 ;
        RECT 1548.210 2399.310 1550.500 2399.450 ;
        RECT 1558.640 2399.450 1558.780 2588.430 ;
        RECT 1559.490 2588.235 1559.770 2588.605 ;
        RECT 1559.030 2587.555 1559.310 2587.925 ;
        RECT 1559.560 2587.730 1559.700 2588.235 ;
        RECT 1566.460 2588.070 1566.600 2589.595 ;
        RECT 1586.240 2588.070 1586.380 2590.955 ;
        RECT 1607.860 2590.790 1608.000 2591.635 ;
        RECT 1608.320 2591.470 1608.460 2592.315 ;
        RECT 1614.700 2592.170 1614.960 2592.490 ;
        RECT 1621.590 2592.315 1621.870 2592.685 ;
        RECT 1621.660 2591.810 1621.800 2592.315 ;
        RECT 1630.800 2592.170 1631.060 2592.490 ;
        RECT 1633.550 2592.315 1633.830 2592.685 ;
        RECT 1639.080 2592.510 1639.340 2592.830 ;
        RECT 1633.560 2592.170 1633.820 2592.315 ;
        RECT 1621.600 2591.490 1621.860 2591.810 ;
        RECT 1608.260 2591.150 1608.520 2591.470 ;
        RECT 1614.690 2590.955 1614.970 2591.325 ;
        RECT 1593.990 2590.275 1594.270 2590.645 ;
        RECT 1607.800 2590.470 1608.060 2590.790 ;
        RECT 1614.760 2590.450 1614.900 2590.955 ;
        RECT 1594.060 2590.110 1594.200 2590.275 ;
        RECT 1614.700 2590.130 1614.960 2590.450 ;
        RECT 1587.090 2589.595 1587.370 2589.965 ;
        RECT 1594.000 2589.790 1594.260 2590.110 ;
        RECT 1600.890 2589.595 1601.170 2589.965 ;
        RECT 1587.100 2589.450 1587.360 2589.595 ;
        RECT 1586.640 2589.110 1586.900 2589.430 ;
        RECT 1566.400 2587.750 1566.660 2588.070 ;
        RECT 1586.180 2587.750 1586.440 2588.070 ;
        RECT 1559.100 2412.290 1559.240 2587.555 ;
        RECT 1559.500 2587.410 1559.760 2587.730 ;
        RECT 1572.840 2587.410 1573.100 2587.730 ;
        RECT 1559.040 2411.970 1559.300 2412.290 ;
        RECT 1559.500 2411.290 1559.760 2411.610 ;
        RECT 1559.560 2410.250 1559.700 2411.290 ;
        RECT 1559.500 2409.930 1559.760 2410.250 ;
        RECT 1559.250 2399.450 1559.530 2400.000 ;
        RECT 1558.640 2399.310 1559.530 2399.450 ;
        RECT 1515.090 2396.000 1515.370 2399.310 ;
        RECT 1526.130 2396.000 1526.410 2399.310 ;
        RECT 1537.170 2396.000 1537.450 2399.310 ;
        RECT 1548.210 2396.000 1548.490 2399.310 ;
        RECT 1559.250 2396.000 1559.530 2399.310 ;
        RECT 1570.290 2398.770 1570.570 2400.000 ;
        RECT 1572.900 2398.770 1573.040 2587.410 ;
        RECT 1586.700 2409.570 1586.840 2589.110 ;
        RECT 1600.960 2589.090 1601.100 2589.595 ;
        RECT 1614.240 2589.450 1614.500 2589.770 ;
        RECT 1600.900 2588.770 1601.160 2589.090 ;
        RECT 1607.340 2588.770 1607.600 2589.090 ;
        RECT 1593.990 2410.075 1594.270 2410.445 ;
        RECT 1594.000 2409.930 1594.260 2410.075 ;
        RECT 1593.540 2409.590 1593.800 2409.910 ;
        RECT 1582.500 2409.250 1582.760 2409.570 ;
        RECT 1586.640 2409.250 1586.900 2409.570 ;
        RECT 1570.290 2398.630 1573.040 2398.770 ;
        RECT 1580.870 2399.450 1581.150 2400.000 ;
        RECT 1582.560 2399.450 1582.700 2409.250 ;
        RECT 1580.870 2399.310 1582.700 2399.450 ;
        RECT 1591.910 2399.450 1592.190 2400.000 ;
        RECT 1593.600 2399.450 1593.740 2409.590 ;
        RECT 1607.400 2409.570 1607.540 2588.770 ;
        RECT 1609.640 2411.290 1609.900 2411.610 ;
        RECT 1609.700 2410.445 1609.840 2411.290 ;
        RECT 1609.630 2410.075 1609.910 2410.445 ;
        RECT 1604.580 2409.250 1604.840 2409.570 ;
        RECT 1607.340 2409.250 1607.600 2409.570 ;
        RECT 1591.910 2399.310 1593.740 2399.450 ;
        RECT 1602.950 2399.450 1603.230 2400.000 ;
        RECT 1604.640 2399.450 1604.780 2409.250 ;
        RECT 1614.300 2400.810 1614.440 2589.450 ;
        RECT 1621.590 2588.235 1621.870 2588.605 ;
        RECT 1621.600 2588.090 1621.860 2588.235 ;
        RECT 1630.860 2588.070 1631.000 2592.170 ;
        RECT 1644.660 2592.150 1644.800 2592.995 ;
        RECT 1644.600 2591.830 1644.860 2592.150 ;
        RECT 1656.160 2591.470 1656.300 2592.995 ;
        RECT 1661.620 2592.850 1661.880 2593.170 ;
        RECT 1667.130 2592.315 1667.410 2592.685 ;
        RECT 1667.200 2591.810 1667.340 2592.315 ;
        RECT 1667.140 2591.490 1667.400 2591.810 ;
        RECT 1669.960 2591.470 1670.100 2593.530 ;
        RECT 1679.550 2592.995 1679.830 2593.365 ;
        RECT 1679.620 2592.490 1679.760 2592.995 ;
        RECT 1685.080 2592.570 1685.340 2592.830 ;
        RECT 1685.530 2592.570 1685.810 2592.685 ;
        RECT 1686.460 2592.570 1686.720 2592.830 ;
        RECT 1685.080 2592.510 1686.720 2592.570 ;
        RECT 1679.560 2592.170 1679.820 2592.490 ;
        RECT 1685.140 2592.430 1686.660 2592.510 ;
        RECT 1685.530 2592.315 1685.810 2592.430 ;
        RECT 1685.600 2592.015 1685.740 2592.315 ;
        RECT 1690.660 2592.150 1690.800 2593.530 ;
        RECT 1698.020 2593.510 1698.160 2593.675 ;
        RECT 1697.960 2593.190 1698.220 2593.510 ;
        RECT 1702.620 2592.685 1702.760 2593.870 ;
        RECT 1738.430 2593.675 1738.710 2594.045 ;
        RECT 1738.440 2593.530 1738.700 2593.675 ;
        RECT 1707.610 2592.995 1707.890 2593.365 ;
        RECT 1732.910 2592.995 1733.190 2593.365 ;
        RECT 1707.620 2592.850 1707.880 2592.995 ;
        RECT 1732.920 2592.850 1733.180 2592.995 ;
        RECT 1702.550 2592.315 1702.830 2592.685 ;
        RECT 1690.600 2591.830 1690.860 2592.150 ;
        RECT 1656.100 2591.150 1656.360 2591.470 ;
        RECT 1669.900 2591.150 1670.160 2591.470 ;
        RECT 1656.090 2590.275 1656.370 2590.645 ;
        RECT 1678.630 2590.275 1678.910 2590.645 ;
        RECT 1642.290 2589.595 1642.570 2589.965 ;
        RECT 1642.360 2589.430 1642.500 2589.595 ;
        RECT 1631.250 2588.915 1631.530 2589.285 ;
        RECT 1642.300 2589.110 1642.560 2589.430 ;
        RECT 1652.420 2589.110 1652.680 2589.430 ;
        RECT 1631.320 2588.750 1631.460 2588.915 ;
        RECT 1631.260 2588.430 1631.520 2588.750 ;
        RECT 1635.390 2588.235 1635.670 2588.605 ;
        RECT 1635.460 2588.070 1635.600 2588.235 ;
        RECT 1641.840 2588.090 1642.100 2588.410 ;
        RECT 1630.800 2587.750 1631.060 2588.070 ;
        RECT 1635.400 2587.750 1635.660 2588.070 ;
        RECT 1638.620 2587.750 1638.880 2588.070 ;
        RECT 1631.720 2587.410 1631.980 2587.730 ;
        RECT 1626.660 2410.270 1626.920 2410.590 ;
        RECT 1614.070 2400.670 1614.440 2400.810 ;
        RECT 1614.070 2400.000 1614.210 2400.670 ;
        RECT 1602.950 2399.310 1604.780 2399.450 ;
        RECT 1570.290 2396.000 1570.570 2398.630 ;
        RECT 1580.870 2396.000 1581.150 2399.310 ;
        RECT 1591.910 2396.000 1592.190 2399.310 ;
        RECT 1602.950 2396.000 1603.230 2399.310 ;
        RECT 1613.990 2396.000 1614.270 2400.000 ;
        RECT 1625.030 2399.450 1625.310 2400.000 ;
        RECT 1626.720 2399.450 1626.860 2410.270 ;
        RECT 1631.780 2409.910 1631.920 2587.410 ;
        RECT 1638.680 2410.590 1638.820 2587.750 ;
        RECT 1638.620 2410.270 1638.880 2410.590 ;
        RECT 1631.720 2409.590 1631.980 2409.910 ;
        RECT 1641.900 2409.570 1642.040 2588.090 ;
        RECT 1649.190 2587.555 1649.470 2587.925 ;
        RECT 1649.200 2587.410 1649.460 2587.555 ;
        RECT 1652.480 2410.590 1652.620 2589.110 ;
        RECT 1656.160 2589.090 1656.300 2590.275 ;
        RECT 1662.990 2589.595 1663.270 2589.965 ;
        RECT 1663.000 2589.450 1663.260 2589.595 ;
        RECT 1678.700 2589.430 1678.840 2590.275 ;
        RECT 1702.620 2590.110 1702.760 2592.315 ;
        RECT 1702.560 2589.790 1702.820 2590.110 ;
        RECT 1707.680 2589.770 1707.820 2592.850 ;
        RECT 1738.500 2592.830 1738.640 2593.530 ;
        RECT 1744.020 2593.510 1744.160 2593.665 ;
        RECT 1743.960 2593.365 1744.220 2593.510 ;
        RECT 1743.950 2592.995 1744.230 2593.365 ;
        RECT 1725.550 2592.315 1725.830 2592.685 ;
        RECT 1738.440 2592.510 1738.700 2592.830 ;
        RECT 1744.020 2592.490 1744.160 2592.995 ;
        RECT 1725.560 2592.170 1725.820 2592.315 ;
        RECT 1731.540 2592.170 1731.800 2592.490 ;
        RECT 1743.960 2592.170 1744.220 2592.490 ;
        RECT 1713.130 2591.635 1713.410 2592.005 ;
        RECT 1718.190 2591.635 1718.470 2592.005 ;
        RECT 1713.140 2591.490 1713.400 2591.635 ;
        RECT 1707.620 2589.450 1707.880 2589.770 ;
        RECT 1678.640 2589.110 1678.900 2589.430 ;
        RECT 1656.100 2588.770 1656.360 2589.090 ;
        RECT 1683.690 2588.915 1683.970 2589.285 ;
        RECT 1690.590 2588.915 1690.870 2589.285 ;
        RECT 1662.990 2588.235 1663.270 2588.605 ;
        RECT 1669.440 2588.430 1669.700 2588.750 ;
        RECT 1663.060 2588.070 1663.200 2588.235 ;
        RECT 1663.000 2587.750 1663.260 2588.070 ;
        RECT 1666.220 2587.410 1666.480 2587.730 ;
        RECT 1656.100 2411.290 1656.360 2411.610 ;
        RECT 1648.740 2410.270 1649.000 2410.590 ;
        RECT 1652.420 2410.270 1652.680 2410.590 ;
        RECT 1637.700 2409.250 1637.960 2409.570 ;
        RECT 1641.840 2409.250 1642.100 2409.570 ;
        RECT 1625.030 2399.310 1626.860 2399.450 ;
        RECT 1636.070 2399.450 1636.350 2400.000 ;
        RECT 1637.760 2399.450 1637.900 2409.250 ;
        RECT 1636.070 2399.310 1637.900 2399.450 ;
        RECT 1647.110 2399.450 1647.390 2400.000 ;
        RECT 1648.800 2399.450 1648.940 2410.270 ;
        RECT 1656.160 2410.250 1656.300 2411.290 ;
        RECT 1666.280 2410.590 1666.420 2587.410 ;
        RECT 1659.780 2410.270 1660.040 2410.590 ;
        RECT 1666.220 2410.270 1666.480 2410.590 ;
        RECT 1656.100 2409.930 1656.360 2410.250 ;
        RECT 1647.110 2399.310 1648.940 2399.450 ;
        RECT 1658.150 2399.450 1658.430 2400.000 ;
        RECT 1659.840 2399.450 1659.980 2410.270 ;
        RECT 1669.500 2400.810 1669.640 2588.430 ;
        RECT 1669.890 2588.235 1670.170 2588.605 ;
        RECT 1669.900 2588.090 1670.160 2588.235 ;
        RECT 1683.760 2587.730 1683.900 2588.915 ;
        RECT 1690.660 2588.750 1690.800 2588.915 ;
        RECT 1690.600 2588.430 1690.860 2588.750 ;
        RECT 1697.490 2588.235 1697.770 2588.605 ;
        RECT 1683.700 2587.410 1683.960 2587.730 ;
        RECT 1686.920 2587.410 1687.180 2587.730 ;
        RECT 1697.030 2587.555 1697.310 2587.925 ;
        RECT 1697.560 2587.730 1697.700 2588.235 ;
        RECT 1713.200 2588.070 1713.340 2591.490 ;
        RECT 1718.260 2591.470 1718.400 2591.635 ;
        RECT 1718.200 2591.150 1718.460 2591.470 ;
        RECT 1718.260 2589.430 1718.400 2591.150 ;
        RECT 1718.200 2589.110 1718.460 2589.430 ;
        RECT 1731.600 2588.410 1731.740 2592.170 ;
        RECT 1779.840 2590.130 1780.100 2590.450 ;
        RECT 1731.540 2588.090 1731.800 2588.410 ;
        RECT 1745.330 2588.235 1745.610 2588.605 ;
        RECT 1686.980 2410.250 1687.120 2587.410 ;
        RECT 1681.860 2409.930 1682.120 2410.250 ;
        RECT 1686.920 2409.930 1687.180 2410.250 ;
        RECT 1669.270 2400.670 1669.640 2400.810 ;
        RECT 1669.270 2400.000 1669.410 2400.670 ;
        RECT 1658.150 2399.310 1659.980 2399.450 ;
        RECT 1625.030 2396.000 1625.310 2399.310 ;
        RECT 1636.070 2396.000 1636.350 2399.310 ;
        RECT 1647.110 2396.000 1647.390 2399.310 ;
        RECT 1658.150 2396.000 1658.430 2399.310 ;
        RECT 1669.190 2396.000 1669.470 2400.000 ;
        RECT 1680.230 2399.450 1680.510 2400.000 ;
        RECT 1681.920 2399.450 1682.060 2409.930 ;
        RECT 1697.100 2408.890 1697.240 2587.555 ;
        RECT 1697.500 2587.410 1697.760 2587.730 ;
        RECT 1703.930 2587.555 1704.210 2587.925 ;
        RECT 1713.140 2587.750 1713.400 2588.070 ;
        RECT 1714.510 2587.555 1714.790 2587.925 ;
        RECT 1721.410 2587.555 1721.690 2587.925 ;
        RECT 1731.530 2587.555 1731.810 2587.925 ;
        RECT 1736.590 2587.555 1736.870 2587.925 ;
        RECT 1703.020 2411.290 1703.280 2411.610 ;
        RECT 1703.080 2410.590 1703.220 2411.290 ;
        RECT 1703.480 2410.950 1703.740 2411.270 ;
        RECT 1703.020 2410.270 1703.280 2410.590 ;
        RECT 1703.540 2410.250 1703.680 2410.950 ;
        RECT 1703.480 2409.930 1703.740 2410.250 ;
        RECT 1692.900 2408.570 1693.160 2408.890 ;
        RECT 1697.040 2408.570 1697.300 2408.890 ;
        RECT 1680.230 2399.310 1682.060 2399.450 ;
        RECT 1691.270 2399.450 1691.550 2400.000 ;
        RECT 1692.960 2399.450 1693.100 2408.570 ;
        RECT 1691.270 2399.310 1693.100 2399.450 ;
        RECT 1702.310 2399.450 1702.590 2400.000 ;
        RECT 1704.000 2399.450 1704.140 2587.555 ;
        RECT 1714.060 2410.950 1714.320 2411.270 ;
        RECT 1714.120 2410.250 1714.260 2410.950 ;
        RECT 1714.060 2409.930 1714.320 2410.250 ;
        RECT 1702.310 2399.310 1704.140 2399.450 ;
        RECT 1713.350 2399.450 1713.630 2400.000 ;
        RECT 1714.580 2399.450 1714.720 2587.555 ;
        RECT 1713.350 2399.310 1714.720 2399.450 ;
        RECT 1680.230 2396.000 1680.510 2399.310 ;
        RECT 1691.270 2396.000 1691.550 2399.310 ;
        RECT 1702.310 2396.000 1702.590 2399.310 ;
        RECT 1713.350 2396.000 1713.630 2399.310 ;
        RECT 1721.480 2398.770 1721.620 2587.555 ;
        RECT 1731.600 2410.590 1731.740 2587.555 ;
        RECT 1736.600 2587.410 1736.860 2587.555 ;
        RECT 1742.120 2587.410 1742.380 2587.730 ;
        RECT 1744.870 2587.555 1745.150 2587.925 ;
        RECT 1742.180 2410.590 1742.320 2587.410 ;
        RECT 1731.540 2410.270 1731.800 2410.590 ;
        RECT 1733.840 2410.270 1734.100 2410.590 ;
        RECT 1742.120 2410.270 1742.380 2410.590 ;
        RECT 1724.390 2398.770 1724.670 2400.000 ;
        RECT 1733.900 2399.450 1734.040 2410.270 ;
        RECT 1744.940 2409.910 1745.080 2587.555 ;
        RECT 1745.400 2411.010 1745.540 2588.235 ;
        RECT 1752.700 2411.290 1752.960 2411.610 ;
        RECT 1745.400 2410.870 1746.460 2411.010 ;
        RECT 1746.320 2410.590 1746.460 2410.870 ;
        RECT 1745.800 2410.270 1746.060 2410.590 ;
        RECT 1746.260 2410.270 1746.520 2410.590 ;
        RECT 1744.880 2409.590 1745.140 2409.910 ;
        RECT 1735.430 2399.450 1735.710 2400.000 ;
        RECT 1733.900 2399.310 1735.710 2399.450 ;
        RECT 1745.860 2399.450 1746.000 2410.270 ;
        RECT 1752.760 2410.250 1752.900 2411.290 ;
        RECT 1755.460 2410.270 1755.720 2410.590 ;
        RECT 1752.700 2409.930 1752.960 2410.250 ;
        RECT 1746.470 2399.450 1746.750 2400.000 ;
        RECT 1745.860 2399.310 1746.750 2399.450 ;
        RECT 1755.520 2399.450 1755.660 2410.270 ;
        RECT 1766.500 2409.590 1766.760 2409.910 ;
        RECT 1757.050 2399.450 1757.330 2400.000 ;
        RECT 1755.520 2399.310 1757.330 2399.450 ;
        RECT 1766.560 2399.450 1766.700 2409.590 ;
        RECT 1768.090 2399.450 1768.370 2400.000 ;
        RECT 1766.560 2399.310 1768.370 2399.450 ;
        RECT 1721.480 2398.630 1724.670 2398.770 ;
        RECT 1724.390 2396.000 1724.670 2398.630 ;
        RECT 1735.430 2396.000 1735.710 2399.310 ;
        RECT 1746.470 2396.000 1746.750 2399.310 ;
        RECT 1757.050 2396.000 1757.330 2399.310 ;
        RECT 1768.090 2396.000 1768.370 2399.310 ;
        RECT 1779.130 2399.450 1779.410 2400.000 ;
        RECT 1779.900 2399.450 1780.040 2590.130 ;
        RECT 1887.940 2414.690 1888.200 2415.010 ;
        RECT 1835.950 2412.115 1836.230 2412.485 ;
        RECT 1877.350 2412.115 1877.630 2412.485 ;
        RECT 1800.540 2411.290 1800.800 2411.610 ;
        RECT 1835.500 2411.520 1835.760 2411.610 ;
        RECT 1836.020 2411.520 1836.160 2412.115 ;
        RECT 1835.500 2411.380 1836.160 2411.520 ;
        RECT 1835.500 2411.290 1835.760 2411.380 ;
        RECT 1791.800 2410.270 1792.060 2410.590 ;
        RECT 1779.130 2399.310 1780.040 2399.450 ;
        RECT 1790.170 2399.450 1790.450 2400.000 ;
        RECT 1791.860 2399.450 1792.000 2410.270 ;
        RECT 1800.600 2410.250 1800.740 2411.290 ;
        RECT 1877.420 2411.270 1877.560 2412.115 ;
        RECT 1876.900 2410.950 1877.160 2411.270 ;
        RECT 1877.360 2410.950 1877.620 2411.270 ;
        RECT 1865.860 2410.610 1866.120 2410.930 ;
        RECT 1800.540 2409.930 1800.800 2410.250 ;
        RECT 1802.840 2409.930 1803.100 2410.250 ;
        RECT 1790.170 2399.310 1792.000 2399.450 ;
        RECT 1801.210 2399.450 1801.490 2400.000 ;
        RECT 1802.900 2399.450 1803.040 2409.930 ;
        RECT 1813.880 2409.590 1814.140 2409.910 ;
        RECT 1801.210 2399.310 1803.040 2399.450 ;
        RECT 1812.250 2399.450 1812.530 2400.000 ;
        RECT 1813.940 2399.450 1814.080 2409.590 ;
        RECT 1824.920 2409.250 1825.180 2409.570 ;
        RECT 1812.250 2399.310 1814.080 2399.450 ;
        RECT 1823.290 2399.450 1823.570 2400.000 ;
        RECT 1824.980 2399.450 1825.120 2409.250 ;
        RECT 1835.040 2408.910 1835.300 2409.230 ;
        RECT 1823.290 2399.310 1825.120 2399.450 ;
        RECT 1834.330 2399.450 1834.610 2400.000 ;
        RECT 1835.100 2399.450 1835.240 2408.910 ;
        RECT 1847.000 2408.570 1847.260 2408.890 ;
        RECT 1834.330 2399.310 1835.240 2399.450 ;
        RECT 1845.370 2399.450 1845.650 2400.000 ;
        RECT 1847.060 2399.450 1847.200 2408.570 ;
        RECT 1858.040 2408.230 1858.300 2408.550 ;
        RECT 1845.370 2399.310 1847.200 2399.450 ;
        RECT 1856.410 2399.450 1856.690 2400.000 ;
        RECT 1858.100 2399.450 1858.240 2408.230 ;
        RECT 1856.410 2399.310 1858.240 2399.450 ;
        RECT 1865.920 2399.450 1866.060 2410.610 ;
        RECT 1867.450 2399.450 1867.730 2400.000 ;
        RECT 1865.920 2399.310 1867.730 2399.450 ;
        RECT 1876.960 2399.450 1877.100 2410.950 ;
        RECT 1878.490 2399.450 1878.770 2400.000 ;
        RECT 1876.960 2399.310 1878.770 2399.450 ;
        RECT 1888.000 2399.450 1888.140 2414.690 ;
        RECT 1898.120 2411.950 1898.260 2704.515 ;
        RECT 1898.060 2411.630 1898.320 2411.950 ;
        RECT 1898.580 2411.125 1898.720 3047.915 ;
        RECT 2087.110 3030.915 2087.390 3031.285 ;
        RECT 2083.890 2699.075 2084.170 2699.445 ;
        RECT 2083.960 2698.230 2084.100 2699.075 ;
        RECT 2048.940 2697.910 2049.200 2698.230 ;
        RECT 2083.900 2697.910 2084.160 2698.230 ;
        RECT 1993.280 2591.830 1993.540 2592.150 ;
        RECT 1979.940 2591.490 1980.200 2591.810 ;
        RECT 1966.140 2591.150 1966.400 2591.470 ;
        RECT 1959.240 2590.470 1959.500 2590.790 ;
        RECT 1898.980 2414.350 1899.240 2414.670 ;
        RECT 1898.510 2410.755 1898.790 2411.125 ;
        RECT 1889.530 2399.450 1889.810 2400.000 ;
        RECT 1888.000 2399.310 1889.810 2399.450 ;
        RECT 1899.040 2399.450 1899.180 2414.350 ;
        RECT 1911.400 2414.010 1911.660 2414.330 ;
        RECT 1911.460 2400.810 1911.600 2414.010 ;
        RECT 1920.600 2413.670 1920.860 2413.990 ;
        RECT 1911.460 2400.670 1911.830 2400.810 ;
        RECT 1911.690 2400.000 1911.830 2400.670 ;
        RECT 1900.570 2399.450 1900.850 2400.000 ;
        RECT 1899.040 2399.310 1900.850 2399.450 ;
        RECT 1779.130 2396.000 1779.410 2399.310 ;
        RECT 1790.170 2396.000 1790.450 2399.310 ;
        RECT 1801.210 2396.000 1801.490 2399.310 ;
        RECT 1812.250 2396.000 1812.530 2399.310 ;
        RECT 1823.290 2396.000 1823.570 2399.310 ;
        RECT 1834.330 2396.000 1834.610 2399.310 ;
        RECT 1845.370 2396.000 1845.650 2399.310 ;
        RECT 1856.410 2396.000 1856.690 2399.310 ;
        RECT 1867.450 2396.000 1867.730 2399.310 ;
        RECT 1878.490 2396.000 1878.770 2399.310 ;
        RECT 1889.530 2396.000 1889.810 2399.310 ;
        RECT 1900.570 2396.000 1900.850 2399.310 ;
        RECT 1911.610 2396.000 1911.890 2400.000 ;
        RECT 1920.660 2399.450 1920.800 2413.670 ;
        RECT 1959.300 2413.650 1959.440 2590.470 ;
        RECT 1932.100 2413.330 1932.360 2413.650 ;
        RECT 1956.940 2413.330 1957.200 2413.650 ;
        RECT 1959.240 2413.330 1959.500 2413.650 ;
        RECT 1922.190 2399.450 1922.470 2400.000 ;
        RECT 1920.660 2399.310 1922.470 2399.450 ;
        RECT 1932.160 2399.450 1932.300 2413.330 ;
        RECT 1932.560 2411.290 1932.820 2411.610 ;
        RECT 1942.670 2411.435 1942.950 2411.805 ;
        RECT 1932.620 2411.125 1932.760 2411.290 ;
        RECT 1932.550 2410.755 1932.830 2411.125 ;
        RECT 1933.230 2399.450 1933.510 2400.000 ;
        RECT 1932.160 2399.310 1933.510 2399.450 ;
        RECT 1942.740 2399.450 1942.880 2411.435 ;
        RECT 1945.900 2411.290 1946.160 2411.610 ;
        RECT 1945.960 2411.125 1946.100 2411.290 ;
        RECT 1945.890 2410.755 1946.170 2411.125 ;
        RECT 1944.270 2399.450 1944.550 2400.000 ;
        RECT 1942.740 2399.310 1944.550 2399.450 ;
        RECT 1922.190 2396.000 1922.470 2399.310 ;
        RECT 1933.230 2396.000 1933.510 2399.310 ;
        RECT 1944.270 2396.000 1944.550 2399.310 ;
        RECT 1955.310 2399.450 1955.590 2400.000 ;
        RECT 1957.000 2399.450 1957.140 2413.330 ;
        RECT 1966.200 2400.130 1966.340 2591.150 ;
        RECT 1980.000 2400.130 1980.140 2591.490 ;
        RECT 1993.340 2413.650 1993.480 2591.830 ;
        RECT 1990.060 2413.330 1990.320 2413.650 ;
        RECT 1993.280 2413.330 1993.540 2413.650 ;
        RECT 1966.200 2400.000 1966.570 2400.130 ;
        RECT 1966.200 2399.990 1966.630 2400.000 ;
        RECT 1955.310 2399.310 1957.140 2399.450 ;
        RECT 1955.310 2396.000 1955.590 2399.310 ;
        RECT 1966.350 2396.000 1966.630 2399.990 ;
        RECT 1977.390 2399.450 1977.670 2400.000 ;
        RECT 1979.080 2399.990 1980.140 2400.130 ;
        RECT 1979.080 2399.450 1979.220 2399.990 ;
        RECT 1977.390 2399.310 1979.220 2399.450 ;
        RECT 1988.430 2399.450 1988.710 2400.000 ;
        RECT 1990.120 2399.450 1990.260 2413.330 ;
        RECT 1997.880 2412.990 1998.140 2413.310 ;
        RECT 1988.430 2399.310 1990.260 2399.450 ;
        RECT 1997.940 2399.450 1998.080 2412.990 ;
        RECT 2049.000 2412.970 2049.140 2697.910 ;
        RECT 2008.920 2412.650 2009.180 2412.970 ;
        RECT 2045.260 2412.650 2045.520 2412.970 ;
        RECT 2048.940 2412.650 2049.200 2412.970 ;
        RECT 1999.470 2399.450 1999.750 2400.000 ;
        RECT 1997.940 2399.310 1999.750 2399.450 ;
        RECT 2008.980 2399.450 2009.120 2412.650 ;
        RECT 2019.960 2412.310 2020.220 2412.630 ;
        RECT 2010.510 2399.450 2010.790 2400.000 ;
        RECT 2008.980 2399.310 2010.790 2399.450 ;
        RECT 2020.020 2399.450 2020.160 2412.310 ;
        RECT 2031.000 2411.970 2031.260 2412.290 ;
        RECT 2021.550 2399.450 2021.830 2400.000 ;
        RECT 2020.020 2399.310 2021.830 2399.450 ;
        RECT 2031.060 2399.450 2031.200 2411.970 ;
        RECT 2032.590 2399.450 2032.870 2400.000 ;
        RECT 2031.060 2399.310 2032.870 2399.450 ;
        RECT 1977.390 2396.000 1977.670 2399.310 ;
        RECT 1988.430 2396.000 1988.710 2399.310 ;
        RECT 1999.470 2396.000 1999.750 2399.310 ;
        RECT 2010.510 2396.000 2010.790 2399.310 ;
        RECT 2021.550 2396.000 2021.830 2399.310 ;
        RECT 2032.590 2396.000 2032.870 2399.310 ;
        RECT 2043.630 2399.450 2043.910 2400.000 ;
        RECT 2045.320 2399.450 2045.460 2412.650 ;
        RECT 2086.660 2411.970 2086.920 2412.290 ;
        RECT 2076.080 2411.630 2076.340 2411.950 ;
        RECT 2067.340 2411.290 2067.600 2411.610 ;
        RECT 2053.080 2410.610 2053.340 2410.930 ;
        RECT 2043.630 2399.310 2045.460 2399.450 ;
        RECT 2053.140 2399.450 2053.280 2410.610 ;
        RECT 2054.670 2399.450 2054.950 2400.000 ;
        RECT 2053.140 2399.310 2054.950 2399.450 ;
        RECT 2043.630 2396.000 2043.910 2399.310 ;
        RECT 2054.670 2396.000 2054.950 2399.310 ;
        RECT 2065.710 2399.450 2065.990 2400.000 ;
        RECT 2067.400 2399.450 2067.540 2411.290 ;
        RECT 2065.710 2399.310 2067.540 2399.450 ;
        RECT 2065.710 2396.000 2065.990 2399.310 ;
        RECT 2076.140 2398.770 2076.280 2411.630 ;
        RECT 2076.750 2398.770 2077.030 2400.000 ;
        RECT 2086.720 2399.450 2086.860 2411.970 ;
        RECT 2087.180 2408.550 2087.320 3030.915 ;
        RECT 2087.570 3024.115 2087.850 3024.485 ;
        RECT 2087.640 2408.890 2087.780 3024.115 ;
        RECT 2088.030 3015.955 2088.310 3016.325 ;
        RECT 2088.100 2409.230 2088.240 3015.955 ;
        RECT 2088.490 3009.835 2088.770 3010.205 ;
        RECT 2088.560 2409.570 2088.700 3009.835 ;
        RECT 2088.950 3001.675 2089.230 3002.045 ;
        RECT 2089.020 2409.910 2089.160 3001.675 ;
        RECT 2089.410 2996.235 2089.690 2996.605 ;
        RECT 2089.480 2410.250 2089.620 2996.235 ;
        RECT 2089.870 2988.075 2090.150 2988.445 ;
        RECT 2089.940 2410.590 2090.080 2988.075 ;
        RECT 2090.330 2691.595 2090.610 2691.965 ;
        RECT 2090.400 2604.730 2090.540 2691.595 ;
      LAYER met2 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
      LAYER met2 ;
        RECT 2482.320 3049.645 2482.460 3051.850 ;
        RECT 2482.250 3049.275 2482.530 3049.645 ;
        RECT 2497.960 2747.725 2498.100 3063.750 ;
        RECT 2497.890 2747.355 2498.170 2747.725 ;
        RECT 2497.890 2709.955 2498.170 2710.325 ;
        RECT 2497.960 2704.885 2498.100 2709.955 ;
        RECT 2497.890 2704.515 2498.170 2704.885 ;
        RECT 2090.340 2604.410 2090.600 2604.730 ;
        RECT 2090.400 2411.125 2090.540 2604.410 ;
        RECT 2126.670 2598.435 2126.950 2598.805 ;
        RECT 2126.740 2590.790 2126.880 2598.435 ;
        RECT 2215.910 2593.675 2216.190 2594.045 ;
        RECT 2256.390 2593.675 2256.670 2594.045 ;
        RECT 2262.830 2593.675 2263.110 2594.045 ;
        RECT 2268.350 2593.675 2268.630 2594.045 ;
        RECT 2297.790 2593.675 2298.070 2594.045 ;
        RECT 2305.150 2593.675 2305.430 2594.045 ;
        RECT 2215.980 2593.510 2216.120 2593.675 ;
        RECT 2256.400 2593.530 2256.660 2593.675 ;
        RECT 2146.450 2592.995 2146.730 2593.365 ;
        RECT 2215.920 2593.190 2216.180 2593.510 ;
        RECT 2145.990 2591.635 2146.270 2592.005 ;
        RECT 2146.520 2591.810 2146.660 2592.995 ;
        RECT 2208.100 2592.850 2208.360 2593.170 ;
        RECT 2152.890 2592.315 2153.170 2592.685 ;
        RECT 2152.960 2592.150 2153.100 2592.315 ;
        RECT 2152.900 2591.830 2153.160 2592.150 ;
        RECT 2146.060 2591.470 2146.200 2591.635 ;
        RECT 2146.460 2591.490 2146.720 2591.810 ;
        RECT 2146.000 2591.150 2146.260 2591.470 ;
        RECT 2126.680 2590.470 2126.940 2590.790 ;
        RECT 2132.190 2590.275 2132.470 2590.645 ;
        RECT 2176.810 2590.275 2177.090 2590.645 ;
        RECT 2179.570 2590.275 2179.850 2590.645 ;
        RECT 2183.710 2590.275 2183.990 2590.645 ;
        RECT 2132.200 2590.130 2132.460 2590.275 ;
        RECT 2152.900 2589.790 2153.160 2590.110 ;
        RECT 2133.120 2414.350 2133.380 2414.670 ;
        RECT 2122.080 2412.990 2122.340 2413.310 ;
        RECT 2111.040 2412.650 2111.300 2412.970 ;
        RECT 2100.000 2412.310 2100.260 2412.630 ;
        RECT 2090.330 2410.755 2090.610 2411.125 ;
        RECT 2089.880 2410.270 2090.140 2410.590 ;
        RECT 2089.420 2409.930 2089.680 2410.250 ;
        RECT 2088.960 2409.590 2089.220 2409.910 ;
        RECT 2088.500 2409.250 2088.760 2409.570 ;
        RECT 2088.040 2408.910 2088.300 2409.230 ;
        RECT 2087.580 2408.570 2087.840 2408.890 ;
        RECT 2087.120 2408.230 2087.380 2408.550 ;
        RECT 2087.790 2399.450 2088.070 2400.000 ;
        RECT 2086.720 2399.310 2088.070 2399.450 ;
        RECT 2076.140 2398.630 2077.030 2398.770 ;
        RECT 2076.750 2396.000 2077.030 2398.630 ;
        RECT 2087.790 2396.000 2088.070 2399.310 ;
        RECT 2098.370 2399.450 2098.650 2400.000 ;
        RECT 2100.060 2399.450 2100.200 2412.310 ;
        RECT 2098.370 2399.310 2100.200 2399.450 ;
        RECT 2109.410 2399.450 2109.690 2400.000 ;
        RECT 2111.100 2399.450 2111.240 2412.650 ;
        RECT 2109.410 2399.310 2111.240 2399.450 ;
        RECT 2120.450 2399.450 2120.730 2400.000 ;
        RECT 2122.140 2399.450 2122.280 2412.990 ;
        RECT 2120.450 2399.310 2122.280 2399.450 ;
        RECT 2098.370 2396.000 2098.650 2399.310 ;
        RECT 2109.410 2396.000 2109.690 2399.310 ;
        RECT 2120.450 2396.000 2120.730 2399.310 ;
        RECT 2131.490 2398.090 2131.770 2400.000 ;
        RECT 2133.180 2398.090 2133.320 2414.350 ;
        RECT 2144.160 2410.950 2144.420 2411.270 ;
        RECT 2131.490 2397.950 2133.320 2398.090 ;
        RECT 2142.530 2399.450 2142.810 2400.000 ;
        RECT 2144.220 2399.450 2144.360 2410.950 ;
        RECT 2142.530 2399.310 2144.360 2399.450 ;
        RECT 2152.960 2399.450 2153.100 2589.790 ;
        RECT 2159.800 2589.450 2160.060 2589.770 ;
        RECT 2170.380 2589.450 2170.640 2589.770 ;
        RECT 2153.570 2399.450 2153.850 2400.000 ;
        RECT 2152.960 2399.310 2153.850 2399.450 ;
        RECT 2159.860 2399.450 2160.000 2589.450 ;
        RECT 2170.440 2589.285 2170.580 2589.450 ;
        RECT 2163.020 2588.770 2163.280 2589.090 ;
        RECT 2170.370 2588.915 2170.650 2589.285 ;
        RECT 2163.080 2588.605 2163.220 2588.770 ;
        RECT 2163.010 2588.235 2163.290 2588.605 ;
        RECT 2166.230 2588.235 2166.510 2588.605 ;
        RECT 2163.080 2411.610 2163.220 2588.235 ;
        RECT 2166.300 2415.010 2166.440 2588.235 ;
        RECT 2170.440 2573.530 2170.580 2588.915 ;
        RECT 2173.130 2588.235 2173.410 2588.605 ;
        RECT 2169.980 2573.390 2170.580 2573.530 ;
        RECT 2169.980 2560.045 2170.120 2573.390 ;
        RECT 2168.990 2559.675 2169.270 2560.045 ;
        RECT 2169.910 2559.675 2170.190 2560.045 ;
        RECT 2169.060 2511.910 2169.200 2559.675 ;
        RECT 2169.000 2511.590 2169.260 2511.910 ;
        RECT 2170.380 2511.590 2170.640 2511.910 ;
        RECT 2170.440 2476.970 2170.580 2511.590 ;
        RECT 2169.520 2476.830 2170.580 2476.970 ;
        RECT 2169.520 2463.290 2169.660 2476.830 ;
        RECT 2168.080 2462.970 2168.340 2463.290 ;
        RECT 2169.460 2462.970 2169.720 2463.290 ;
        RECT 2168.140 2415.205 2168.280 2462.970 ;
        RECT 2166.240 2414.690 2166.500 2415.010 ;
        RECT 2168.070 2414.835 2168.350 2415.205 ;
        RECT 2168.990 2414.835 2169.270 2415.205 ;
        RECT 2169.060 2411.950 2169.200 2414.835 ;
        RECT 2173.200 2414.330 2173.340 2588.235 ;
        RECT 2173.600 2587.750 2173.860 2588.070 ;
        RECT 2173.140 2414.010 2173.400 2414.330 ;
        RECT 2169.000 2411.630 2169.260 2411.950 ;
        RECT 2163.020 2411.290 2163.280 2411.610 ;
        RECT 2164.610 2399.450 2164.890 2400.000 ;
        RECT 2159.860 2399.310 2164.890 2399.450 ;
        RECT 2173.660 2399.450 2173.800 2587.750 ;
        RECT 2176.880 2412.290 2177.020 2590.275 ;
        RECT 2179.580 2590.130 2179.840 2590.275 ;
        RECT 2183.780 2590.110 2183.920 2590.275 ;
        RECT 2183.720 2589.790 2183.980 2590.110 ;
        RECT 2180.500 2589.110 2180.760 2589.430 ;
        RECT 2180.030 2588.235 2180.310 2588.605 ;
        RECT 2180.100 2413.650 2180.240 2588.235 ;
        RECT 2180.560 2414.410 2180.700 2589.110 ;
        RECT 2180.560 2414.270 2182.540 2414.410 ;
        RECT 2180.500 2413.670 2180.760 2413.990 ;
        RECT 2180.040 2413.330 2180.300 2413.650 ;
        RECT 2180.560 2412.630 2180.700 2413.670 ;
        RECT 2180.500 2412.310 2180.760 2412.630 ;
        RECT 2176.820 2411.970 2177.080 2412.290 ;
        RECT 2182.400 2400.130 2182.540 2414.270 ;
        RECT 2183.780 2413.990 2183.920 2589.790 ;
        RECT 2186.470 2589.595 2186.750 2589.965 ;
        RECT 2186.540 2589.430 2186.680 2589.595 ;
        RECT 2184.640 2589.110 2184.900 2589.430 ;
        RECT 2186.480 2589.110 2186.740 2589.430 ;
        RECT 2183.720 2413.670 2183.980 2413.990 ;
        RECT 2184.700 2412.970 2184.840 2589.110 ;
        RECT 2186.930 2588.235 2187.210 2588.605 ;
        RECT 2190.620 2588.430 2190.880 2588.750 ;
        RECT 2187.000 2413.990 2187.140 2588.235 ;
        RECT 2190.680 2587.925 2190.820 2588.430 ;
        RECT 2193.830 2588.235 2194.110 2588.605 ;
        RECT 2190.610 2587.555 2190.890 2587.925 ;
        RECT 2193.370 2587.555 2193.650 2587.925 ;
        RECT 2186.940 2413.670 2187.200 2413.990 ;
        RECT 2190.680 2413.310 2190.820 2587.555 ;
        RECT 2190.620 2412.990 2190.880 2413.310 ;
        RECT 2193.440 2412.970 2193.580 2587.555 ;
        RECT 2193.900 2413.310 2194.040 2588.235 ;
        RECT 2194.300 2588.090 2194.560 2588.410 ;
        RECT 2197.510 2588.235 2197.790 2588.605 ;
        RECT 2204.410 2588.235 2204.690 2588.605 ;
        RECT 2193.840 2412.990 2194.100 2413.310 ;
        RECT 2184.640 2412.650 2184.900 2412.970 ;
        RECT 2193.380 2412.650 2193.640 2412.970 ;
        RECT 2175.650 2399.450 2175.930 2400.000 ;
        RECT 2182.400 2399.990 2184.840 2400.130 ;
        RECT 2173.660 2399.310 2175.930 2399.450 ;
        RECT 2184.700 2399.450 2184.840 2399.990 ;
        RECT 2186.690 2399.450 2186.970 2400.000 ;
        RECT 2184.700 2399.310 2186.970 2399.450 ;
        RECT 2131.490 2396.000 2131.770 2397.950 ;
        RECT 2142.530 2396.000 2142.810 2399.310 ;
        RECT 2153.570 2396.000 2153.850 2399.310 ;
        RECT 2164.610 2396.000 2164.890 2399.310 ;
        RECT 2175.650 2396.000 2175.930 2399.310 ;
        RECT 2186.690 2396.000 2186.970 2399.310 ;
        RECT 2194.360 2398.770 2194.500 2588.090 ;
        RECT 2197.580 2588.070 2197.720 2588.235 ;
        RECT 2204.420 2588.090 2204.680 2588.235 ;
        RECT 2197.520 2587.750 2197.780 2588.070 ;
        RECT 2197.580 2414.670 2197.720 2587.750 ;
        RECT 2200.730 2587.555 2201.010 2587.925 ;
        RECT 2197.520 2414.350 2197.780 2414.670 ;
        RECT 2200.800 2412.290 2200.940 2587.555 ;
        RECT 2200.740 2411.970 2201.000 2412.290 ;
        RECT 2204.480 2411.270 2204.620 2588.090 ;
        RECT 2207.630 2587.555 2207.910 2587.925 ;
        RECT 2207.700 2411.950 2207.840 2587.555 ;
        RECT 2207.640 2411.630 2207.900 2411.950 ;
        RECT 2204.420 2410.950 2204.680 2411.270 ;
        RECT 2197.730 2398.770 2198.010 2400.000 ;
        RECT 2208.160 2399.450 2208.300 2592.850 ;
        RECT 2215.000 2592.510 2215.260 2592.830 ;
        RECT 2209.470 2590.955 2209.750 2591.325 ;
        RECT 2209.540 2589.090 2209.680 2590.955 ;
        RECT 2214.540 2590.810 2214.800 2591.130 ;
        RECT 2214.600 2589.090 2214.740 2590.810 ;
        RECT 2209.480 2588.770 2209.740 2589.090 ;
        RECT 2214.540 2588.770 2214.800 2589.090 ;
        RECT 2214.530 2587.555 2214.810 2587.925 ;
        RECT 2214.600 2412.630 2214.740 2587.555 ;
        RECT 2214.540 2412.310 2214.800 2412.630 ;
        RECT 2208.770 2399.450 2209.050 2400.000 ;
        RECT 2208.160 2399.310 2209.050 2399.450 ;
        RECT 2194.360 2398.630 2198.010 2398.770 ;
        RECT 2197.730 2396.000 2198.010 2398.630 ;
        RECT 2208.770 2396.000 2209.050 2399.310 ;
        RECT 2215.060 2398.770 2215.200 2592.510 ;
        RECT 2215.980 2589.770 2216.120 2593.190 ;
        RECT 2220.510 2592.995 2220.790 2593.365 ;
        RECT 2220.520 2592.850 2220.780 2592.995 ;
        RECT 2220.580 2590.450 2220.720 2592.850 ;
        RECT 2228.800 2592.170 2229.060 2592.490 ;
        RECT 2235.690 2592.315 2235.970 2592.685 ;
        RECT 2243.980 2592.510 2244.240 2592.830 ;
        RECT 2227.870 2590.955 2228.150 2591.325 ;
        RECT 2220.520 2590.130 2220.780 2590.450 ;
        RECT 2227.940 2590.110 2228.080 2590.955 ;
        RECT 2227.880 2589.790 2228.140 2590.110 ;
        RECT 2215.920 2589.450 2216.180 2589.770 ;
        RECT 2228.330 2588.235 2228.610 2588.605 ;
        RECT 2221.430 2587.555 2221.710 2587.925 ;
        RECT 2227.870 2587.555 2228.150 2587.925 ;
        RECT 2221.500 2411.610 2221.640 2587.555 ;
        RECT 2221.440 2411.290 2221.700 2411.610 ;
        RECT 2227.940 2408.890 2228.080 2587.555 ;
        RECT 2227.880 2408.570 2228.140 2408.890 ;
        RECT 2228.400 2408.550 2228.540 2588.235 ;
        RECT 2228.340 2408.230 2228.600 2408.550 ;
        RECT 2219.810 2398.770 2220.090 2400.000 ;
        RECT 2228.860 2399.450 2229.000 2592.170 ;
        RECT 2235.760 2592.150 2235.900 2592.315 ;
        RECT 2232.930 2591.635 2233.210 2592.005 ;
        RECT 2235.700 2591.830 2235.960 2592.150 ;
        RECT 2244.040 2592.005 2244.180 2592.510 ;
        RECT 2249.490 2592.315 2249.770 2592.685 ;
        RECT 2249.500 2592.170 2249.760 2592.315 ;
        RECT 2232.940 2591.490 2233.200 2591.635 ;
        RECT 2233.000 2589.430 2233.140 2591.490 ;
        RECT 2232.940 2589.110 2233.200 2589.430 ;
        RECT 2235.760 2588.750 2235.900 2591.830 ;
        RECT 2243.970 2591.635 2244.250 2592.005 ;
        RECT 2235.700 2588.430 2235.960 2588.750 ;
        RECT 2244.040 2588.070 2244.180 2591.635 ;
        RECT 2249.560 2588.410 2249.700 2592.170 ;
        RECT 2256.460 2591.130 2256.600 2593.530 ;
        RECT 2262.900 2593.510 2263.040 2593.675 ;
        RECT 2262.840 2593.190 2263.100 2593.510 ;
        RECT 2268.420 2593.170 2268.560 2593.675 ;
        RECT 2297.800 2593.530 2298.060 2593.675 ;
        RECT 2305.220 2593.510 2305.360 2593.675 ;
        RECT 2268.360 2592.850 2268.620 2593.170 ;
        RECT 2291.810 2592.995 2292.090 2593.365 ;
        RECT 2297.790 2592.995 2298.070 2593.365 ;
        RECT 2305.160 2593.190 2305.420 2593.510 ;
        RECT 2311.590 2592.995 2311.870 2593.365 ;
        RECT 2332.290 2592.995 2332.570 2593.365 ;
        RECT 2291.880 2592.830 2292.020 2592.995 ;
        RECT 2280.310 2592.315 2280.590 2592.685 ;
        RECT 2285.370 2592.315 2285.650 2592.685 ;
        RECT 2291.820 2592.510 2292.080 2592.830 ;
        RECT 2276.170 2591.635 2276.450 2592.005 ;
        RECT 2280.380 2591.810 2280.520 2592.315 ;
        RECT 2285.440 2592.150 2285.580 2592.315 ;
        RECT 2297.860 2592.150 2298.000 2592.995 ;
        RECT 2311.600 2592.850 2311.860 2592.995 ;
        RECT 2332.360 2592.830 2332.500 2592.995 ;
        RECT 2332.300 2592.510 2332.560 2592.830 ;
        RECT 2339.190 2592.315 2339.470 2592.685 ;
        RECT 2339.260 2592.150 2339.400 2592.315 ;
        RECT 2285.380 2591.830 2285.640 2592.150 ;
        RECT 2297.800 2591.830 2298.060 2592.150 ;
        RECT 2276.240 2591.470 2276.380 2591.635 ;
        RECT 2280.320 2591.490 2280.580 2591.810 ;
        RECT 2318.490 2591.635 2318.770 2592.005 ;
        RECT 2332.290 2591.635 2332.570 2592.005 ;
        RECT 2339.200 2591.830 2339.460 2592.150 ;
        RECT 2276.180 2591.150 2276.440 2591.470 ;
        RECT 2256.400 2590.810 2256.660 2591.130 ;
        RECT 2276.240 2590.110 2276.380 2591.150 ;
        RECT 2280.380 2591.130 2280.520 2591.490 ;
        RECT 2318.560 2591.470 2318.700 2591.635 ;
        RECT 2332.300 2591.490 2332.560 2591.635 ;
        RECT 2318.500 2591.150 2318.760 2591.470 ;
        RECT 2280.320 2590.810 2280.580 2591.130 ;
        RECT 2325.390 2590.955 2325.670 2591.325 ;
        RECT 2325.400 2590.810 2325.660 2590.955 ;
        RECT 2276.180 2589.790 2276.440 2590.110 ;
        RECT 2249.500 2588.090 2249.760 2588.410 ;
        RECT 2269.270 2588.235 2269.550 2588.605 ;
        RECT 2303.770 2588.235 2304.050 2588.605 ;
        RECT 2345.170 2588.235 2345.450 2588.605 ;
        RECT 2235.230 2587.555 2235.510 2587.925 ;
        RECT 2242.130 2587.555 2242.410 2587.925 ;
        RECT 2243.980 2587.750 2244.240 2588.070 ;
        RECT 2249.030 2587.555 2249.310 2587.925 ;
        RECT 2255.930 2587.555 2256.210 2587.925 ;
        RECT 2262.830 2587.555 2263.110 2587.925 ;
        RECT 2235.300 2409.570 2235.440 2587.555 ;
        RECT 2240.300 2414.690 2240.560 2415.010 ;
        RECT 2235.240 2409.250 2235.500 2409.570 ;
        RECT 2230.850 2399.450 2231.130 2400.000 ;
        RECT 2228.860 2399.310 2231.130 2399.450 ;
        RECT 2240.360 2399.450 2240.500 2414.690 ;
        RECT 2242.200 2409.230 2242.340 2587.555 ;
        RECT 2249.100 2409.910 2249.240 2587.555 ;
        RECT 2251.340 2414.010 2251.600 2414.330 ;
        RECT 2249.040 2409.590 2249.300 2409.910 ;
        RECT 2242.140 2408.910 2242.400 2409.230 ;
        RECT 2241.890 2399.450 2242.170 2400.000 ;
        RECT 2240.360 2399.310 2242.170 2399.450 ;
        RECT 2251.400 2399.450 2251.540 2414.010 ;
        RECT 2256.000 2410.250 2256.140 2587.555 ;
        RECT 2262.900 2410.590 2263.040 2587.555 ;
        RECT 2263.300 2413.330 2263.560 2413.650 ;
        RECT 2262.840 2410.270 2263.100 2410.590 ;
        RECT 2255.940 2409.930 2256.200 2410.250 ;
        RECT 2263.360 2400.810 2263.500 2413.330 ;
        RECT 2269.340 2410.930 2269.480 2588.235 ;
        RECT 2269.730 2587.555 2270.010 2587.925 ;
        RECT 2276.630 2587.555 2276.910 2587.925 ;
        RECT 2283.530 2587.555 2283.810 2587.925 ;
        RECT 2290.430 2587.555 2290.710 2587.925 ;
        RECT 2297.330 2587.555 2297.610 2587.925 ;
        RECT 2269.800 2411.270 2269.940 2587.555 ;
        RECT 2276.700 2415.010 2276.840 2587.555 ;
        RECT 2276.640 2414.690 2276.900 2415.010 ;
        RECT 2283.600 2414.670 2283.740 2587.555 ;
        RECT 2283.540 2414.350 2283.800 2414.670 ;
        RECT 2290.500 2414.330 2290.640 2587.555 ;
        RECT 2290.440 2414.010 2290.700 2414.330 ;
        RECT 2297.400 2413.990 2297.540 2587.555 ;
        RECT 2272.960 2413.670 2273.220 2413.990 ;
        RECT 2297.340 2413.670 2297.600 2413.990 ;
        RECT 2269.740 2410.950 2270.000 2411.270 ;
        RECT 2269.280 2410.610 2269.540 2410.930 ;
        RECT 2263.360 2400.670 2263.730 2400.810 ;
        RECT 2263.590 2400.000 2263.730 2400.670 ;
        RECT 2252.930 2399.450 2253.210 2400.000 ;
        RECT 2251.400 2399.310 2253.210 2399.450 ;
        RECT 2215.060 2398.630 2220.090 2398.770 ;
        RECT 2219.810 2396.000 2220.090 2398.630 ;
        RECT 2230.850 2396.000 2231.130 2399.310 ;
        RECT 2241.890 2396.000 2242.170 2399.310 ;
        RECT 2252.930 2396.000 2253.210 2399.310 ;
        RECT 2263.510 2396.000 2263.790 2400.000 ;
        RECT 2273.020 2399.450 2273.160 2413.670 ;
        RECT 2303.840 2413.650 2303.980 2588.235 ;
        RECT 2304.230 2587.555 2304.510 2587.925 ;
        RECT 2311.130 2587.555 2311.410 2587.925 ;
        RECT 2318.030 2587.555 2318.310 2587.925 ;
        RECT 2324.930 2587.555 2325.210 2587.925 ;
        RECT 2331.830 2587.555 2332.110 2587.925 ;
        RECT 2338.730 2587.555 2339.010 2587.925 ;
        RECT 2303.780 2413.330 2304.040 2413.650 ;
        RECT 2284.460 2412.990 2284.720 2413.310 ;
        RECT 2274.550 2399.450 2274.830 2400.000 ;
        RECT 2273.020 2399.310 2274.830 2399.450 ;
        RECT 2284.520 2399.450 2284.660 2412.990 ;
        RECT 2304.300 2412.970 2304.440 2587.555 ;
        RECT 2311.200 2413.310 2311.340 2587.555 ;
        RECT 2311.140 2412.990 2311.400 2413.310 ;
        RECT 2295.040 2412.650 2295.300 2412.970 ;
        RECT 2304.240 2412.650 2304.500 2412.970 ;
        RECT 2285.590 2399.450 2285.870 2400.000 ;
        RECT 2284.520 2399.310 2285.870 2399.450 ;
        RECT 2295.100 2399.450 2295.240 2412.650 ;
        RECT 2318.100 2412.370 2318.240 2587.555 ;
        RECT 2325.000 2412.630 2325.140 2587.555 ;
        RECT 2318.100 2412.290 2319.620 2412.370 ;
        RECT 2324.940 2412.310 2325.200 2412.630 ;
        RECT 2306.080 2411.970 2306.340 2412.290 ;
        RECT 2318.100 2412.230 2319.680 2412.290 ;
        RECT 2319.420 2411.970 2319.680 2412.230 ;
        RECT 2296.630 2399.450 2296.910 2400.000 ;
        RECT 2295.100 2399.310 2296.910 2399.450 ;
        RECT 2306.140 2399.450 2306.280 2411.970 ;
        RECT 2331.900 2411.950 2332.040 2587.555 ;
        RECT 2338.800 2412.485 2338.940 2587.555 ;
        RECT 2338.730 2412.115 2339.010 2412.485 ;
        RECT 2318.500 2411.630 2318.760 2411.950 ;
        RECT 2328.160 2411.630 2328.420 2411.950 ;
        RECT 2331.840 2411.630 2332.100 2411.950 ;
        RECT 2318.560 2400.810 2318.700 2411.630 ;
        RECT 2318.560 2400.670 2318.930 2400.810 ;
        RECT 2318.790 2400.000 2318.930 2400.670 ;
        RECT 2307.670 2399.450 2307.950 2400.000 ;
        RECT 2306.140 2399.310 2307.950 2399.450 ;
        RECT 2274.550 2396.000 2274.830 2399.310 ;
        RECT 2285.590 2396.000 2285.870 2399.310 ;
        RECT 2296.630 2396.000 2296.910 2399.310 ;
        RECT 2307.670 2396.000 2307.950 2399.310 ;
        RECT 2318.710 2396.000 2318.990 2400.000 ;
        RECT 2328.220 2399.450 2328.360 2411.630 ;
        RECT 2345.240 2411.610 2345.380 2588.235 ;
        RECT 2345.630 2587.555 2345.910 2587.925 ;
        RECT 2345.700 2411.805 2345.840 2587.555 ;
        RECT 2449.600 2414.690 2449.860 2415.010 ;
        RECT 2340.120 2411.290 2340.380 2411.610 ;
        RECT 2345.180 2411.290 2345.440 2411.610 ;
        RECT 2345.630 2411.435 2345.910 2411.805 ;
        RECT 2329.750 2399.450 2330.030 2400.000 ;
        RECT 2328.220 2399.310 2330.030 2399.450 ;
        RECT 2340.180 2399.450 2340.320 2411.290 ;
        RECT 2438.100 2410.950 2438.360 2411.270 ;
        RECT 2428.900 2410.610 2429.160 2410.930 ;
        RECT 2416.480 2410.270 2416.740 2410.590 ;
        RECT 2405.440 2409.930 2405.700 2410.250 ;
        RECT 2394.400 2409.590 2394.660 2409.910 ;
        RECT 2373.700 2409.250 2373.960 2409.570 ;
        RECT 2361.280 2408.570 2361.540 2408.890 ;
        RECT 2350.240 2408.230 2350.500 2408.550 ;
        RECT 2340.790 2399.450 2341.070 2400.000 ;
        RECT 2340.180 2399.310 2341.070 2399.450 ;
        RECT 2350.300 2399.450 2350.440 2408.230 ;
        RECT 2351.830 2399.450 2352.110 2400.000 ;
        RECT 2350.300 2399.310 2352.110 2399.450 ;
        RECT 2361.340 2399.450 2361.480 2408.570 ;
        RECT 2373.760 2400.810 2373.900 2409.250 ;
        RECT 2383.360 2408.910 2383.620 2409.230 ;
        RECT 2373.760 2400.670 2374.130 2400.810 ;
        RECT 2373.990 2400.000 2374.130 2400.670 ;
        RECT 2362.870 2399.450 2363.150 2400.000 ;
        RECT 2361.340 2399.310 2363.150 2399.450 ;
        RECT 2329.750 2396.000 2330.030 2399.310 ;
        RECT 2340.790 2396.000 2341.070 2399.310 ;
        RECT 2351.830 2396.000 2352.110 2399.310 ;
        RECT 2362.870 2396.000 2363.150 2399.310 ;
        RECT 2373.910 2396.000 2374.190 2400.000 ;
        RECT 2383.420 2399.450 2383.560 2408.910 ;
        RECT 2384.950 2399.450 2385.230 2400.000 ;
        RECT 2383.420 2399.310 2385.230 2399.450 ;
        RECT 2394.460 2399.450 2394.600 2409.590 ;
        RECT 2395.990 2399.450 2396.270 2400.000 ;
        RECT 2394.460 2399.310 2396.270 2399.450 ;
        RECT 2405.500 2399.450 2405.640 2409.930 ;
        RECT 2407.030 2399.450 2407.310 2400.000 ;
        RECT 2405.500 2399.310 2407.310 2399.450 ;
        RECT 2416.540 2399.450 2416.680 2410.270 ;
        RECT 2428.960 2400.810 2429.100 2410.610 ;
        RECT 2428.960 2400.670 2429.330 2400.810 ;
        RECT 2429.190 2400.000 2429.330 2400.670 ;
        RECT 2418.070 2399.450 2418.350 2400.000 ;
        RECT 2416.540 2399.310 2418.350 2399.450 ;
        RECT 2384.950 2396.000 2385.230 2399.310 ;
        RECT 2395.990 2396.000 2396.270 2399.310 ;
        RECT 2407.030 2396.000 2407.310 2399.310 ;
        RECT 2418.070 2396.000 2418.350 2399.310 ;
        RECT 2429.110 2396.000 2429.390 2400.000 ;
        RECT 2438.160 2399.450 2438.300 2410.950 ;
        RECT 2439.690 2399.450 2439.970 2400.000 ;
        RECT 2438.160 2399.310 2439.970 2399.450 ;
        RECT 2449.660 2399.450 2449.800 2414.690 ;
        RECT 2460.180 2414.350 2460.440 2414.670 ;
        RECT 2450.730 2399.450 2451.010 2400.000 ;
        RECT 2449.660 2399.310 2451.010 2399.450 ;
        RECT 2460.240 2399.450 2460.380 2414.350 ;
        RECT 2471.220 2414.010 2471.480 2414.330 ;
        RECT 2461.770 2399.450 2462.050 2400.000 ;
        RECT 2460.240 2399.310 2462.050 2399.450 ;
        RECT 2471.280 2399.450 2471.420 2414.010 ;
        RECT 2482.260 2413.670 2482.520 2413.990 ;
        RECT 2472.810 2399.450 2473.090 2400.000 ;
        RECT 2471.280 2399.310 2473.090 2399.450 ;
        RECT 2482.320 2399.450 2482.460 2413.670 ;
        RECT 2493.300 2413.330 2493.560 2413.650 ;
        RECT 2483.850 2399.450 2484.130 2400.000 ;
        RECT 2482.320 2399.310 2484.130 2399.450 ;
        RECT 2493.360 2399.450 2493.500 2413.330 ;
        RECT 2515.380 2412.990 2515.640 2413.310 ;
        RECT 2504.800 2412.650 2505.060 2412.970 ;
        RECT 2494.890 2399.450 2495.170 2400.000 ;
        RECT 2493.360 2399.310 2495.170 2399.450 ;
        RECT 2504.860 2399.450 2505.000 2412.650 ;
        RECT 2505.930 2399.450 2506.210 2400.000 ;
        RECT 2504.860 2399.310 2506.210 2399.450 ;
        RECT 2515.440 2399.450 2515.580 2412.990 ;
        RECT 2537.460 2412.310 2537.720 2412.630 ;
        RECT 2526.420 2411.970 2526.680 2412.290 ;
        RECT 2516.970 2399.450 2517.250 2400.000 ;
        RECT 2515.440 2399.310 2517.250 2399.450 ;
        RECT 2526.480 2399.450 2526.620 2411.970 ;
        RECT 2528.010 2399.450 2528.290 2400.000 ;
        RECT 2526.480 2399.310 2528.290 2399.450 ;
        RECT 2537.520 2399.450 2537.660 2412.310 ;
        RECT 2559.990 2412.115 2560.270 2412.485 ;
        RECT 2548.500 2411.630 2548.760 2411.950 ;
        RECT 2539.050 2399.450 2539.330 2400.000 ;
        RECT 2537.520 2399.310 2539.330 2399.450 ;
        RECT 2548.560 2399.450 2548.700 2411.630 ;
        RECT 2550.090 2399.450 2550.370 2400.000 ;
        RECT 2548.560 2399.310 2550.370 2399.450 ;
        RECT 2560.060 2399.450 2560.200 2412.115 ;
        RECT 2570.580 2411.290 2570.840 2411.610 ;
        RECT 2581.610 2411.435 2581.890 2411.805 ;
        RECT 2561.130 2399.450 2561.410 2400.000 ;
        RECT 2560.060 2399.310 2561.410 2399.450 ;
        RECT 2570.640 2399.450 2570.780 2411.290 ;
        RECT 2572.170 2399.450 2572.450 2400.000 ;
        RECT 2570.640 2399.310 2572.450 2399.450 ;
        RECT 2581.680 2399.450 2581.820 2411.435 ;
        RECT 2592.650 2410.755 2592.930 2411.125 ;
        RECT 2583.210 2399.450 2583.490 2400.000 ;
        RECT 2581.680 2399.310 2583.490 2399.450 ;
        RECT 2592.720 2399.450 2592.860 2410.755 ;
        RECT 2594.250 2399.450 2594.530 2400.000 ;
        RECT 2592.720 2399.310 2594.530 2399.450 ;
        RECT 2439.690 2396.000 2439.970 2399.310 ;
        RECT 2450.730 2396.000 2451.010 2399.310 ;
        RECT 2461.770 2396.000 2462.050 2399.310 ;
        RECT 2472.810 2396.000 2473.090 2399.310 ;
        RECT 2483.850 2396.000 2484.130 2399.310 ;
        RECT 2494.890 2396.000 2495.170 2399.310 ;
        RECT 2505.930 2396.000 2506.210 2399.310 ;
        RECT 2516.970 2396.000 2517.250 2399.310 ;
        RECT 2528.010 2396.000 2528.290 2399.310 ;
        RECT 2539.050 2396.000 2539.330 2399.310 ;
        RECT 2550.090 2396.000 2550.370 2399.310 ;
        RECT 2561.130 2396.000 2561.410 2399.310 ;
        RECT 2572.170 2396.000 2572.450 2399.310 ;
        RECT 2583.210 2396.000 2583.490 2399.310 ;
        RECT 2594.250 2396.000 2594.530 2399.310 ;
      LAYER met2 ;
        RECT 1404.690 2395.720 1404.870 2396.000 ;
        RECT 1405.710 2395.720 1415.450 2396.000 ;
        RECT 1416.290 2395.720 1426.490 2396.000 ;
        RECT 1427.330 2395.720 1437.530 2396.000 ;
        RECT 1438.370 2395.720 1448.570 2396.000 ;
        RECT 1449.410 2395.720 1459.610 2396.000 ;
        RECT 1460.450 2395.720 1470.650 2396.000 ;
        RECT 1471.490 2395.720 1481.690 2396.000 ;
        RECT 1482.530 2395.720 1492.730 2396.000 ;
        RECT 1493.570 2395.720 1503.770 2396.000 ;
        RECT 1504.610 2395.720 1514.810 2396.000 ;
        RECT 1515.650 2395.720 1525.850 2396.000 ;
        RECT 1526.690 2395.720 1536.890 2396.000 ;
        RECT 1537.730 2395.720 1547.930 2396.000 ;
        RECT 1548.770 2395.720 1558.970 2396.000 ;
        RECT 1559.810 2395.720 1570.010 2396.000 ;
        RECT 1570.850 2395.720 1580.590 2396.000 ;
        RECT 1581.430 2395.720 1591.630 2396.000 ;
        RECT 1592.470 2395.720 1602.670 2396.000 ;
        RECT 1603.510 2395.720 1613.710 2396.000 ;
        RECT 1614.550 2395.720 1624.750 2396.000 ;
        RECT 1625.590 2395.720 1635.790 2396.000 ;
        RECT 1636.630 2395.720 1646.830 2396.000 ;
        RECT 1647.670 2395.720 1657.870 2396.000 ;
        RECT 1658.710 2395.720 1668.910 2396.000 ;
        RECT 1669.750 2395.720 1679.950 2396.000 ;
        RECT 1680.790 2395.720 1690.990 2396.000 ;
        RECT 1691.830 2395.720 1702.030 2396.000 ;
        RECT 1702.870 2395.720 1713.070 2396.000 ;
        RECT 1713.910 2395.720 1724.110 2396.000 ;
        RECT 1724.950 2395.720 1735.150 2396.000 ;
        RECT 1735.990 2395.720 1746.190 2396.000 ;
        RECT 1747.030 2395.720 1756.770 2396.000 ;
        RECT 1757.610 2395.720 1767.810 2396.000 ;
        RECT 1768.650 2395.720 1778.850 2396.000 ;
        RECT 1779.690 2395.720 1789.890 2396.000 ;
        RECT 1790.730 2395.720 1800.930 2396.000 ;
        RECT 1801.770 2395.720 1811.970 2396.000 ;
        RECT 1812.810 2395.720 1823.010 2396.000 ;
        RECT 1823.850 2395.720 1834.050 2396.000 ;
        RECT 1834.890 2395.720 1845.090 2396.000 ;
        RECT 1845.930 2395.720 1856.130 2396.000 ;
        RECT 1856.970 2395.720 1867.170 2396.000 ;
        RECT 1868.010 2395.720 1878.210 2396.000 ;
        RECT 1879.050 2395.720 1889.250 2396.000 ;
        RECT 1890.090 2395.720 1900.290 2396.000 ;
        RECT 1901.130 2395.720 1911.330 2396.000 ;
        RECT 1912.170 2395.720 1921.910 2396.000 ;
        RECT 1922.750 2395.720 1932.950 2396.000 ;
        RECT 1933.790 2395.720 1943.990 2396.000 ;
        RECT 1944.830 2395.720 1955.030 2396.000 ;
        RECT 1955.870 2395.720 1966.070 2396.000 ;
        RECT 1966.910 2395.720 1977.110 2396.000 ;
        RECT 1977.950 2395.720 1988.150 2396.000 ;
        RECT 1988.990 2395.720 1999.190 2396.000 ;
        RECT 2000.030 2395.720 2010.230 2396.000 ;
        RECT 2011.070 2395.720 2021.270 2396.000 ;
        RECT 2022.110 2395.720 2032.310 2396.000 ;
        RECT 2033.150 2395.720 2043.350 2396.000 ;
        RECT 2044.190 2395.720 2054.390 2396.000 ;
        RECT 2055.230 2395.720 2065.430 2396.000 ;
        RECT 2066.270 2395.720 2076.470 2396.000 ;
        RECT 2077.310 2395.720 2087.510 2396.000 ;
        RECT 2088.350 2395.720 2098.090 2396.000 ;
        RECT 2098.930 2395.720 2109.130 2396.000 ;
        RECT 2109.970 2395.720 2120.170 2396.000 ;
        RECT 2121.010 2395.720 2131.210 2396.000 ;
        RECT 2132.050 2395.720 2142.250 2396.000 ;
        RECT 2143.090 2395.720 2153.290 2396.000 ;
        RECT 2154.130 2395.720 2164.330 2396.000 ;
        RECT 2165.170 2395.720 2175.370 2396.000 ;
        RECT 2176.210 2395.720 2186.410 2396.000 ;
        RECT 2187.250 2395.720 2197.450 2396.000 ;
        RECT 2198.290 2395.720 2208.490 2396.000 ;
        RECT 2209.330 2395.720 2219.530 2396.000 ;
        RECT 2220.370 2395.720 2230.570 2396.000 ;
        RECT 2231.410 2395.720 2241.610 2396.000 ;
        RECT 2242.450 2395.720 2252.650 2396.000 ;
        RECT 2253.490 2395.720 2263.230 2396.000 ;
        RECT 2264.070 2395.720 2274.270 2396.000 ;
        RECT 2275.110 2395.720 2285.310 2396.000 ;
        RECT 2286.150 2395.720 2296.350 2396.000 ;
        RECT 2297.190 2395.720 2307.390 2396.000 ;
        RECT 2308.230 2395.720 2318.430 2396.000 ;
        RECT 2319.270 2395.720 2329.470 2396.000 ;
        RECT 2330.310 2395.720 2340.510 2396.000 ;
        RECT 2341.350 2395.720 2351.550 2396.000 ;
        RECT 2352.390 2395.720 2362.590 2396.000 ;
        RECT 2363.430 2395.720 2373.630 2396.000 ;
        RECT 2374.470 2395.720 2384.670 2396.000 ;
        RECT 2385.510 2395.720 2395.710 2396.000 ;
        RECT 2396.550 2395.720 2406.750 2396.000 ;
        RECT 2407.590 2395.720 2417.790 2396.000 ;
        RECT 2418.630 2395.720 2428.830 2396.000 ;
        RECT 2429.670 2395.720 2439.410 2396.000 ;
        RECT 2440.250 2395.720 2450.450 2396.000 ;
        RECT 2451.290 2395.720 2461.490 2396.000 ;
        RECT 2462.330 2395.720 2472.530 2396.000 ;
        RECT 2473.370 2395.720 2483.570 2396.000 ;
        RECT 2484.410 2395.720 2494.610 2396.000 ;
        RECT 2495.450 2395.720 2505.650 2396.000 ;
        RECT 2506.490 2395.720 2516.690 2396.000 ;
        RECT 2517.530 2395.720 2527.730 2396.000 ;
        RECT 2528.570 2395.720 2538.770 2396.000 ;
        RECT 2539.610 2395.720 2549.810 2396.000 ;
        RECT 2550.650 2395.720 2560.850 2396.000 ;
        RECT 2561.690 2395.720 2571.890 2396.000 ;
        RECT 2572.730 2395.720 2582.930 2396.000 ;
        RECT 2583.770 2395.720 2593.970 2396.000 ;
        RECT 2594.810 2395.720 2594.990 2396.000 ;
        RECT 1404.690 1204.280 2594.990 2395.720 ;
        RECT 1404.690 1204.000 1404.870 1204.280 ;
        RECT 1405.710 1204.000 1415.450 1204.280 ;
        RECT 1416.290 1204.000 1426.490 1204.280 ;
        RECT 1427.330 1204.000 1437.530 1204.280 ;
        RECT 1438.370 1204.000 1448.570 1204.280 ;
        RECT 1449.410 1204.000 1459.610 1204.280 ;
        RECT 1460.450 1204.000 1470.650 1204.280 ;
        RECT 1471.490 1204.000 1481.690 1204.280 ;
        RECT 1482.530 1204.000 1492.730 1204.280 ;
        RECT 1493.570 1204.000 1503.770 1204.280 ;
        RECT 1504.610 1204.000 1514.810 1204.280 ;
        RECT 1515.650 1204.000 1525.850 1204.280 ;
        RECT 1526.690 1204.000 1536.890 1204.280 ;
        RECT 1537.730 1204.000 1547.930 1204.280 ;
        RECT 1548.770 1204.000 1558.970 1204.280 ;
        RECT 1559.810 1204.000 1570.010 1204.280 ;
        RECT 1570.850 1204.000 1580.590 1204.280 ;
        RECT 1581.430 1204.000 1591.630 1204.280 ;
        RECT 1592.470 1204.000 1602.670 1204.280 ;
        RECT 1603.510 1204.000 1613.710 1204.280 ;
        RECT 1614.550 1204.000 1624.750 1204.280 ;
        RECT 1625.590 1204.000 1635.790 1204.280 ;
        RECT 1636.630 1204.000 1646.830 1204.280 ;
        RECT 1647.670 1204.000 1657.870 1204.280 ;
        RECT 1658.710 1204.000 1668.910 1204.280 ;
        RECT 1669.750 1204.000 1679.950 1204.280 ;
        RECT 1680.790 1204.000 1690.990 1204.280 ;
        RECT 1691.830 1204.000 1702.030 1204.280 ;
        RECT 1702.870 1204.000 1713.070 1204.280 ;
        RECT 1713.910 1204.000 1724.110 1204.280 ;
        RECT 1724.950 1204.000 1735.150 1204.280 ;
        RECT 1735.990 1204.000 1746.190 1204.280 ;
        RECT 1747.030 1204.000 1756.770 1204.280 ;
        RECT 1757.610 1204.000 1767.810 1204.280 ;
        RECT 1768.650 1204.000 1778.850 1204.280 ;
        RECT 1779.690 1204.000 1789.890 1204.280 ;
        RECT 1790.730 1204.000 1800.930 1204.280 ;
        RECT 1801.770 1204.000 1811.970 1204.280 ;
        RECT 1812.810 1204.000 1823.010 1204.280 ;
        RECT 1823.850 1204.000 1834.050 1204.280 ;
        RECT 1834.890 1204.000 1845.090 1204.280 ;
        RECT 1845.930 1204.000 1856.130 1204.280 ;
        RECT 1856.970 1204.000 1867.170 1204.280 ;
        RECT 1868.010 1204.000 1878.210 1204.280 ;
        RECT 1879.050 1204.000 1889.250 1204.280 ;
        RECT 1890.090 1204.000 1900.290 1204.280 ;
        RECT 1901.130 1204.000 1911.330 1204.280 ;
        RECT 1912.170 1204.000 1921.910 1204.280 ;
        RECT 1922.750 1204.000 1932.950 1204.280 ;
        RECT 1933.790 1204.000 1943.990 1204.280 ;
        RECT 1944.830 1204.000 1955.030 1204.280 ;
        RECT 1955.870 1204.000 1966.070 1204.280 ;
        RECT 1966.910 1204.000 1977.110 1204.280 ;
        RECT 1977.950 1204.000 1988.150 1204.280 ;
        RECT 1988.990 1204.000 1999.190 1204.280 ;
        RECT 2000.030 1204.000 2010.230 1204.280 ;
        RECT 2011.070 1204.000 2021.270 1204.280 ;
        RECT 2022.110 1204.000 2032.310 1204.280 ;
        RECT 2033.150 1204.000 2043.350 1204.280 ;
        RECT 2044.190 1204.000 2054.390 1204.280 ;
        RECT 2055.230 1204.000 2065.430 1204.280 ;
        RECT 2066.270 1204.000 2076.470 1204.280 ;
        RECT 2077.310 1204.000 2087.510 1204.280 ;
        RECT 2088.350 1204.000 2098.090 1204.280 ;
        RECT 2098.930 1204.000 2109.130 1204.280 ;
        RECT 2109.970 1204.000 2120.170 1204.280 ;
        RECT 2121.010 1204.000 2131.210 1204.280 ;
        RECT 2132.050 1204.000 2142.250 1204.280 ;
        RECT 2143.090 1204.000 2153.290 1204.280 ;
        RECT 2154.130 1204.000 2164.330 1204.280 ;
        RECT 2165.170 1204.000 2175.370 1204.280 ;
        RECT 2176.210 1204.000 2186.410 1204.280 ;
        RECT 2187.250 1204.000 2197.450 1204.280 ;
        RECT 2198.290 1204.000 2208.490 1204.280 ;
        RECT 2209.330 1204.000 2219.530 1204.280 ;
        RECT 2220.370 1204.000 2230.570 1204.280 ;
        RECT 2231.410 1204.000 2241.610 1204.280 ;
        RECT 2242.450 1204.000 2252.650 1204.280 ;
        RECT 2253.490 1204.000 2263.230 1204.280 ;
        RECT 2264.070 1204.000 2274.270 1204.280 ;
        RECT 2275.110 1204.000 2285.310 1204.280 ;
        RECT 2286.150 1204.000 2296.350 1204.280 ;
        RECT 2297.190 1204.000 2307.390 1204.280 ;
        RECT 2308.230 1204.000 2318.430 1204.280 ;
        RECT 2319.270 1204.000 2329.470 1204.280 ;
        RECT 2330.310 1204.000 2340.510 1204.280 ;
        RECT 2341.350 1204.000 2351.550 1204.280 ;
        RECT 2352.390 1204.000 2362.590 1204.280 ;
        RECT 2363.430 1204.000 2373.630 1204.280 ;
        RECT 2374.470 1204.000 2384.670 1204.280 ;
        RECT 2385.510 1204.000 2395.710 1204.280 ;
        RECT 2396.550 1204.000 2406.750 1204.280 ;
        RECT 2407.590 1204.000 2417.790 1204.280 ;
        RECT 2418.630 1204.000 2428.830 1204.280 ;
        RECT 2429.670 1204.000 2439.410 1204.280 ;
        RECT 2440.250 1204.000 2450.450 1204.280 ;
        RECT 2451.290 1204.000 2461.490 1204.280 ;
        RECT 2462.330 1204.000 2472.530 1204.280 ;
        RECT 2473.370 1204.000 2483.570 1204.280 ;
        RECT 2484.410 1204.000 2494.610 1204.280 ;
        RECT 2495.450 1204.000 2505.650 1204.280 ;
        RECT 2506.490 1204.000 2516.690 1204.280 ;
        RECT 2517.530 1204.000 2527.730 1204.280 ;
        RECT 2528.570 1204.000 2538.770 1204.280 ;
        RECT 2539.610 1204.000 2549.810 1204.280 ;
        RECT 2550.650 1204.000 2560.850 1204.280 ;
        RECT 2561.690 1204.000 2571.890 1204.280 ;
        RECT 2572.730 1204.000 2582.930 1204.280 ;
        RECT 2583.770 1204.000 2593.970 1204.280 ;
        RECT 2594.810 1204.000 2594.990 1204.280 ;
      LAYER met2 ;
        RECT 1415.730 1200.610 1416.010 1204.000 ;
        RECT 1426.770 1200.610 1427.050 1204.000 ;
        RECT 1437.810 1200.610 1438.090 1204.000 ;
        RECT 1415.730 1200.470 1417.560 1200.610 ;
        RECT 1415.730 1200.000 1416.010 1200.470 ;
        RECT 1417.420 1191.010 1417.560 1200.470 ;
        RECT 1426.770 1200.470 1428.140 1200.610 ;
        RECT 1426.770 1200.000 1427.050 1200.470 ;
        RECT 1417.360 1190.690 1417.620 1191.010 ;
        RECT 1428.000 1190.330 1428.140 1200.470 ;
        RECT 1437.810 1200.470 1439.640 1200.610 ;
        RECT 1437.810 1200.000 1438.090 1200.470 ;
        RECT 1427.940 1190.010 1428.200 1190.330 ;
        RECT 1439.500 1187.270 1439.640 1200.470 ;
        RECT 1448.850 1200.000 1449.130 1204.000 ;
        RECT 1459.890 1200.610 1460.170 1204.000 ;
        RECT 1470.930 1200.610 1471.210 1204.000 ;
        RECT 1481.970 1200.610 1482.250 1204.000 ;
        RECT 1493.010 1200.610 1493.290 1204.000 ;
        RECT 1459.890 1200.470 1462.640 1200.610 ;
        RECT 1459.890 1200.000 1460.170 1200.470 ;
        RECT 1448.930 1199.250 1449.070 1200.000 ;
        RECT 1448.700 1199.110 1449.070 1199.250 ;
        RECT 1439.440 1186.950 1439.700 1187.270 ;
        RECT 1441.740 1186.950 1442.000 1187.270 ;
        RECT 1441.800 1019.845 1441.940 1186.950 ;
        RECT 1441.730 1019.475 1442.010 1019.845 ;
        RECT 1448.700 1019.165 1448.840 1199.110 ;
        RECT 1462.500 1051.950 1462.640 1200.470 ;
        RECT 1470.930 1200.470 1472.760 1200.610 ;
        RECT 1470.930 1200.000 1471.210 1200.470 ;
        RECT 1472.620 1192.370 1472.760 1200.470 ;
        RECT 1481.970 1200.470 1483.340 1200.610 ;
        RECT 1481.970 1200.000 1482.250 1200.470 ;
        RECT 1472.560 1192.050 1472.820 1192.370 ;
        RECT 1476.240 1192.050 1476.500 1192.370 ;
        RECT 1462.440 1051.630 1462.700 1051.950 ;
        RECT 1448.630 1018.795 1448.910 1019.165 ;
        RECT 1476.300 1014.550 1476.440 1192.050 ;
        RECT 1483.200 1014.890 1483.340 1200.470 ;
        RECT 1493.010 1200.470 1494.840 1200.610 ;
        RECT 1493.010 1200.000 1493.290 1200.470 ;
        RECT 1490.040 1190.690 1490.300 1191.010 ;
        RECT 1483.140 1014.570 1483.400 1014.890 ;
        RECT 1476.240 1014.230 1476.500 1014.550 ;
        RECT 1490.100 558.805 1490.240 1190.690 ;
        RECT 1494.700 1187.270 1494.840 1200.470 ;
        RECT 1504.050 1200.000 1504.330 1204.000 ;
        RECT 1515.090 1200.610 1515.370 1204.000 ;
        RECT 1526.130 1200.610 1526.410 1204.000 ;
        RECT 1537.170 1200.610 1537.450 1204.000 ;
        RECT 1548.210 1200.610 1548.490 1204.000 ;
        RECT 1515.090 1200.470 1516.920 1200.610 ;
        RECT 1515.090 1200.000 1515.370 1200.470 ;
        RECT 1504.130 1199.250 1504.270 1200.000 ;
        RECT 1503.900 1199.110 1504.270 1199.250 ;
        RECT 1494.640 1186.950 1494.900 1187.270 ;
        RECT 1496.940 1186.950 1497.200 1187.270 ;
        RECT 1496.480 1051.630 1496.740 1051.950 ;
        RECT 1496.540 1020.410 1496.680 1051.630 ;
        RECT 1497.000 1021.010 1497.140 1186.950 ;
        RECT 1496.940 1020.690 1497.200 1021.010 ;
        RECT 1496.930 1020.410 1497.210 1020.525 ;
        RECT 1496.540 1020.270 1497.210 1020.410 ;
        RECT 1503.900 1020.330 1504.040 1199.110 ;
        RECT 1516.780 1191.010 1516.920 1200.470 ;
        RECT 1526.130 1200.470 1527.960 1200.610 ;
        RECT 1526.130 1200.000 1526.410 1200.470 ;
        RECT 1527.820 1191.350 1527.960 1200.470 ;
        RECT 1537.170 1200.470 1538.540 1200.610 ;
        RECT 1537.170 1200.000 1537.450 1200.470 ;
        RECT 1527.760 1191.030 1528.020 1191.350 ;
        RECT 1516.720 1190.690 1516.980 1191.010 ;
        RECT 1538.400 1190.670 1538.540 1200.470 ;
        RECT 1548.210 1200.470 1550.040 1200.610 ;
        RECT 1548.210 1200.000 1548.490 1200.470 ;
        RECT 1549.900 1191.690 1550.040 1200.470 ;
        RECT 1559.250 1200.000 1559.530 1204.000 ;
        RECT 1570.290 1200.610 1570.570 1204.000 ;
        RECT 1580.870 1200.610 1581.150 1204.000 ;
        RECT 1591.910 1200.610 1592.190 1204.000 ;
        RECT 1602.950 1200.610 1603.230 1204.000 ;
        RECT 1570.290 1200.470 1573.040 1200.610 ;
        RECT 1570.290 1200.000 1570.570 1200.470 ;
        RECT 1559.330 1199.250 1559.470 1200.000 ;
        RECT 1559.100 1199.110 1559.470 1199.250 ;
        RECT 1559.100 1192.030 1559.240 1199.110 ;
        RECT 1559.040 1191.710 1559.300 1192.030 ;
        RECT 1549.840 1191.370 1550.100 1191.690 ;
        RECT 1538.340 1190.350 1538.600 1190.670 ;
        RECT 1496.930 1020.155 1497.210 1020.270 ;
        RECT 1503.840 1020.010 1504.100 1020.330 ;
        RECT 1572.900 1019.990 1573.040 1200.470 ;
        RECT 1580.870 1200.470 1582.700 1200.610 ;
        RECT 1580.870 1200.000 1581.150 1200.470 ;
        RECT 1582.560 1192.710 1582.700 1200.470 ;
        RECT 1591.910 1200.470 1593.740 1200.610 ;
        RECT 1591.910 1200.000 1592.190 1200.470 ;
        RECT 1582.500 1192.390 1582.760 1192.710 ;
        RECT 1586.640 1192.390 1586.900 1192.710 ;
        RECT 1572.840 1019.670 1573.100 1019.990 ;
        RECT 1586.700 1019.650 1586.840 1192.390 ;
        RECT 1586.640 1019.330 1586.900 1019.650 ;
        RECT 1593.600 1019.310 1593.740 1200.470 ;
        RECT 1602.950 1200.470 1604.780 1200.610 ;
        RECT 1602.950 1200.000 1603.230 1200.470 ;
        RECT 1604.640 1187.270 1604.780 1200.470 ;
        RECT 1613.990 1200.000 1614.270 1204.000 ;
        RECT 1625.030 1200.610 1625.310 1204.000 ;
        RECT 1636.070 1200.610 1636.350 1204.000 ;
        RECT 1647.110 1200.610 1647.390 1204.000 ;
        RECT 1658.150 1200.610 1658.430 1204.000 ;
        RECT 1625.030 1200.470 1628.240 1200.610 ;
        RECT 1625.030 1200.000 1625.310 1200.470 ;
        RECT 1614.070 1199.250 1614.210 1200.000 ;
        RECT 1614.070 1199.110 1614.440 1199.250 ;
        RECT 1604.580 1186.950 1604.840 1187.270 ;
        RECT 1607.340 1186.950 1607.600 1187.270 ;
        RECT 1593.540 1018.990 1593.800 1019.310 ;
        RECT 1607.400 1018.970 1607.540 1186.950 ;
        RECT 1607.340 1018.650 1607.600 1018.970 ;
        RECT 1614.300 1018.630 1614.440 1199.110 ;
        RECT 1614.240 1018.310 1614.500 1018.630 ;
        RECT 1628.100 1018.290 1628.240 1200.470 ;
        RECT 1636.070 1200.470 1637.900 1200.610 ;
        RECT 1636.070 1200.000 1636.350 1200.470 ;
        RECT 1637.760 1187.270 1637.900 1200.470 ;
        RECT 1647.110 1200.470 1648.940 1200.610 ;
        RECT 1647.110 1200.000 1647.390 1200.470 ;
        RECT 1641.380 1192.050 1641.640 1192.370 ;
        RECT 1637.700 1186.950 1637.960 1187.270 ;
        RECT 1628.040 1017.970 1628.300 1018.290 ;
        RECT 1641.440 1016.445 1641.580 1192.050 ;
        RECT 1648.800 1187.270 1648.940 1200.470 ;
        RECT 1658.150 1200.470 1659.980 1200.610 ;
        RECT 1658.150 1200.000 1658.430 1200.470 ;
        RECT 1655.640 1192.730 1655.900 1193.050 ;
        RECT 1641.840 1186.950 1642.100 1187.270 ;
        RECT 1648.740 1186.950 1649.000 1187.270 ;
        RECT 1641.900 1021.010 1642.040 1186.950 ;
        RECT 1648.740 1159.070 1649.000 1159.390 ;
        RECT 1648.800 1124.450 1648.940 1159.070 ;
        RECT 1647.420 1124.310 1648.940 1124.450 ;
        RECT 1647.420 1076.850 1647.560 1124.310 ;
        RECT 1646.960 1076.710 1647.560 1076.850 ;
        RECT 1646.960 1062.685 1647.100 1076.710 ;
        RECT 1646.890 1062.315 1647.170 1062.685 ;
        RECT 1641.840 1020.690 1642.100 1021.010 ;
        RECT 1641.840 1017.290 1642.100 1017.610 ;
        RECT 1641.900 1017.125 1642.040 1017.290 ;
        RECT 1654.720 1017.125 1654.980 1017.270 ;
        RECT 1641.830 1016.755 1642.110 1017.125 ;
        RECT 1654.710 1016.755 1654.990 1017.125 ;
        RECT 1655.700 1016.445 1655.840 1192.730 ;
        RECT 1659.840 1188.630 1659.980 1200.470 ;
        RECT 1669.190 1200.000 1669.470 1204.000 ;
        RECT 1680.230 1200.610 1680.510 1204.000 ;
        RECT 1691.270 1200.610 1691.550 1204.000 ;
        RECT 1702.310 1200.610 1702.590 1204.000 ;
        RECT 1713.350 1200.610 1713.630 1204.000 ;
        RECT 1724.390 1200.610 1724.670 1204.000 ;
        RECT 1735.430 1200.610 1735.710 1204.000 ;
        RECT 1746.470 1200.610 1746.750 1204.000 ;
        RECT 1757.050 1200.610 1757.330 1204.000 ;
        RECT 1768.090 1200.610 1768.370 1204.000 ;
        RECT 1680.230 1200.470 1683.440 1200.610 ;
        RECT 1680.230 1200.000 1680.510 1200.470 ;
        RECT 1669.270 1199.250 1669.410 1200.000 ;
        RECT 1669.270 1199.110 1669.640 1199.250 ;
        RECT 1668.520 1193.410 1668.780 1193.730 ;
        RECT 1662.540 1193.070 1662.800 1193.390 ;
        RECT 1659.780 1188.310 1660.040 1188.630 ;
        RECT 1641.370 1016.075 1641.650 1016.445 ;
        RECT 1655.630 1016.075 1655.910 1016.445 ;
        RECT 1662.080 1016.270 1662.340 1016.590 ;
        RECT 1662.600 1016.445 1662.740 1193.070 ;
        RECT 1667.600 1192.390 1667.860 1192.710 ;
        RECT 1667.660 1159.390 1667.800 1192.390 ;
        RECT 1668.580 1187.270 1668.720 1193.410 ;
        RECT 1669.500 1187.950 1669.640 1199.110 ;
        RECT 1675.880 1188.990 1676.140 1189.310 ;
        RECT 1669.440 1187.630 1669.700 1187.950 ;
        RECT 1668.520 1186.950 1668.780 1187.270 ;
        RECT 1669.440 1186.950 1669.700 1187.270 ;
        RECT 1667.600 1159.070 1667.860 1159.390 ;
        RECT 1669.500 1016.445 1669.640 1186.950 ;
        RECT 1675.940 1017.125 1676.080 1188.990 ;
        RECT 1676.340 1187.970 1676.600 1188.290 ;
        RECT 1675.420 1016.610 1675.680 1016.930 ;
        RECT 1675.870 1016.755 1676.150 1017.125 ;
        RECT 1662.140 1015.765 1662.280 1016.270 ;
        RECT 1662.530 1016.075 1662.810 1016.445 ;
        RECT 1668.980 1015.930 1669.240 1016.250 ;
        RECT 1669.430 1016.075 1669.710 1016.445 ;
        RECT 1669.040 1015.765 1669.180 1015.930 ;
        RECT 1675.480 1015.765 1675.620 1016.610 ;
        RECT 1676.400 1016.445 1676.540 1187.970 ;
        RECT 1683.300 1187.010 1683.440 1200.470 ;
        RECT 1690.660 1200.470 1691.550 1200.610 ;
        RECT 1686.920 1187.290 1687.180 1187.610 ;
        RECT 1683.300 1186.870 1683.900 1187.010 ;
        RECT 1684.160 1186.950 1684.420 1187.270 ;
        RECT 1682.320 1159.070 1682.580 1159.390 ;
        RECT 1682.380 1128.530 1682.520 1159.070 ;
        RECT 1682.380 1128.390 1682.980 1128.530 ;
        RECT 1682.840 1104.310 1682.980 1128.390 ;
        RECT 1682.780 1103.990 1683.040 1104.310 ;
        RECT 1683.240 1103.990 1683.500 1104.310 ;
        RECT 1683.300 1077.110 1683.440 1103.990 ;
        RECT 1683.240 1076.790 1683.500 1077.110 ;
        RECT 1683.240 1076.110 1683.500 1076.430 ;
        RECT 1683.300 1038.885 1683.440 1076.110 ;
        RECT 1683.230 1038.515 1683.510 1038.885 ;
        RECT 1680.020 1018.990 1680.280 1019.310 ;
        RECT 1680.080 1017.950 1680.220 1018.990 ;
        RECT 1680.020 1017.630 1680.280 1017.950 ;
        RECT 1683.760 1017.125 1683.900 1186.870 ;
        RECT 1684.220 1159.390 1684.360 1186.950 ;
        RECT 1684.160 1159.070 1684.420 1159.390 ;
        RECT 1686.980 1021.350 1687.120 1187.290 ;
        RECT 1690.660 1187.270 1690.800 1200.470 ;
        RECT 1691.270 1200.000 1691.550 1200.470 ;
        RECT 1700.780 1200.470 1702.590 1200.610 ;
        RECT 1697.960 1188.310 1698.220 1188.630 ;
        RECT 1691.060 1187.630 1691.320 1187.950 ;
        RECT 1690.600 1186.950 1690.860 1187.270 ;
        RECT 1686.920 1021.030 1687.180 1021.350 ;
        RECT 1689.680 1017.290 1689.940 1017.610 ;
        RECT 1683.690 1016.755 1683.970 1017.125 ;
        RECT 1676.330 1016.075 1676.610 1016.445 ;
        RECT 1683.240 1015.765 1683.500 1015.910 ;
        RECT 1648.740 1015.250 1649.000 1015.570 ;
        RECT 1662.070 1015.395 1662.350 1015.765 ;
        RECT 1668.970 1015.395 1669.250 1015.765 ;
        RECT 1675.410 1015.395 1675.690 1015.765 ;
        RECT 1683.230 1015.395 1683.510 1015.765 ;
        RECT 1648.800 1015.085 1648.940 1015.250 ;
        RECT 1683.240 1015.085 1683.500 1015.230 ;
        RECT 1689.740 1015.085 1689.880 1017.290 ;
        RECT 1691.120 1016.445 1691.260 1187.630 ;
        RECT 1698.020 1016.445 1698.160 1188.310 ;
        RECT 1700.780 1188.290 1700.920 1200.470 ;
        RECT 1702.310 1200.000 1702.590 1200.470 ;
        RECT 1711.820 1200.470 1713.630 1200.610 ;
        RECT 1707.620 1190.690 1707.880 1191.010 ;
        RECT 1700.720 1187.970 1700.980 1188.290 ;
        RECT 1704.400 1021.205 1704.660 1021.350 ;
        RECT 1704.390 1020.835 1704.670 1021.205 ;
        RECT 1706.240 1021.030 1706.500 1021.350 ;
        RECT 1706.300 1017.610 1706.440 1021.030 ;
        RECT 1707.680 1018.290 1707.820 1190.690 ;
        RECT 1711.820 1189.310 1711.960 1200.470 ;
        RECT 1713.350 1200.000 1713.630 1200.470 ;
        RECT 1722.860 1200.470 1724.670 1200.610 ;
        RECT 1722.860 1193.730 1723.000 1200.470 ;
        RECT 1724.390 1200.000 1724.670 1200.470 ;
        RECT 1733.900 1200.470 1735.710 1200.610 ;
        RECT 1722.800 1193.410 1723.060 1193.730 ;
        RECT 1733.900 1193.390 1734.040 1200.470 ;
        RECT 1735.430 1200.000 1735.710 1200.470 ;
        RECT 1745.860 1200.470 1746.750 1200.610 ;
        RECT 1733.840 1193.070 1734.100 1193.390 ;
        RECT 1745.860 1193.050 1746.000 1200.470 ;
        RECT 1746.470 1200.000 1746.750 1200.470 ;
        RECT 1755.520 1200.470 1757.330 1200.610 ;
        RECT 1745.800 1192.730 1746.060 1193.050 ;
        RECT 1755.520 1192.710 1755.660 1200.470 ;
        RECT 1757.050 1200.000 1757.330 1200.470 ;
        RECT 1766.560 1200.470 1768.370 1200.610 ;
        RECT 1755.460 1192.390 1755.720 1192.710 ;
        RECT 1766.560 1192.370 1766.700 1200.470 ;
        RECT 1768.090 1200.000 1768.370 1200.470 ;
        RECT 1779.130 1200.610 1779.410 1204.000 ;
        RECT 1790.170 1200.610 1790.450 1204.000 ;
        RECT 1801.210 1200.610 1801.490 1204.000 ;
        RECT 1812.250 1200.610 1812.530 1204.000 ;
        RECT 1823.290 1200.610 1823.570 1204.000 ;
        RECT 1779.130 1200.470 1780.040 1200.610 ;
        RECT 1779.130 1200.000 1779.410 1200.470 ;
        RECT 1766.500 1192.050 1766.760 1192.370 ;
        RECT 1714.520 1191.710 1714.780 1192.030 ;
        RECT 1711.760 1188.990 1712.020 1189.310 ;
        RECT 1711.300 1020.690 1711.560 1021.010 ;
        RECT 1711.360 1018.485 1711.500 1020.690 ;
        RECT 1707.620 1017.970 1707.880 1018.290 ;
        RECT 1711.290 1018.115 1711.570 1018.485 ;
        RECT 1711.300 1017.805 1711.560 1017.950 ;
        RECT 1706.240 1017.290 1706.500 1017.610 ;
        RECT 1711.290 1017.435 1711.570 1017.805 ;
        RECT 1712.280 1017.610 1713.800 1017.690 ;
        RECT 1712.220 1017.550 1713.860 1017.610 ;
        RECT 1712.220 1017.290 1712.480 1017.550 ;
        RECT 1713.600 1017.290 1713.860 1017.550 ;
        RECT 1700.720 1016.950 1700.980 1017.270 ;
        RECT 1691.050 1016.075 1691.330 1016.445 ;
        RECT 1697.950 1016.075 1698.230 1016.445 ;
        RECT 1696.120 1015.250 1696.380 1015.570 ;
        RECT 1696.180 1015.085 1696.320 1015.250 ;
        RECT 1700.780 1015.085 1700.920 1016.950 ;
        RECT 1714.580 1016.590 1714.720 1191.710 ;
        RECT 1721.420 1191.370 1721.680 1191.690 ;
        RECT 1714.980 1191.030 1715.240 1191.350 ;
        RECT 1715.040 1019.310 1715.180 1191.030 ;
        RECT 1717.280 1020.690 1717.540 1021.010 ;
        RECT 1714.980 1018.990 1715.240 1019.310 ;
        RECT 1707.160 1016.270 1707.420 1016.590 ;
        RECT 1714.520 1016.270 1714.780 1016.590 ;
        RECT 1707.220 1015.085 1707.360 1016.270 ;
        RECT 1713.600 1015.930 1713.860 1016.250 ;
        RECT 1713.660 1015.085 1713.800 1015.930 ;
        RECT 1717.340 1015.570 1717.480 1020.690 ;
        RECT 1718.200 1018.485 1718.460 1018.630 ;
        RECT 1718.190 1018.115 1718.470 1018.485 ;
        RECT 1718.200 1016.950 1718.460 1017.270 ;
        RECT 1717.740 1015.930 1718.000 1016.250 ;
        RECT 1717.800 1015.570 1717.940 1015.930 ;
        RECT 1717.280 1015.250 1717.540 1015.570 ;
        RECT 1717.740 1015.250 1718.000 1015.570 ;
        RECT 1718.260 1015.085 1718.400 1016.950 ;
        RECT 1721.480 1016.250 1721.620 1191.370 ;
        RECT 1735.220 1190.350 1735.480 1190.670 ;
        RECT 1728.320 1190.010 1728.580 1190.330 ;
        RECT 1728.380 1018.970 1728.520 1190.010 ;
        RECT 1735.280 1021.350 1735.420 1190.350 ;
        RECT 1732.000 1021.030 1732.260 1021.350 ;
        RECT 1735.220 1021.030 1735.480 1021.350 ;
        RECT 1725.100 1018.650 1725.360 1018.970 ;
        RECT 1728.320 1018.650 1728.580 1018.970 ;
        RECT 1725.160 1016.445 1725.300 1018.650 ;
        RECT 1732.060 1018.290 1732.200 1021.030 ;
        RECT 1741.660 1020.690 1741.920 1021.010 ;
        RECT 1748.100 1020.690 1748.360 1021.010 ;
        RECT 1752.230 1020.835 1752.510 1021.205 ;
        RECT 1759.600 1021.030 1759.860 1021.350 ;
        RECT 1752.240 1020.690 1752.500 1020.835 ;
        RECT 1738.900 1019.330 1739.160 1019.650 ;
        RECT 1732.000 1017.970 1732.260 1018.290 ;
        RECT 1735.680 1017.970 1735.940 1018.290 ;
        RECT 1732.000 1017.290 1732.260 1017.610 ;
        RECT 1732.060 1016.445 1732.200 1017.290 ;
        RECT 1721.420 1015.930 1721.680 1016.250 ;
        RECT 1725.090 1016.075 1725.370 1016.445 ;
        RECT 1731.990 1016.075 1732.270 1016.445 ;
        RECT 1729.700 1015.590 1729.960 1015.910 ;
        RECT 1724.640 1015.085 1724.900 1015.230 ;
        RECT 1729.760 1015.085 1729.900 1015.590 ;
        RECT 1735.740 1015.085 1735.880 1017.970 ;
        RECT 1738.960 1015.765 1739.100 1019.330 ;
        RECT 1738.890 1015.395 1739.170 1015.765 ;
        RECT 1741.720 1015.085 1741.860 1020.690 ;
        RECT 1745.800 1019.670 1746.060 1019.990 ;
        RECT 1745.860 1018.485 1746.000 1019.670 ;
        RECT 1745.790 1018.115 1746.070 1018.485 ;
        RECT 1748.160 1017.950 1748.300 1020.690 ;
        RECT 1759.140 1019.670 1759.400 1019.990 ;
        RECT 1748.100 1017.630 1748.360 1017.950 ;
        RECT 1748.100 1016.950 1748.360 1017.270 ;
        RECT 1745.800 1016.445 1746.060 1016.590 ;
        RECT 1745.790 1016.075 1746.070 1016.445 ;
        RECT 1748.160 1015.085 1748.300 1016.950 ;
        RECT 1755.460 1015.930 1755.720 1016.250 ;
        RECT 1755.920 1015.930 1756.180 1016.250 ;
        RECT 1755.520 1015.765 1755.660 1015.930 ;
        RECT 1755.450 1015.395 1755.730 1015.765 ;
        RECT 1755.980 1015.085 1756.120 1015.930 ;
        RECT 1759.200 1015.570 1759.340 1019.670 ;
        RECT 1759.660 1018.485 1759.800 1021.030 ;
        RECT 1776.610 1019.475 1776.890 1019.845 ;
        RECT 1766.500 1018.990 1766.760 1019.310 ;
        RECT 1772.940 1018.990 1773.200 1019.310 ;
        RECT 1759.590 1018.115 1759.870 1018.485 ;
        RECT 1766.040 1017.970 1766.300 1018.290 ;
        RECT 1766.100 1016.930 1766.240 1017.970 ;
        RECT 1766.040 1016.610 1766.300 1016.930 ;
        RECT 1759.140 1015.250 1759.400 1015.570 ;
        RECT 1759.200 1015.085 1759.340 1015.250 ;
        RECT 1766.100 1015.085 1766.240 1016.610 ;
        RECT 1766.560 1015.765 1766.700 1018.990 ;
        RECT 1766.490 1015.395 1766.770 1015.765 ;
        RECT 1773.000 1015.230 1773.140 1018.990 ;
        RECT 1773.400 1018.485 1773.660 1018.630 ;
        RECT 1773.390 1018.115 1773.670 1018.485 ;
        RECT 1776.680 1017.125 1776.820 1019.475 ;
        RECT 1778.000 1017.970 1778.260 1018.290 ;
        RECT 1776.610 1016.755 1776.890 1017.125 ;
        RECT 1778.060 1015.910 1778.200 1017.970 ;
        RECT 1779.900 1017.805 1780.040 1200.470 ;
        RECT 1790.170 1200.470 1793.840 1200.610 ;
        RECT 1790.170 1200.000 1790.450 1200.470 ;
        RECT 1786.730 1020.835 1787.010 1021.205 ;
        RECT 1786.740 1020.690 1787.000 1020.835 ;
        RECT 1787.660 1020.690 1787.920 1021.010 ;
        RECT 1787.200 1020.350 1787.460 1020.670 ;
        RECT 1780.300 1020.010 1780.560 1020.330 ;
        RECT 1779.830 1017.435 1780.110 1017.805 ;
        RECT 1780.360 1016.445 1780.500 1020.010 ;
        RECT 1787.260 1019.845 1787.400 1020.350 ;
        RECT 1787.190 1019.475 1787.470 1019.845 ;
        RECT 1787.720 1017.950 1787.860 1020.690 ;
        RECT 1790.420 1020.350 1790.680 1020.670 ;
        RECT 1787.660 1017.630 1787.920 1017.950 ;
        RECT 1782.140 1017.290 1782.400 1017.610 ;
        RECT 1780.290 1016.075 1780.570 1016.445 ;
        RECT 1778.000 1015.590 1778.260 1015.910 ;
        RECT 1772.940 1015.085 1773.200 1015.230 ;
        RECT 1778.060 1015.085 1778.200 1015.590 ;
        RECT 1782.200 1015.085 1782.340 1017.290 ;
        RECT 1787.720 1015.765 1787.860 1017.630 ;
        RECT 1790.480 1017.270 1790.620 1020.350 ;
        RECT 1793.700 1018.485 1793.840 1200.470 ;
        RECT 1801.210 1200.470 1803.040 1200.610 ;
        RECT 1801.210 1200.000 1801.490 1200.470 ;
        RECT 1802.900 1190.670 1803.040 1200.470 ;
        RECT 1812.250 1200.470 1814.540 1200.610 ;
        RECT 1812.250 1200.000 1812.530 1200.470 ;
        RECT 1802.840 1190.350 1803.100 1190.670 ;
        RECT 1800.080 1020.010 1800.340 1020.330 ;
        RECT 1793.630 1018.115 1793.910 1018.485 ;
        RECT 1790.420 1016.950 1790.680 1017.270 ;
        RECT 1787.650 1015.395 1787.930 1015.765 ;
        RECT 1790.480 1015.085 1790.620 1016.950 ;
        RECT 1800.140 1016.250 1800.280 1020.010 ;
        RECT 1806.060 1019.670 1806.320 1019.990 ;
        RECT 1800.080 1015.930 1800.340 1016.250 ;
        RECT 1800.140 1015.085 1800.280 1015.930 ;
        RECT 1806.120 1015.085 1806.260 1019.670 ;
        RECT 1807.900 1019.330 1808.160 1019.650 ;
        RECT 1812.960 1019.330 1813.220 1019.650 ;
        RECT 1807.960 1018.630 1808.100 1019.330 ;
        RECT 1807.900 1018.310 1808.160 1018.630 ;
        RECT 1813.020 1015.085 1813.160 1019.330 ;
        RECT 1814.400 1019.165 1814.540 1200.470 ;
        RECT 1823.290 1200.470 1825.120 1200.610 ;
        RECT 1823.290 1200.000 1823.570 1200.470 ;
        RECT 1824.980 1187.270 1825.120 1200.470 ;
        RECT 1834.330 1200.000 1834.610 1204.000 ;
        RECT 1845.370 1200.610 1845.650 1204.000 ;
        RECT 1843.840 1200.470 1845.650 1200.610 ;
        RECT 1834.410 1199.250 1834.550 1200.000 ;
        RECT 1834.410 1199.110 1834.780 1199.250 ;
        RECT 1834.120 1187.290 1834.380 1187.610 ;
        RECT 1824.920 1186.950 1825.180 1187.270 ;
        RECT 1831.820 1186.950 1832.080 1187.270 ;
        RECT 1831.880 1021.350 1832.020 1186.950 ;
        RECT 1831.820 1021.030 1832.080 1021.350 ;
        RECT 1834.180 1021.205 1834.320 1187.290 ;
        RECT 1834.110 1020.835 1834.390 1021.205 ;
        RECT 1834.640 1020.525 1834.780 1199.110 ;
        RECT 1843.840 1187.610 1843.980 1200.470 ;
        RECT 1845.370 1200.000 1845.650 1200.470 ;
        RECT 1856.410 1200.000 1856.690 1204.000 ;
        RECT 1867.450 1200.610 1867.730 1204.000 ;
        RECT 1878.490 1200.610 1878.770 1204.000 ;
        RECT 1889.530 1200.610 1889.810 1204.000 ;
        RECT 1900.570 1200.610 1900.850 1204.000 ;
        RECT 1911.610 1200.610 1911.890 1204.000 ;
        RECT 1922.190 1200.610 1922.470 1204.000 ;
        RECT 1933.230 1200.610 1933.510 1204.000 ;
        RECT 1944.270 1200.610 1944.550 1204.000 ;
        RECT 1955.310 1200.610 1955.590 1204.000 ;
        RECT 1966.350 1201.290 1966.630 1204.000 ;
        RECT 1965.740 1201.150 1966.630 1201.290 ;
        RECT 1867.450 1200.470 1869.280 1200.610 ;
        RECT 1867.450 1200.000 1867.730 1200.470 ;
        RECT 1856.490 1199.250 1856.630 1200.000 ;
        RECT 1856.260 1199.110 1856.630 1199.250 ;
        RECT 1855.740 1191.370 1856.000 1191.690 ;
        RECT 1843.780 1187.290 1844.040 1187.610 ;
        RECT 1835.040 1186.950 1835.300 1187.270 ;
        RECT 1821.700 1020.010 1821.960 1020.330 ;
        RECT 1834.570 1020.155 1834.850 1020.525 ;
        RECT 1821.760 1019.730 1821.900 1020.010 ;
        RECT 1835.100 1019.845 1835.240 1186.950 ;
        RECT 1842.400 1021.205 1842.660 1021.350 ;
        RECT 1855.800 1021.205 1855.940 1191.370 ;
        RECT 1856.260 1187.270 1856.400 1199.110 ;
        RECT 1869.140 1190.330 1869.280 1200.470 ;
        RECT 1878.490 1200.470 1880.320 1200.610 ;
        RECT 1878.490 1200.000 1878.770 1200.470 ;
        RECT 1869.080 1190.010 1869.340 1190.330 ;
        RECT 1880.180 1188.630 1880.320 1200.470 ;
        RECT 1889.530 1200.470 1890.440 1200.610 ;
        RECT 1889.530 1200.000 1889.810 1200.470 ;
        RECT 1880.120 1188.310 1880.380 1188.630 ;
        RECT 1884.260 1188.310 1884.520 1188.630 ;
        RECT 1856.200 1186.950 1856.460 1187.270 ;
        RECT 1842.390 1020.835 1842.670 1021.205 ;
        RECT 1855.730 1020.835 1856.010 1021.205 ;
        RECT 1869.540 1020.010 1869.800 1020.330 ;
        RECT 1821.760 1019.590 1822.360 1019.730 ;
        RECT 1814.330 1018.795 1814.610 1019.165 ;
        RECT 1817.560 1018.990 1817.820 1019.310 ;
        RECT 1817.620 1015.085 1817.760 1018.990 ;
        RECT 1821.700 1018.650 1821.960 1018.970 ;
        RECT 1821.760 1017.125 1821.900 1018.650 ;
        RECT 1822.220 1017.950 1822.360 1019.590 ;
        RECT 1835.030 1019.475 1835.310 1019.845 ;
        RECT 1824.000 1018.650 1824.260 1018.970 ;
        RECT 1822.160 1017.630 1822.420 1017.950 ;
        RECT 1821.690 1016.755 1821.970 1017.125 ;
        RECT 1824.060 1015.085 1824.200 1018.650 ;
        RECT 1869.600 1017.950 1869.740 1020.010 ;
        RECT 1869.540 1017.630 1869.800 1017.950 ;
        RECT 1648.730 1014.715 1649.010 1015.085 ;
        RECT 1683.230 1014.715 1683.510 1015.085 ;
        RECT 1689.670 1014.715 1689.950 1015.085 ;
        RECT 1696.110 1014.715 1696.390 1015.085 ;
        RECT 1700.710 1014.715 1700.990 1015.085 ;
        RECT 1707.150 1014.715 1707.430 1015.085 ;
        RECT 1713.590 1014.715 1713.870 1015.085 ;
        RECT 1718.190 1014.715 1718.470 1015.085 ;
        RECT 1724.630 1014.715 1724.910 1015.085 ;
        RECT 1729.690 1014.715 1729.970 1015.085 ;
        RECT 1735.670 1014.715 1735.950 1015.085 ;
        RECT 1741.650 1014.715 1741.930 1015.085 ;
        RECT 1748.090 1014.715 1748.370 1015.085 ;
        RECT 1755.910 1014.715 1756.190 1015.085 ;
        RECT 1759.130 1014.715 1759.410 1015.085 ;
        RECT 1766.030 1014.715 1766.310 1015.085 ;
        RECT 1772.930 1014.715 1773.210 1015.085 ;
        RECT 1777.990 1014.715 1778.270 1015.085 ;
        RECT 1782.130 1014.715 1782.410 1015.085 ;
        RECT 1787.190 1014.715 1787.470 1015.085 ;
        RECT 1790.410 1014.715 1790.690 1015.085 ;
        RECT 1794.090 1014.715 1794.370 1015.085 ;
        RECT 1800.070 1014.715 1800.350 1015.085 ;
        RECT 1806.050 1014.715 1806.330 1015.085 ;
        RECT 1812.950 1014.715 1813.230 1015.085 ;
        RECT 1817.550 1014.715 1817.830 1015.085 ;
        RECT 1823.990 1014.715 1824.270 1015.085 ;
        RECT 1787.200 1014.570 1787.460 1014.715 ;
        RECT 1794.160 1014.550 1794.300 1014.715 ;
        RECT 1794.100 1014.230 1794.360 1014.550 ;
        RECT 1490.030 558.435 1490.310 558.805 ;
        RECT 1503.830 556.395 1504.110 556.765 ;
        RECT 1503.900 554.870 1504.040 556.395 ;
      LAYER met2 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
      LAYER met2 ;
        RECT 1884.320 908.325 1884.460 1188.310 ;
        RECT 1890.300 1024.750 1890.440 1200.470 ;
        RECT 1900.570 1200.470 1904.240 1200.610 ;
        RECT 1900.570 1200.000 1900.850 1200.470 ;
        RECT 1902.200 1192.390 1902.460 1192.710 ;
        RECT 1901.740 1192.050 1902.000 1192.370 ;
        RECT 1901.280 1191.710 1901.540 1192.030 ;
        RECT 1900.820 1190.690 1901.080 1191.010 ;
        RECT 1890.240 1024.430 1890.500 1024.750 ;
        RECT 1898.980 917.330 1899.240 917.650 ;
        RECT 1899.040 913.765 1899.180 917.330 ;
        RECT 1898.970 913.395 1899.250 913.765 ;
        RECT 1884.250 907.955 1884.530 908.325 ;
        RECT 1899.900 620.510 1900.160 620.830 ;
        RECT 1899.960 615.925 1900.100 620.510 ;
        RECT 1899.890 615.555 1900.170 615.925 ;
        RECT 1900.360 592.970 1900.620 593.290 ;
        RECT 1900.420 590.765 1900.560 592.970 ;
        RECT 1900.350 590.395 1900.630 590.765 ;
        RECT 1900.360 579.370 1900.620 579.690 ;
        RECT 1900.420 579.205 1900.560 579.370 ;
        RECT 1900.350 578.835 1900.630 579.205 ;
        RECT 1900.880 573.765 1901.020 1190.690 ;
        RECT 1901.340 593.485 1901.480 1191.710 ;
        RECT 1901.800 601.645 1901.940 1192.050 ;
        RECT 1902.260 610.485 1902.400 1192.390 ;
        RECT 1904.100 1006.050 1904.240 1200.470 ;
        RECT 1911.610 1200.470 1913.440 1200.610 ;
        RECT 1911.610 1200.000 1911.890 1200.470 ;
        RECT 1913.300 1187.270 1913.440 1200.470 ;
        RECT 1922.190 1200.470 1924.940 1200.610 ;
        RECT 1922.190 1200.000 1922.470 1200.470 ;
        RECT 1913.240 1186.950 1913.500 1187.270 ;
        RECT 1917.840 1186.950 1918.100 1187.270 ;
        RECT 1917.900 1006.390 1918.040 1186.950 ;
        RECT 1918.300 1021.030 1918.560 1021.350 ;
        RECT 1918.360 1020.330 1918.500 1021.030 ;
        RECT 1918.300 1020.010 1918.560 1020.330 ;
        RECT 1924.800 1006.730 1924.940 1200.470 ;
        RECT 1933.230 1200.470 1935.060 1200.610 ;
        RECT 1933.230 1200.000 1933.510 1200.470 ;
        RECT 1934.920 1187.270 1935.060 1200.470 ;
        RECT 1944.270 1200.470 1945.640 1200.610 ;
        RECT 1944.270 1200.000 1944.550 1200.470 ;
        RECT 1934.860 1186.950 1935.120 1187.270 ;
        RECT 1938.540 1186.950 1938.800 1187.270 ;
        RECT 1938.600 1007.070 1938.740 1186.950 ;
        RECT 1945.500 1007.410 1945.640 1200.470 ;
        RECT 1955.310 1200.470 1957.140 1200.610 ;
        RECT 1955.310 1200.000 1955.590 1200.470 ;
        RECT 1957.000 1187.270 1957.140 1200.470 ;
        RECT 1965.740 1191.350 1965.880 1201.150 ;
        RECT 1966.350 1200.000 1966.630 1201.150 ;
        RECT 1977.390 1200.610 1977.670 1204.000 ;
        RECT 1988.430 1200.610 1988.710 1204.000 ;
        RECT 1999.470 1200.610 1999.750 1204.000 ;
        RECT 2010.510 1200.610 2010.790 1204.000 ;
        RECT 2021.550 1200.610 2021.830 1204.000 ;
        RECT 2032.590 1200.610 2032.870 1204.000 ;
        RECT 2043.630 1200.610 2043.910 1204.000 ;
        RECT 2054.670 1200.610 2054.950 1204.000 ;
        RECT 1975.860 1200.470 1977.670 1200.610 ;
        RECT 1969.820 1192.730 1970.080 1193.050 ;
        RECT 1965.680 1191.030 1965.940 1191.350 ;
        RECT 1956.940 1186.950 1957.200 1187.270 ;
        RECT 1959.240 1186.950 1959.500 1187.270 ;
        RECT 1945.440 1007.090 1945.700 1007.410 ;
        RECT 1938.540 1006.750 1938.800 1007.070 ;
        RECT 1924.740 1006.410 1925.000 1006.730 ;
        RECT 1917.840 1006.070 1918.100 1006.390 ;
        RECT 1904.040 1005.730 1904.300 1006.050 ;
        RECT 1959.300 1003.670 1959.440 1186.950 ;
        RECT 1966.140 1021.030 1966.400 1021.350 ;
        RECT 1966.200 1020.330 1966.340 1021.030 ;
        RECT 1966.140 1020.010 1966.400 1020.330 ;
        RECT 1959.240 1003.350 1959.500 1003.670 ;
        RECT 1902.190 610.115 1902.470 610.485 ;
        RECT 1901.730 601.275 1902.010 601.645 ;
        RECT 1901.270 593.115 1901.550 593.485 ;
        RECT 1969.880 593.290 1970.020 1192.730 ;
        RECT 1975.860 1191.690 1976.000 1200.470 ;
        RECT 1977.390 1200.000 1977.670 1200.470 ;
        RECT 1987.360 1200.470 1988.710 1200.610 ;
        RECT 1975.800 1191.370 1976.060 1191.690 ;
        RECT 1987.360 1187.270 1987.500 1200.470 ;
        RECT 1988.430 1200.000 1988.710 1200.470 ;
        RECT 1997.940 1200.470 1999.750 1200.610 ;
        RECT 1997.940 1192.710 1998.080 1200.470 ;
        RECT 1999.470 1200.000 1999.750 1200.470 ;
        RECT 2008.980 1200.470 2010.790 1200.610 ;
        RECT 1997.880 1192.390 1998.140 1192.710 ;
        RECT 2008.980 1192.370 2009.120 1200.470 ;
        RECT 2010.510 1200.000 2010.790 1200.470 ;
        RECT 2020.020 1200.470 2021.830 1200.610 ;
        RECT 2008.920 1192.050 2009.180 1192.370 ;
        RECT 2020.020 1192.030 2020.160 1200.470 ;
        RECT 2021.550 1200.000 2021.830 1200.470 ;
        RECT 2031.060 1200.470 2032.870 1200.610 ;
        RECT 2031.060 1193.050 2031.200 1200.470 ;
        RECT 2032.590 1200.000 2032.870 1200.470 ;
        RECT 2042.560 1200.470 2043.910 1200.610 ;
        RECT 2031.000 1192.730 2031.260 1193.050 ;
        RECT 2019.960 1191.710 2020.220 1192.030 ;
        RECT 2042.560 1191.690 2042.700 1200.470 ;
        RECT 2043.630 1200.000 2043.910 1200.470 ;
        RECT 2053.140 1200.470 2054.950 1200.610 ;
        RECT 1997.420 1191.370 1997.680 1191.690 ;
        RECT 2042.500 1191.370 2042.760 1191.690 ;
        RECT 1976.720 1186.950 1976.980 1187.270 ;
        RECT 1987.300 1186.950 1987.560 1187.270 ;
        RECT 1976.780 620.830 1976.920 1186.950 ;
        RECT 1976.720 620.510 1976.980 620.830 ;
        RECT 1969.820 592.970 1970.080 593.290 ;
        RECT 1997.480 579.690 1997.620 1191.370 ;
        RECT 2053.140 1191.010 2053.280 1200.470 ;
        RECT 2054.670 1200.000 2054.950 1200.470 ;
        RECT 2065.710 1200.610 2065.990 1204.000 ;
        RECT 2065.710 1200.470 2067.540 1200.610 ;
        RECT 2065.710 1200.000 2065.990 1200.470 ;
        RECT 2067.400 1192.030 2067.540 1200.470 ;
        RECT 2076.750 1200.000 2077.030 1204.000 ;
        RECT 2087.790 1200.610 2088.070 1204.000 ;
        RECT 2098.370 1200.610 2098.650 1204.000 ;
        RECT 2109.410 1200.610 2109.690 1204.000 ;
        RECT 2120.450 1200.610 2120.730 1204.000 ;
        RECT 2087.790 1200.470 2089.620 1200.610 ;
        RECT 2087.790 1200.000 2088.070 1200.470 ;
        RECT 2076.830 1199.250 2076.970 1200.000 ;
        RECT 2076.600 1199.110 2076.970 1199.250 ;
        RECT 2076.600 1192.370 2076.740 1199.110 ;
        RECT 2076.540 1192.050 2076.800 1192.370 ;
        RECT 2067.340 1191.710 2067.600 1192.030 ;
        RECT 2089.480 1191.690 2089.620 1200.470 ;
        RECT 2098.370 1200.470 2100.200 1200.610 ;
        RECT 2098.370 1200.000 2098.650 1200.470 ;
        RECT 2100.060 1192.710 2100.200 1200.470 ;
        RECT 2109.410 1200.470 2111.240 1200.610 ;
        RECT 2109.410 1200.000 2109.690 1200.470 ;
        RECT 2111.100 1193.050 2111.240 1200.470 ;
        RECT 2120.450 1200.470 2122.280 1200.610 ;
        RECT 2120.450 1200.000 2120.730 1200.470 ;
        RECT 2122.140 1193.390 2122.280 1200.470 ;
        RECT 2131.490 1200.000 2131.770 1204.000 ;
        RECT 2142.530 1200.610 2142.810 1204.000 ;
        RECT 2153.570 1200.610 2153.850 1204.000 ;
        RECT 2164.610 1200.610 2164.890 1204.000 ;
        RECT 2175.650 1200.610 2175.930 1204.000 ;
        RECT 2186.690 1200.610 2186.970 1204.000 ;
        RECT 2197.730 1200.610 2198.010 1204.000 ;
        RECT 2208.770 1200.610 2209.050 1204.000 ;
        RECT 2219.810 1200.610 2220.090 1204.000 ;
        RECT 2230.850 1200.610 2231.130 1204.000 ;
        RECT 2142.530 1200.470 2144.360 1200.610 ;
        RECT 2142.530 1200.000 2142.810 1200.470 ;
        RECT 2131.570 1199.250 2131.710 1200.000 ;
        RECT 2131.570 1199.110 2131.940 1199.250 ;
        RECT 2131.800 1193.730 2131.940 1199.110 ;
        RECT 2131.740 1193.410 2132.000 1193.730 ;
        RECT 2122.080 1193.070 2122.340 1193.390 ;
        RECT 2111.040 1192.730 2111.300 1193.050 ;
        RECT 2100.000 1192.390 2100.260 1192.710 ;
        RECT 2089.420 1191.370 2089.680 1191.690 ;
        RECT 2144.220 1191.010 2144.360 1200.470 ;
        RECT 2152.960 1200.470 2153.850 1200.610 ;
        RECT 2053.080 1190.690 2053.340 1191.010 ;
        RECT 2144.160 1190.690 2144.420 1191.010 ;
        RECT 2014.900 1021.030 2015.160 1021.350 ;
        RECT 2062.740 1021.030 2063.000 1021.350 ;
        RECT 2111.500 1021.030 2111.760 1021.350 ;
        RECT 2014.960 1020.330 2015.100 1021.030 ;
        RECT 2062.800 1020.330 2062.940 1021.030 ;
        RECT 2111.560 1020.330 2111.700 1021.030 ;
        RECT 2014.900 1020.010 2015.160 1020.330 ;
        RECT 2062.740 1020.010 2063.000 1020.330 ;
        RECT 2111.500 1020.010 2111.760 1020.330 ;
        RECT 2152.960 1018.970 2153.100 1200.470 ;
        RECT 2153.570 1200.000 2153.850 1200.470 ;
        RECT 2159.860 1200.470 2164.890 1200.610 ;
        RECT 2159.340 1021.030 2159.600 1021.350 ;
        RECT 2159.400 1020.330 2159.540 1021.030 ;
        RECT 2159.340 1020.010 2159.600 1020.330 ;
        RECT 2159.860 1019.310 2160.000 1200.470 ;
        RECT 2164.610 1200.000 2164.890 1200.470 ;
        RECT 2173.660 1200.470 2175.930 1200.610 ;
        RECT 2173.660 1019.650 2173.800 1200.470 ;
        RECT 2175.650 1200.000 2175.930 1200.470 ;
        RECT 2180.560 1200.470 2186.970 1200.610 ;
        RECT 2180.560 1019.990 2180.700 1200.470 ;
        RECT 2186.690 1200.000 2186.970 1200.470 ;
        RECT 2194.360 1200.470 2198.010 1200.610 ;
        RECT 2194.360 1020.330 2194.500 1200.470 ;
        RECT 2197.730 1200.000 2198.010 1200.470 ;
        RECT 2208.160 1200.470 2209.050 1200.610 ;
        RECT 2208.160 1020.670 2208.300 1200.470 ;
        RECT 2208.770 1200.000 2209.050 1200.470 ;
        RECT 2215.060 1200.470 2220.090 1200.610 ;
        RECT 2215.060 1021.010 2215.200 1200.470 ;
        RECT 2219.810 1200.000 2220.090 1200.470 ;
        RECT 2228.860 1200.470 2231.130 1200.610 ;
        RECT 2215.000 1020.690 2215.260 1021.010 ;
        RECT 2208.100 1020.350 2208.360 1020.670 ;
        RECT 2194.300 1020.010 2194.560 1020.330 ;
        RECT 2180.500 1019.670 2180.760 1019.990 ;
        RECT 2173.600 1019.330 2173.860 1019.650 ;
        RECT 2159.800 1018.990 2160.060 1019.310 ;
        RECT 2152.900 1018.650 2153.160 1018.970 ;
        RECT 2228.860 1017.610 2229.000 1200.470 ;
        RECT 2230.850 1200.000 2231.130 1200.470 ;
        RECT 2241.890 1200.000 2242.170 1204.000 ;
        RECT 2252.930 1200.610 2253.210 1204.000 ;
        RECT 2263.510 1200.610 2263.790 1204.000 ;
        RECT 2274.550 1200.610 2274.830 1204.000 ;
        RECT 2285.590 1200.610 2285.870 1204.000 ;
        RECT 2296.630 1200.610 2296.910 1204.000 ;
        RECT 2307.670 1200.610 2307.950 1204.000 ;
        RECT 2318.710 1200.610 2318.990 1204.000 ;
        RECT 2329.750 1200.610 2330.030 1204.000 ;
        RECT 2340.790 1200.610 2341.070 1204.000 ;
        RECT 2252.930 1200.470 2256.140 1200.610 ;
        RECT 2252.930 1200.000 2253.210 1200.470 ;
        RECT 2241.970 1199.250 2242.110 1200.000 ;
        RECT 2241.740 1199.110 2242.110 1199.250 ;
        RECT 2238.920 1190.690 2239.180 1191.010 ;
        RECT 2238.980 1019.650 2239.120 1190.690 ;
        RECT 2241.740 1025.090 2241.880 1199.110 ;
        RECT 2245.820 1193.410 2246.080 1193.730 ;
        RECT 2242.140 1190.690 2242.400 1191.010 ;
        RECT 2241.680 1024.770 2241.940 1025.090 ;
        RECT 2242.200 1021.205 2242.340 1190.690 ;
        RECT 2242.130 1020.835 2242.410 1021.205 ;
        RECT 2245.880 1020.670 2246.020 1193.410 ;
        RECT 2252.720 1193.070 2252.980 1193.390 ;
        RECT 2252.780 1021.350 2252.920 1193.070 ;
        RECT 2256.000 1025.430 2256.140 1200.470 ;
        RECT 2263.510 1200.470 2265.340 1200.610 ;
        RECT 2263.510 1200.000 2263.790 1200.470 ;
        RECT 2259.620 1192.730 2259.880 1193.050 ;
        RECT 2255.940 1025.110 2256.200 1025.430 ;
        RECT 2252.720 1021.030 2252.980 1021.350 ;
        RECT 2254.560 1021.030 2254.820 1021.350 ;
        RECT 2259.680 1021.205 2259.820 1192.730 ;
        RECT 2265.200 1192.710 2265.340 1200.470 ;
        RECT 2274.550 1200.470 2276.380 1200.610 ;
        RECT 2274.550 1200.000 2274.830 1200.470 ;
        RECT 2276.240 1193.390 2276.380 1200.470 ;
        RECT 2285.590 1200.470 2287.420 1200.610 ;
        RECT 2285.590 1200.000 2285.870 1200.470 ;
        RECT 2276.180 1193.070 2276.440 1193.390 ;
        RECT 2287.280 1193.050 2287.420 1200.470 ;
        RECT 2296.630 1200.470 2297.540 1200.610 ;
        RECT 2296.630 1200.000 2296.910 1200.470 ;
        RECT 2287.220 1192.730 2287.480 1193.050 ;
        RECT 2290.440 1192.730 2290.700 1193.050 ;
        RECT 2265.140 1192.390 2265.400 1192.710 ;
        RECT 2266.520 1192.050 2266.780 1192.370 ;
        RECT 2260.540 1191.710 2260.800 1192.030 ;
        RECT 2260.600 1191.350 2260.740 1191.710 ;
        RECT 2260.080 1191.030 2260.340 1191.350 ;
        RECT 2260.540 1191.030 2260.800 1191.350 ;
        RECT 2260.140 1189.990 2260.280 1191.030 ;
        RECT 2260.080 1189.670 2260.340 1189.990 ;
        RECT 2266.580 1021.205 2266.720 1192.050 ;
        RECT 2280.320 1191.710 2280.580 1192.030 ;
        RECT 2283.540 1191.710 2283.800 1192.030 ;
        RECT 2273.420 1191.370 2273.680 1191.690 ;
        RECT 2276.640 1191.370 2276.900 1191.690 ;
        RECT 2245.820 1020.525 2246.080 1020.670 ;
        RECT 2254.620 1020.525 2254.760 1021.030 ;
        RECT 2259.610 1020.835 2259.890 1021.205 ;
        RECT 2266.510 1020.835 2266.790 1021.205 ;
        RECT 2245.810 1020.155 2246.090 1020.525 ;
        RECT 2254.550 1020.155 2254.830 1020.525 ;
        RECT 2238.920 1019.330 2239.180 1019.650 ;
        RECT 2242.140 1019.330 2242.400 1019.650 ;
        RECT 2228.800 1017.290 2229.060 1017.610 ;
        RECT 2242.200 1006.925 2242.340 1019.330 ;
        RECT 2259.680 1018.290 2259.820 1020.835 ;
        RECT 2266.520 1020.690 2266.780 1020.835 ;
        RECT 2266.580 1020.535 2266.720 1020.690 ;
        RECT 2269.740 1020.010 2270.000 1020.330 ;
        RECT 2259.620 1017.970 2259.880 1018.290 ;
        RECT 2269.800 1017.125 2269.940 1020.010 ;
        RECT 2273.480 1019.845 2273.620 1191.370 ;
        RECT 2276.700 1021.205 2276.840 1191.370 ;
        RECT 2276.630 1020.835 2276.910 1021.205 ;
        RECT 2276.640 1019.845 2276.900 1019.990 ;
        RECT 2273.410 1019.475 2273.690 1019.845 ;
        RECT 2276.630 1019.475 2276.910 1019.845 ;
        RECT 2273.480 1017.950 2273.620 1019.475 ;
        RECT 2273.420 1017.630 2273.680 1017.950 ;
        RECT 2280.380 1017.125 2280.520 1191.710 ;
        RECT 2281.240 1191.030 2281.500 1191.350 ;
        RECT 2281.300 1020.525 2281.440 1191.030 ;
        RECT 2283.600 1021.205 2283.740 1191.710 ;
        RECT 2287.220 1189.670 2287.480 1189.990 ;
        RECT 2287.280 1172.730 2287.420 1189.670 ;
        RECT 2287.280 1172.590 2287.880 1172.730 ;
        RECT 2287.740 1125.130 2287.880 1172.590 ;
        RECT 2287.740 1124.990 2288.340 1125.130 ;
        RECT 2288.200 1028.490 2288.340 1124.990 ;
        RECT 2287.220 1028.170 2287.480 1028.490 ;
        RECT 2288.140 1028.170 2288.400 1028.490 ;
        RECT 2283.530 1020.835 2283.810 1021.205 ;
        RECT 2281.230 1020.155 2281.510 1020.525 ;
        RECT 2287.280 1020.410 2287.420 1028.170 ;
        RECT 2287.280 1020.270 2287.880 1020.410 ;
        RECT 2269.730 1016.755 2270.010 1017.125 ;
        RECT 2280.310 1016.755 2280.590 1017.125 ;
        RECT 2281.300 1016.590 2281.440 1020.155 ;
        RECT 2287.220 1019.330 2287.480 1019.650 ;
        RECT 2283.540 1017.290 2283.800 1017.610 ;
        RECT 2283.600 1017.125 2283.740 1017.290 ;
        RECT 2283.530 1016.755 2283.810 1017.125 ;
        RECT 2281.240 1016.270 2281.500 1016.590 ;
        RECT 2287.280 1016.445 2287.420 1019.330 ;
        RECT 2287.210 1016.075 2287.490 1016.445 ;
        RECT 2287.220 1015.930 2287.480 1016.075 ;
        RECT 2287.280 1015.775 2287.420 1015.930 ;
        RECT 2255.020 1015.250 2255.280 1015.570 ;
        RECT 2249.040 1015.085 2249.300 1015.230 ;
        RECT 2255.080 1015.085 2255.220 1015.250 ;
        RECT 2249.030 1014.715 2249.310 1015.085 ;
        RECT 2255.010 1014.715 2255.290 1015.085 ;
        RECT 2262.830 1014.715 2263.110 1015.085 ;
        RECT 2262.900 1014.550 2263.040 1014.715 ;
        RECT 2262.840 1014.230 2263.100 1014.550 ;
        RECT 2242.130 1006.555 2242.410 1006.925 ;
        RECT 2287.740 1003.330 2287.880 1020.270 ;
        RECT 2289.980 1019.330 2290.240 1019.650 ;
        RECT 2290.040 1015.085 2290.180 1019.330 ;
        RECT 2290.500 1019.310 2290.640 1192.730 ;
        RECT 2296.880 1191.030 2297.140 1191.350 ;
        RECT 2293.660 1020.350 2293.920 1020.670 ;
        RECT 2290.440 1018.990 2290.700 1019.310 ;
        RECT 2293.720 1016.930 2293.860 1020.350 ;
        RECT 2293.660 1016.610 2293.920 1016.930 ;
        RECT 2293.720 1015.085 2293.860 1016.610 ;
        RECT 2296.940 1016.445 2297.080 1191.030 ;
        RECT 2297.400 1018.970 2297.540 1200.470 ;
        RECT 2307.670 1200.470 2309.500 1200.610 ;
        RECT 2307.670 1200.000 2307.950 1200.470 ;
        RECT 2309.360 1188.970 2309.500 1200.470 ;
        RECT 2318.710 1200.470 2320.540 1200.610 ;
        RECT 2318.710 1200.000 2318.990 1200.470 ;
        RECT 2317.580 1192.390 2317.840 1192.710 ;
        RECT 2311.140 1192.050 2311.400 1192.370 ;
        RECT 2309.300 1188.650 2309.560 1188.970 ;
        RECT 2303.320 1021.030 2303.580 1021.350 ;
        RECT 2297.340 1018.650 2297.600 1018.970 ;
        RECT 2303.380 1017.270 2303.520 1021.030 ;
        RECT 2304.240 1018.310 2304.500 1018.630 ;
        RECT 2303.320 1016.950 2303.580 1017.270 ;
        RECT 2304.300 1017.125 2304.440 1018.310 ;
        RECT 2307.920 1017.970 2308.180 1018.290 ;
        RECT 2296.870 1016.075 2297.150 1016.445 ;
        RECT 2303.380 1015.085 2303.520 1016.950 ;
        RECT 2304.230 1016.755 2304.510 1017.125 ;
        RECT 2307.980 1015.085 2308.120 1017.970 ;
        RECT 2311.200 1016.445 2311.340 1192.050 ;
        RECT 2312.060 1020.690 2312.320 1021.010 ;
        RECT 2311.130 1016.075 2311.410 1016.445 ;
        RECT 2312.120 1015.910 2312.260 1020.690 ;
        RECT 2317.120 1017.630 2317.380 1017.950 ;
        RECT 2312.060 1015.590 2312.320 1015.910 ;
        RECT 2312.120 1015.085 2312.260 1015.590 ;
        RECT 2317.180 1015.085 2317.320 1017.630 ;
        RECT 2317.640 1017.125 2317.780 1192.390 ;
        RECT 2320.400 1187.270 2320.540 1200.470 ;
        RECT 2329.750 1200.470 2331.580 1200.610 ;
        RECT 2329.750 1200.000 2330.030 1200.470 ;
        RECT 2324.480 1189.670 2324.740 1189.990 ;
        RECT 2320.340 1186.950 2320.600 1187.270 ;
        RECT 2318.040 1020.690 2318.300 1021.010 ;
        RECT 2317.570 1016.755 2317.850 1017.125 ;
        RECT 2318.100 1016.445 2318.240 1020.690 ;
        RECT 2323.560 1017.290 2323.820 1017.610 ;
        RECT 2318.030 1016.075 2318.310 1016.445 ;
        RECT 2323.620 1015.085 2323.760 1017.290 ;
        RECT 2324.540 1016.445 2324.680 1189.670 ;
        RECT 2331.440 1187.610 2331.580 1200.470 ;
        RECT 2340.790 1200.470 2342.620 1200.610 ;
        RECT 2340.790 1200.000 2341.070 1200.470 ;
        RECT 2338.740 1188.990 2339.000 1189.310 ;
        RECT 2331.380 1187.290 2331.640 1187.610 ;
        RECT 2324.940 1186.950 2325.200 1187.270 ;
        RECT 2325.000 1021.350 2325.140 1186.950 ;
        RECT 2330.920 1025.790 2331.180 1026.110 ;
        RECT 2324.940 1021.030 2325.200 1021.350 ;
        RECT 2330.980 1021.205 2331.120 1025.790 ;
        RECT 2338.800 1021.205 2338.940 1188.990 ;
        RECT 2342.480 1187.270 2342.620 1200.470 ;
        RECT 2351.830 1200.000 2352.110 1204.000 ;
        RECT 2362.870 1200.610 2363.150 1204.000 ;
        RECT 2359.960 1200.470 2363.150 1200.610 ;
        RECT 2351.910 1199.250 2352.050 1200.000 ;
        RECT 2351.910 1199.110 2352.280 1199.250 ;
        RECT 2351.620 1188.310 2351.880 1188.630 ;
        RECT 2342.420 1186.950 2342.680 1187.270 ;
        RECT 2345.640 1186.950 2345.900 1187.270 ;
        RECT 2345.180 1025.450 2345.440 1025.770 ;
        RECT 2345.240 1021.205 2345.380 1025.450 ;
        RECT 2330.910 1020.835 2331.190 1021.205 ;
        RECT 2338.730 1020.835 2339.010 1021.205 ;
        RECT 2345.170 1020.835 2345.450 1021.205 ;
        RECT 2342.420 1016.610 2342.680 1016.930 ;
        RECT 2324.470 1016.075 2324.750 1016.445 ;
        RECT 2329.540 1016.270 2329.800 1016.590 ;
        RECT 2329.600 1015.085 2329.740 1016.270 ;
        RECT 2335.520 1015.930 2335.780 1016.250 ;
        RECT 2335.580 1015.085 2335.720 1015.930 ;
        RECT 2342.480 1015.085 2342.620 1016.610 ;
        RECT 2289.970 1014.715 2290.250 1015.085 ;
        RECT 2293.650 1014.715 2293.930 1015.085 ;
        RECT 2303.310 1014.715 2303.590 1015.085 ;
        RECT 2307.910 1014.715 2308.190 1015.085 ;
        RECT 2312.050 1014.715 2312.330 1015.085 ;
        RECT 2317.110 1014.715 2317.390 1015.085 ;
        RECT 2323.550 1014.715 2323.830 1015.085 ;
        RECT 2329.530 1014.715 2329.810 1015.085 ;
        RECT 2335.510 1014.715 2335.790 1015.085 ;
        RECT 2342.410 1014.715 2342.690 1015.085 ;
        RECT 2345.700 1014.890 2345.840 1186.950 ;
        RECT 2351.680 1020.525 2351.820 1188.310 ;
        RECT 2352.140 1028.150 2352.280 1199.110 ;
        RECT 2359.960 1187.010 2360.100 1200.470 ;
        RECT 2362.870 1200.000 2363.150 1200.470 ;
        RECT 2373.910 1200.000 2374.190 1204.000 ;
        RECT 2384.950 1200.610 2385.230 1204.000 ;
        RECT 2395.990 1200.610 2396.270 1204.000 ;
        RECT 2407.030 1200.610 2407.310 1204.000 ;
        RECT 2418.070 1200.610 2418.350 1204.000 ;
        RECT 2383.420 1200.470 2385.230 1200.610 ;
        RECT 2373.990 1199.250 2374.130 1200.000 ;
        RECT 2373.760 1199.110 2374.130 1199.250 ;
        RECT 2363.120 1193.410 2363.380 1193.730 ;
        RECT 2359.500 1186.870 2360.100 1187.010 ;
        RECT 2352.080 1027.830 2352.340 1028.150 ;
        RECT 2352.540 1026.130 2352.800 1026.450 ;
        RECT 2352.600 1021.205 2352.740 1026.130 ;
        RECT 2359.500 1021.205 2359.640 1186.870 ;
        RECT 2359.900 1027.830 2360.160 1028.150 ;
        RECT 2352.530 1020.835 2352.810 1021.205 ;
        RECT 2359.430 1020.835 2359.710 1021.205 ;
        RECT 2351.610 1020.155 2351.890 1020.525 ;
        RECT 2353.920 1020.350 2354.180 1020.670 ;
        RECT 2359.960 1020.525 2360.100 1027.830 ;
        RECT 2353.980 1017.950 2354.120 1020.350 ;
        RECT 2359.890 1020.155 2360.170 1020.525 ;
        RECT 2363.180 1018.630 2363.320 1193.410 ;
        RECT 2370.020 1190.350 2370.280 1190.670 ;
        RECT 2364.040 1189.330 2364.300 1189.650 ;
        RECT 2363.580 1187.290 2363.840 1187.610 ;
        RECT 2363.640 1022.030 2363.780 1187.290 ;
        RECT 2363.580 1021.710 2363.840 1022.030 ;
        RECT 2364.100 1021.010 2364.240 1189.330 ;
        RECT 2364.500 1188.650 2364.760 1188.970 ;
        RECT 2364.040 1020.690 2364.300 1021.010 ;
        RECT 2364.560 1020.670 2364.700 1188.650 ;
        RECT 2363.580 1020.350 2363.840 1020.670 ;
        RECT 2364.500 1020.350 2364.760 1020.670 ;
        RECT 2363.120 1018.310 2363.380 1018.630 ;
        RECT 2355.760 1017.970 2356.020 1018.290 ;
        RECT 2353.920 1017.630 2354.180 1017.950 ;
        RECT 2347.020 1016.950 2347.280 1017.270 ;
        RECT 2347.080 1015.085 2347.220 1016.950 ;
        RECT 2355.290 1016.075 2355.570 1016.445 ;
        RECT 2355.360 1015.910 2355.500 1016.075 ;
        RECT 2355.820 1015.910 2355.960 1017.970 ;
        RECT 2358.060 1017.290 2358.320 1017.610 ;
        RECT 2358.120 1016.590 2358.260 1017.290 ;
        RECT 2363.640 1016.590 2363.780 1020.350 ;
        RECT 2370.080 1018.630 2370.220 1190.350 ;
        RECT 2373.760 1026.450 2373.900 1199.110 ;
        RECT 2383.420 1188.630 2383.560 1200.470 ;
        RECT 2384.950 1200.000 2385.230 1200.470 ;
        RECT 2394.460 1200.470 2396.270 1200.610 ;
        RECT 2383.820 1193.070 2384.080 1193.390 ;
        RECT 2383.360 1188.310 2383.620 1188.630 ;
        RECT 2373.700 1026.130 2373.960 1026.450 ;
        RECT 2383.880 1021.350 2384.020 1193.070 ;
        RECT 2384.280 1192.730 2384.540 1193.050 ;
        RECT 2373.700 1021.205 2373.960 1021.350 ;
        RECT 2373.690 1020.835 2373.970 1021.205 ;
        RECT 2383.820 1021.030 2384.080 1021.350 ;
        RECT 2384.340 1021.010 2384.480 1192.730 ;
        RECT 2394.460 1025.770 2394.600 1200.470 ;
        RECT 2395.990 1200.000 2396.270 1200.470 ;
        RECT 2405.500 1200.470 2407.310 1200.610 ;
        RECT 2405.500 1189.310 2405.640 1200.470 ;
        RECT 2407.030 1200.000 2407.310 1200.470 ;
        RECT 2415.160 1200.470 2418.350 1200.610 ;
        RECT 2405.440 1188.990 2405.700 1189.310 ;
        RECT 2415.160 1026.110 2415.300 1200.470 ;
        RECT 2418.070 1200.000 2418.350 1200.470 ;
        RECT 2429.110 1200.000 2429.390 1204.000 ;
        RECT 2439.690 1200.610 2439.970 1204.000 ;
        RECT 2450.730 1200.610 2451.010 1204.000 ;
        RECT 2461.770 1200.610 2462.050 1204.000 ;
        RECT 2472.810 1200.610 2473.090 1204.000 ;
        RECT 2483.850 1200.610 2484.130 1204.000 ;
        RECT 2494.890 1200.610 2495.170 1204.000 ;
        RECT 2505.930 1200.610 2506.210 1204.000 ;
        RECT 2516.970 1200.610 2517.250 1204.000 ;
        RECT 2528.010 1200.610 2528.290 1204.000 ;
        RECT 2539.050 1200.610 2539.330 1204.000 ;
        RECT 2550.090 1200.610 2550.370 1204.000 ;
        RECT 2561.130 1200.610 2561.410 1204.000 ;
        RECT 2572.170 1200.610 2572.450 1204.000 ;
        RECT 2583.210 1200.610 2583.490 1204.000 ;
        RECT 2594.250 1200.610 2594.530 1204.000 ;
        RECT 2438.160 1200.470 2439.970 1200.610 ;
        RECT 2429.190 1199.250 2429.330 1200.000 ;
        RECT 2428.960 1199.110 2429.330 1199.250 ;
        RECT 2428.960 1189.990 2429.100 1199.110 ;
        RECT 2428.900 1189.670 2429.160 1189.990 ;
        RECT 2438.160 1189.650 2438.300 1200.470 ;
        RECT 2439.690 1200.000 2439.970 1200.470 ;
        RECT 2449.660 1200.470 2451.010 1200.610 ;
        RECT 2449.660 1192.710 2449.800 1200.470 ;
        RECT 2450.730 1200.000 2451.010 1200.470 ;
        RECT 2460.240 1200.470 2462.050 1200.610 ;
        RECT 2449.600 1192.390 2449.860 1192.710 ;
        RECT 2460.240 1192.370 2460.380 1200.470 ;
        RECT 2461.770 1200.000 2462.050 1200.470 ;
        RECT 2471.280 1200.470 2473.090 1200.610 ;
        RECT 2471.280 1193.730 2471.420 1200.470 ;
        RECT 2472.810 1200.000 2473.090 1200.470 ;
        RECT 2482.320 1200.470 2484.130 1200.610 ;
        RECT 2471.220 1193.410 2471.480 1193.730 ;
        RECT 2460.180 1192.050 2460.440 1192.370 ;
        RECT 2482.320 1191.350 2482.460 1200.470 ;
        RECT 2483.850 1200.000 2484.130 1200.470 ;
        RECT 2491.060 1200.470 2495.170 1200.610 ;
        RECT 2482.260 1191.030 2482.520 1191.350 ;
        RECT 2481.800 1190.010 2482.060 1190.330 ;
        RECT 2438.100 1189.330 2438.360 1189.650 ;
        RECT 2415.100 1025.790 2415.360 1026.110 ;
        RECT 2394.400 1025.450 2394.660 1025.770 ;
        RECT 2415.100 1025.110 2415.360 1025.430 ;
        RECT 2403.140 1021.205 2403.400 1021.350 ;
        RECT 2380.600 1020.690 2380.860 1021.010 ;
        RECT 2384.280 1020.690 2384.540 1021.010 ;
        RECT 2403.130 1020.835 2403.410 1021.205 ;
        RECT 2408.200 1020.690 2408.460 1021.010 ;
        RECT 2380.660 1020.525 2380.800 1020.690 ;
        RECT 2387.500 1020.525 2387.760 1020.670 ;
        RECT 2380.590 1020.155 2380.870 1020.525 ;
        RECT 2387.490 1020.155 2387.770 1020.525 ;
        RECT 2394.400 1018.990 2394.660 1019.310 ;
        RECT 2388.420 1018.650 2388.680 1018.970 ;
        RECT 2370.020 1018.310 2370.280 1018.630 ;
        RECT 2373.240 1017.630 2373.500 1017.950 ;
        RECT 2373.700 1017.630 2373.960 1017.950 ;
        RECT 2358.060 1016.270 2358.320 1016.590 ;
        RECT 2363.580 1016.270 2363.840 1016.590 ;
        RECT 2355.300 1015.590 2355.560 1015.910 ;
        RECT 2355.760 1015.590 2356.020 1015.910 ;
        RECT 2355.820 1015.085 2355.960 1015.590 ;
        RECT 2363.640 1015.085 2363.780 1016.270 ;
        RECT 2373.300 1015.085 2373.440 1017.630 ;
        RECT 2373.760 1016.590 2373.900 1017.630 ;
        RECT 2377.840 1017.290 2378.100 1017.610 ;
        RECT 2373.700 1016.270 2373.960 1016.590 ;
        RECT 2377.900 1015.085 2378.040 1017.290 ;
        RECT 2387.960 1017.125 2388.220 1017.270 ;
        RECT 2387.500 1016.610 2387.760 1016.930 ;
        RECT 2387.950 1016.755 2388.230 1017.125 ;
        RECT 2380.600 1015.930 2380.860 1016.250 ;
        RECT 2381.050 1016.075 2381.330 1016.445 ;
        RECT 2381.060 1015.930 2381.320 1016.075 ;
        RECT 2380.660 1015.085 2380.800 1015.930 ;
        RECT 2387.560 1015.085 2387.700 1016.610 ;
        RECT 2388.480 1016.445 2388.620 1018.650 ;
        RECT 2394.460 1017.125 2394.600 1018.990 ;
        RECT 2408.260 1018.485 2408.400 1020.690 ;
        RECT 2408.190 1018.115 2408.470 1018.485 ;
        RECT 2408.200 1017.805 2408.460 1017.950 ;
        RECT 2408.190 1017.435 2408.470 1017.805 ;
        RECT 2415.160 1017.125 2415.300 1025.110 ;
        RECT 2422.000 1024.770 2422.260 1025.090 ;
        RECT 2422.060 1021.205 2422.200 1024.770 ;
        RECT 2450.980 1024.430 2451.240 1024.750 ;
        RECT 2421.990 1020.835 2422.270 1021.205 ;
        RECT 2451.040 1020.525 2451.180 1024.430 ;
        RECT 2450.970 1020.155 2451.250 1020.525 ;
        RECT 2428.900 1018.485 2429.160 1018.630 ;
        RECT 2428.890 1018.115 2429.170 1018.485 ;
        RECT 2422.000 1017.290 2422.260 1017.610 ;
        RECT 2422.060 1017.125 2422.200 1017.290 ;
        RECT 2394.390 1016.755 2394.670 1017.125 ;
        RECT 2415.090 1016.755 2415.370 1017.125 ;
        RECT 2421.990 1016.755 2422.270 1017.125 ;
        RECT 2388.410 1016.075 2388.690 1016.445 ;
        RECT 2394.400 1015.590 2394.660 1015.910 ;
        RECT 2402.220 1015.590 2402.480 1015.910 ;
        RECT 2394.460 1015.085 2394.600 1015.590 ;
        RECT 2402.280 1015.085 2402.420 1015.590 ;
        RECT 2345.640 1014.570 2345.900 1014.890 ;
        RECT 2347.010 1014.715 2347.290 1015.085 ;
        RECT 2355.750 1014.715 2356.030 1015.085 ;
        RECT 2363.570 1014.715 2363.850 1015.085 ;
        RECT 2366.790 1014.715 2367.070 1015.085 ;
        RECT 2373.230 1014.715 2373.510 1015.085 ;
        RECT 2377.830 1014.715 2378.110 1015.085 ;
        RECT 2380.590 1014.715 2380.870 1015.085 ;
        RECT 2387.490 1014.715 2387.770 1015.085 ;
        RECT 2394.390 1014.715 2394.670 1015.085 ;
        RECT 2402.210 1014.715 2402.490 1015.085 ;
        RECT 2415.090 1014.715 2415.370 1015.085 ;
        RECT 2366.800 1014.570 2367.060 1014.715 ;
        RECT 2373.240 1014.570 2373.500 1014.715 ;
        RECT 2415.100 1014.570 2415.360 1014.715 ;
        RECT 2287.680 1003.010 2287.940 1003.330 ;
        RECT 2094.020 1001.310 2094.280 1001.630 ;
        RECT 2094.080 917.650 2094.220 1001.310 ;
        RECT 2094.020 917.330 2094.280 917.650 ;
        RECT 1997.420 579.370 1997.680 579.690 ;
        RECT 1900.810 573.395 1901.090 573.765 ;
        RECT 2083.890 556.395 2084.170 556.765 ;
        RECT 2083.960 554.870 2084.100 556.395 ;
      LAYER met2 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met2 ;
        RECT 2481.860 906.850 2482.000 1190.010 ;
        RECT 2491.060 1019.650 2491.200 1200.470 ;
        RECT 2494.890 1200.000 2495.170 1200.470 ;
        RECT 2504.860 1200.470 2506.210 1200.610 ;
        RECT 2504.860 1192.030 2505.000 1200.470 ;
        RECT 2505.930 1200.000 2506.210 1200.470 ;
        RECT 2511.760 1200.470 2517.250 1200.610 ;
        RECT 2504.800 1191.710 2505.060 1192.030 ;
        RECT 2511.760 1019.990 2511.900 1200.470 ;
        RECT 2516.970 1200.000 2517.250 1200.470 ;
        RECT 2526.480 1200.470 2528.290 1200.610 ;
        RECT 2526.480 1191.690 2526.620 1200.470 ;
        RECT 2528.010 1200.000 2528.290 1200.470 ;
        RECT 2532.460 1200.470 2539.330 1200.610 ;
        RECT 2526.420 1191.370 2526.680 1191.690 ;
        RECT 2532.460 1020.330 2532.600 1200.470 ;
        RECT 2539.050 1200.000 2539.330 1200.470 ;
        RECT 2546.260 1200.470 2550.370 1200.610 ;
        RECT 2532.400 1020.010 2532.660 1020.330 ;
        RECT 2511.700 1019.670 2511.960 1019.990 ;
        RECT 2491.000 1019.330 2491.260 1019.650 ;
        RECT 2546.260 1014.550 2546.400 1200.470 ;
        RECT 2550.090 1200.000 2550.370 1200.470 ;
        RECT 2560.060 1200.470 2561.410 1200.610 ;
        RECT 2560.060 1015.570 2560.200 1200.470 ;
        RECT 2561.130 1200.000 2561.410 1200.470 ;
        RECT 2566.960 1200.470 2572.450 1200.610 ;
        RECT 2560.000 1015.250 2560.260 1015.570 ;
        RECT 2566.960 1015.230 2567.100 1200.470 ;
        RECT 2572.170 1200.000 2572.450 1200.470 ;
        RECT 2581.680 1200.470 2583.490 1200.610 ;
        RECT 2581.680 1191.010 2581.820 1200.470 ;
        RECT 2583.210 1200.000 2583.490 1200.470 ;
        RECT 2593.640 1200.470 2594.530 1200.610 ;
        RECT 2593.640 1197.130 2593.780 1200.470 ;
        RECT 2594.250 1200.000 2594.530 1200.470 ;
        RECT 2587.600 1196.810 2587.860 1197.130 ;
        RECT 2593.580 1196.810 2593.840 1197.130 ;
        RECT 2581.620 1190.690 2581.880 1191.010 ;
        RECT 2566.900 1014.910 2567.160 1015.230 ;
        RECT 2546.200 1014.230 2546.460 1014.550 ;
        RECT 2498.820 1007.090 2499.080 1007.410 ;
        RECT 2498.360 1003.350 2498.620 1003.670 ;
        RECT 2497.900 1003.010 2498.160 1003.330 ;
        RECT 2482.250 906.850 2482.530 906.965 ;
        RECT 2481.860 906.710 2482.530 906.850 ;
        RECT 2482.250 906.595 2482.530 906.710 ;
        RECT 2497.960 576.485 2498.100 1003.010 ;
        RECT 2498.420 579.205 2498.560 1003.350 ;
        RECT 2498.880 590.765 2499.020 1007.090 ;
        RECT 2499.280 1006.750 2499.540 1007.070 ;
        RECT 2499.340 593.485 2499.480 1006.750 ;
        RECT 2499.740 1006.410 2500.000 1006.730 ;
        RECT 2499.800 604.365 2499.940 1006.410 ;
        RECT 2500.200 1006.070 2500.460 1006.390 ;
        RECT 2500.260 610.485 2500.400 1006.070 ;
        RECT 2500.660 1005.730 2500.920 1006.050 ;
        RECT 2500.720 618.645 2500.860 1005.730 ;
        RECT 2587.660 1001.630 2587.800 1196.810 ;
        RECT 2587.600 1001.310 2587.860 1001.630 ;
        RECT 2587.660 917.650 2587.800 1001.310 ;
        RECT 2504.340 917.330 2504.600 917.650 ;
        RECT 2587.600 917.330 2587.860 917.650 ;
        RECT 2504.400 915.805 2504.540 917.330 ;
        RECT 2504.330 915.435 2504.610 915.805 ;
        RECT 2500.650 618.275 2500.930 618.645 ;
        RECT 2500.190 610.115 2500.470 610.485 ;
        RECT 2499.730 603.995 2500.010 604.365 ;
        RECT 2499.270 593.115 2499.550 593.485 ;
        RECT 2498.810 590.395 2499.090 590.765 ;
        RECT 2498.350 578.835 2498.630 579.205 ;
        RECT 2497.890 576.115 2498.170 576.485 ;
        RECT 1503.840 554.550 1504.100 554.870 ;
        RECT 2083.900 554.550 2084.160 554.870 ;
      LAYER via2 ;
        RECT 1868.150 3063.600 1868.430 3063.880 ;
        RECT 1490.030 3033.000 1490.310 3033.280 ;
        RECT 1489.570 3026.880 1489.850 3027.160 ;
        RECT 1489.110 3018.720 1489.390 3019.000 ;
        RECT 1488.650 3012.600 1488.930 3012.880 ;
        RECT 1488.190 3004.440 1488.470 3004.720 ;
        RECT 1487.730 2999.000 1488.010 2999.280 ;
        RECT 1487.270 2990.160 1487.550 2990.440 ;
        RECT 1486.810 2701.160 1487.090 2701.440 ;
        RECT 1486.350 2692.320 1486.630 2692.600 ;
        RECT 1417.350 2410.800 1417.630 2411.080 ;
        RECT 2442.690 3063.600 2442.970 3063.880 ;
        RECT 2469.830 3063.600 2470.110 3063.880 ;
        RECT 1898.510 3047.960 1898.790 3048.240 ;
        RECT 1899.890 3047.960 1900.170 3048.240 ;
        RECT 1898.050 2746.720 1898.330 2747.000 ;
        RECT 1898.050 2704.560 1898.330 2704.840 ;
        RECT 1490.030 2411.480 1490.310 2411.760 ;
        RECT 1569.610 2593.720 1569.890 2594.000 ;
        RECT 1573.750 2593.720 1574.030 2594.000 ;
        RECT 1586.630 2593.720 1586.910 2594.000 ;
        RECT 1591.230 2593.720 1591.510 2594.000 ;
        RECT 1598.590 2593.720 1598.870 2594.000 ;
        RECT 1604.110 2593.720 1604.390 2594.000 ;
        RECT 1614.690 2593.720 1614.970 2594.000 ;
        RECT 1621.590 2593.720 1621.870 2594.000 ;
        RECT 1626.650 2593.720 1626.930 2594.000 ;
        RECT 1651.030 2593.720 1651.310 2594.000 ;
        RECT 1565.470 2592.360 1565.750 2592.640 ;
        RECT 1573.290 2592.360 1573.570 2592.640 ;
        RECT 1581.110 2593.040 1581.390 2593.320 ;
        RECT 1587.090 2593.040 1587.370 2593.320 ;
        RECT 1608.250 2592.360 1608.530 2592.640 ;
        RECT 1639.070 2593.040 1639.350 2593.320 ;
        RECT 1644.590 2593.040 1644.870 2593.320 ;
        RECT 1661.610 2593.720 1661.890 2594.000 ;
        RECT 1669.890 2593.720 1670.170 2594.000 ;
        RECT 1690.590 2593.720 1690.870 2594.000 ;
        RECT 1697.950 2593.720 1698.230 2594.000 ;
        RECT 1656.090 2593.040 1656.370 2593.320 ;
        RECT 1607.790 2591.680 1608.070 2591.960 ;
        RECT 1586.170 2591.000 1586.450 2591.280 ;
        RECT 1566.390 2589.640 1566.670 2589.920 ;
        RECT 1552.130 2588.280 1552.410 2588.560 ;
        RECT 1538.330 2587.600 1538.610 2587.880 ;
        RECT 1545.230 2587.600 1545.510 2587.880 ;
        RECT 1551.210 2587.600 1551.490 2587.880 ;
        RECT 1559.490 2588.280 1559.770 2588.560 ;
        RECT 1559.030 2587.600 1559.310 2587.880 ;
        RECT 1621.590 2592.360 1621.870 2592.640 ;
        RECT 1633.550 2592.360 1633.830 2592.640 ;
        RECT 1614.690 2591.000 1614.970 2591.280 ;
        RECT 1593.990 2590.320 1594.270 2590.600 ;
        RECT 1587.090 2589.640 1587.370 2589.920 ;
        RECT 1600.890 2589.640 1601.170 2589.920 ;
        RECT 1593.990 2410.120 1594.270 2410.400 ;
        RECT 1609.630 2410.120 1609.910 2410.400 ;
        RECT 1621.590 2588.280 1621.870 2588.560 ;
        RECT 1667.130 2592.360 1667.410 2592.640 ;
        RECT 1679.550 2593.040 1679.830 2593.320 ;
        RECT 1685.530 2592.360 1685.810 2592.640 ;
        RECT 1738.430 2593.720 1738.710 2594.000 ;
        RECT 1707.610 2593.040 1707.890 2593.320 ;
        RECT 1732.910 2593.040 1733.190 2593.320 ;
        RECT 1702.550 2592.360 1702.830 2592.640 ;
        RECT 1656.090 2590.320 1656.370 2590.600 ;
        RECT 1678.630 2590.320 1678.910 2590.600 ;
        RECT 1642.290 2589.640 1642.570 2589.920 ;
        RECT 1631.250 2588.960 1631.530 2589.240 ;
        RECT 1635.390 2588.280 1635.670 2588.560 ;
        RECT 1649.190 2587.600 1649.470 2587.880 ;
        RECT 1662.990 2589.640 1663.270 2589.920 ;
        RECT 1743.950 2593.040 1744.230 2593.320 ;
        RECT 1725.550 2592.360 1725.830 2592.640 ;
        RECT 1713.130 2591.680 1713.410 2591.960 ;
        RECT 1718.190 2591.680 1718.470 2591.960 ;
        RECT 1683.690 2588.960 1683.970 2589.240 ;
        RECT 1690.590 2588.960 1690.870 2589.240 ;
        RECT 1662.990 2588.280 1663.270 2588.560 ;
        RECT 1669.890 2588.280 1670.170 2588.560 ;
        RECT 1697.490 2588.280 1697.770 2588.560 ;
        RECT 1697.030 2587.600 1697.310 2587.880 ;
        RECT 1745.330 2588.280 1745.610 2588.560 ;
        RECT 1703.930 2587.600 1704.210 2587.880 ;
        RECT 1714.510 2587.600 1714.790 2587.880 ;
        RECT 1721.410 2587.600 1721.690 2587.880 ;
        RECT 1731.530 2587.600 1731.810 2587.880 ;
        RECT 1736.590 2587.600 1736.870 2587.880 ;
        RECT 1744.870 2587.600 1745.150 2587.880 ;
        RECT 1835.950 2412.160 1836.230 2412.440 ;
        RECT 1877.350 2412.160 1877.630 2412.440 ;
        RECT 2087.110 3030.960 2087.390 3031.240 ;
        RECT 2083.890 2699.120 2084.170 2699.400 ;
        RECT 1898.510 2410.800 1898.790 2411.080 ;
        RECT 1942.670 2411.480 1942.950 2411.760 ;
        RECT 1932.550 2410.800 1932.830 2411.080 ;
        RECT 1945.890 2410.800 1946.170 2411.080 ;
        RECT 2087.570 3024.160 2087.850 3024.440 ;
        RECT 2088.030 3016.000 2088.310 3016.280 ;
        RECT 2088.490 3009.880 2088.770 3010.160 ;
        RECT 2088.950 3001.720 2089.230 3002.000 ;
        RECT 2089.410 2996.280 2089.690 2996.560 ;
        RECT 2089.870 2988.120 2090.150 2988.400 ;
        RECT 2090.330 2691.640 2090.610 2691.920 ;
        RECT 2482.250 3049.320 2482.530 3049.600 ;
        RECT 2497.890 2747.400 2498.170 2747.680 ;
        RECT 2497.890 2710.000 2498.170 2710.280 ;
        RECT 2497.890 2704.560 2498.170 2704.840 ;
        RECT 2126.670 2598.480 2126.950 2598.760 ;
        RECT 2215.910 2593.720 2216.190 2594.000 ;
        RECT 2256.390 2593.720 2256.670 2594.000 ;
        RECT 2262.830 2593.720 2263.110 2594.000 ;
        RECT 2268.350 2593.720 2268.630 2594.000 ;
        RECT 2297.790 2593.720 2298.070 2594.000 ;
        RECT 2305.150 2593.720 2305.430 2594.000 ;
        RECT 2146.450 2593.040 2146.730 2593.320 ;
        RECT 2145.990 2591.680 2146.270 2591.960 ;
        RECT 2152.890 2592.360 2153.170 2592.640 ;
        RECT 2132.190 2590.320 2132.470 2590.600 ;
        RECT 2176.810 2590.320 2177.090 2590.600 ;
        RECT 2179.570 2590.320 2179.850 2590.600 ;
        RECT 2183.710 2590.320 2183.990 2590.600 ;
        RECT 2090.330 2410.800 2090.610 2411.080 ;
        RECT 2170.370 2588.960 2170.650 2589.240 ;
        RECT 2163.010 2588.280 2163.290 2588.560 ;
        RECT 2166.230 2588.280 2166.510 2588.560 ;
        RECT 2173.130 2588.280 2173.410 2588.560 ;
        RECT 2168.990 2559.720 2169.270 2560.000 ;
        RECT 2169.910 2559.720 2170.190 2560.000 ;
        RECT 2168.070 2414.880 2168.350 2415.160 ;
        RECT 2168.990 2414.880 2169.270 2415.160 ;
        RECT 2180.030 2588.280 2180.310 2588.560 ;
        RECT 2186.470 2589.640 2186.750 2589.920 ;
        RECT 2186.930 2588.280 2187.210 2588.560 ;
        RECT 2193.830 2588.280 2194.110 2588.560 ;
        RECT 2190.610 2587.600 2190.890 2587.880 ;
        RECT 2193.370 2587.600 2193.650 2587.880 ;
        RECT 2197.510 2588.280 2197.790 2588.560 ;
        RECT 2204.410 2588.280 2204.690 2588.560 ;
        RECT 2200.730 2587.600 2201.010 2587.880 ;
        RECT 2207.630 2587.600 2207.910 2587.880 ;
        RECT 2209.470 2591.000 2209.750 2591.280 ;
        RECT 2214.530 2587.600 2214.810 2587.880 ;
        RECT 2220.510 2593.040 2220.790 2593.320 ;
        RECT 2235.690 2592.360 2235.970 2592.640 ;
        RECT 2227.870 2591.000 2228.150 2591.280 ;
        RECT 2228.330 2588.280 2228.610 2588.560 ;
        RECT 2221.430 2587.600 2221.710 2587.880 ;
        RECT 2227.870 2587.600 2228.150 2587.880 ;
        RECT 2232.930 2591.680 2233.210 2591.960 ;
        RECT 2249.490 2592.360 2249.770 2592.640 ;
        RECT 2243.970 2591.680 2244.250 2591.960 ;
        RECT 2291.810 2593.040 2292.090 2593.320 ;
        RECT 2297.790 2593.040 2298.070 2593.320 ;
        RECT 2311.590 2593.040 2311.870 2593.320 ;
        RECT 2332.290 2593.040 2332.570 2593.320 ;
        RECT 2280.310 2592.360 2280.590 2592.640 ;
        RECT 2285.370 2592.360 2285.650 2592.640 ;
        RECT 2276.170 2591.680 2276.450 2591.960 ;
        RECT 2339.190 2592.360 2339.470 2592.640 ;
        RECT 2318.490 2591.680 2318.770 2591.960 ;
        RECT 2332.290 2591.680 2332.570 2591.960 ;
        RECT 2325.390 2591.000 2325.670 2591.280 ;
        RECT 2269.270 2588.280 2269.550 2588.560 ;
        RECT 2303.770 2588.280 2304.050 2588.560 ;
        RECT 2345.170 2588.280 2345.450 2588.560 ;
        RECT 2235.230 2587.600 2235.510 2587.880 ;
        RECT 2242.130 2587.600 2242.410 2587.880 ;
        RECT 2249.030 2587.600 2249.310 2587.880 ;
        RECT 2255.930 2587.600 2256.210 2587.880 ;
        RECT 2262.830 2587.600 2263.110 2587.880 ;
        RECT 2269.730 2587.600 2270.010 2587.880 ;
        RECT 2276.630 2587.600 2276.910 2587.880 ;
        RECT 2283.530 2587.600 2283.810 2587.880 ;
        RECT 2290.430 2587.600 2290.710 2587.880 ;
        RECT 2297.330 2587.600 2297.610 2587.880 ;
        RECT 2304.230 2587.600 2304.510 2587.880 ;
        RECT 2311.130 2587.600 2311.410 2587.880 ;
        RECT 2318.030 2587.600 2318.310 2587.880 ;
        RECT 2324.930 2587.600 2325.210 2587.880 ;
        RECT 2331.830 2587.600 2332.110 2587.880 ;
        RECT 2338.730 2587.600 2339.010 2587.880 ;
        RECT 2338.730 2412.160 2339.010 2412.440 ;
        RECT 2345.630 2587.600 2345.910 2587.880 ;
        RECT 2345.630 2411.480 2345.910 2411.760 ;
        RECT 2559.990 2412.160 2560.270 2412.440 ;
        RECT 2581.610 2411.480 2581.890 2411.760 ;
        RECT 2592.650 2410.800 2592.930 2411.080 ;
        RECT 1441.730 1019.520 1442.010 1019.800 ;
        RECT 1448.630 1018.840 1448.910 1019.120 ;
        RECT 1496.930 1020.200 1497.210 1020.480 ;
        RECT 1646.890 1062.360 1647.170 1062.640 ;
        RECT 1641.830 1016.800 1642.110 1017.080 ;
        RECT 1654.710 1016.800 1654.990 1017.080 ;
        RECT 1641.370 1016.120 1641.650 1016.400 ;
        RECT 1655.630 1016.120 1655.910 1016.400 ;
        RECT 1675.870 1016.800 1676.150 1017.080 ;
        RECT 1662.530 1016.120 1662.810 1016.400 ;
        RECT 1669.430 1016.120 1669.710 1016.400 ;
        RECT 1683.230 1038.560 1683.510 1038.840 ;
        RECT 1683.690 1016.800 1683.970 1017.080 ;
        RECT 1676.330 1016.120 1676.610 1016.400 ;
        RECT 1662.070 1015.440 1662.350 1015.720 ;
        RECT 1668.970 1015.440 1669.250 1015.720 ;
        RECT 1675.410 1015.440 1675.690 1015.720 ;
        RECT 1683.230 1015.440 1683.510 1015.720 ;
        RECT 1704.390 1020.880 1704.670 1021.160 ;
        RECT 1711.290 1018.160 1711.570 1018.440 ;
        RECT 1711.290 1017.480 1711.570 1017.760 ;
        RECT 1691.050 1016.120 1691.330 1016.400 ;
        RECT 1697.950 1016.120 1698.230 1016.400 ;
        RECT 1718.190 1018.160 1718.470 1018.440 ;
        RECT 1752.230 1020.880 1752.510 1021.160 ;
        RECT 1725.090 1016.120 1725.370 1016.400 ;
        RECT 1731.990 1016.120 1732.270 1016.400 ;
        RECT 1738.890 1015.440 1739.170 1015.720 ;
        RECT 1745.790 1018.160 1746.070 1018.440 ;
        RECT 1745.790 1016.120 1746.070 1016.400 ;
        RECT 1755.450 1015.440 1755.730 1015.720 ;
        RECT 1776.610 1019.520 1776.890 1019.800 ;
        RECT 1759.590 1018.160 1759.870 1018.440 ;
        RECT 1766.490 1015.440 1766.770 1015.720 ;
        RECT 1773.390 1018.160 1773.670 1018.440 ;
        RECT 1776.610 1016.800 1776.890 1017.080 ;
        RECT 1786.730 1020.880 1787.010 1021.160 ;
        RECT 1779.830 1017.480 1780.110 1017.760 ;
        RECT 1787.190 1019.520 1787.470 1019.800 ;
        RECT 1780.290 1016.120 1780.570 1016.400 ;
        RECT 1793.630 1018.160 1793.910 1018.440 ;
        RECT 1787.650 1015.440 1787.930 1015.720 ;
        RECT 1834.110 1020.880 1834.390 1021.160 ;
        RECT 1834.570 1020.200 1834.850 1020.480 ;
        RECT 1842.390 1020.880 1842.670 1021.160 ;
        RECT 1855.730 1020.880 1856.010 1021.160 ;
        RECT 1814.330 1018.840 1814.610 1019.120 ;
        RECT 1835.030 1019.520 1835.310 1019.800 ;
        RECT 1821.690 1016.800 1821.970 1017.080 ;
        RECT 1648.730 1014.760 1649.010 1015.040 ;
        RECT 1683.230 1014.760 1683.510 1015.040 ;
        RECT 1689.670 1014.760 1689.950 1015.040 ;
        RECT 1696.110 1014.760 1696.390 1015.040 ;
        RECT 1700.710 1014.760 1700.990 1015.040 ;
        RECT 1707.150 1014.760 1707.430 1015.040 ;
        RECT 1713.590 1014.760 1713.870 1015.040 ;
        RECT 1718.190 1014.760 1718.470 1015.040 ;
        RECT 1724.630 1014.760 1724.910 1015.040 ;
        RECT 1729.690 1014.760 1729.970 1015.040 ;
        RECT 1735.670 1014.760 1735.950 1015.040 ;
        RECT 1741.650 1014.760 1741.930 1015.040 ;
        RECT 1748.090 1014.760 1748.370 1015.040 ;
        RECT 1755.910 1014.760 1756.190 1015.040 ;
        RECT 1759.130 1014.760 1759.410 1015.040 ;
        RECT 1766.030 1014.760 1766.310 1015.040 ;
        RECT 1772.930 1014.760 1773.210 1015.040 ;
        RECT 1777.990 1014.760 1778.270 1015.040 ;
        RECT 1782.130 1014.760 1782.410 1015.040 ;
        RECT 1787.190 1014.760 1787.470 1015.040 ;
        RECT 1790.410 1014.760 1790.690 1015.040 ;
        RECT 1794.090 1014.760 1794.370 1015.040 ;
        RECT 1800.070 1014.760 1800.350 1015.040 ;
        RECT 1806.050 1014.760 1806.330 1015.040 ;
        RECT 1812.950 1014.760 1813.230 1015.040 ;
        RECT 1817.550 1014.760 1817.830 1015.040 ;
        RECT 1823.990 1014.760 1824.270 1015.040 ;
        RECT 1490.030 558.480 1490.310 558.760 ;
        RECT 1503.830 556.440 1504.110 556.720 ;
        RECT 1898.970 913.440 1899.250 913.720 ;
        RECT 1884.250 908.000 1884.530 908.280 ;
        RECT 1899.890 615.600 1900.170 615.880 ;
        RECT 1900.350 590.440 1900.630 590.720 ;
        RECT 1900.350 578.880 1900.630 579.160 ;
        RECT 1902.190 610.160 1902.470 610.440 ;
        RECT 1901.730 601.320 1902.010 601.600 ;
        RECT 1901.270 593.160 1901.550 593.440 ;
        RECT 2242.130 1020.880 2242.410 1021.160 ;
        RECT 2259.610 1020.880 2259.890 1021.160 ;
        RECT 2266.510 1020.880 2266.790 1021.160 ;
        RECT 2245.810 1020.200 2246.090 1020.480 ;
        RECT 2254.550 1020.200 2254.830 1020.480 ;
        RECT 2276.630 1020.880 2276.910 1021.160 ;
        RECT 2273.410 1019.520 2273.690 1019.800 ;
        RECT 2276.630 1019.520 2276.910 1019.800 ;
        RECT 2283.530 1020.880 2283.810 1021.160 ;
        RECT 2281.230 1020.200 2281.510 1020.480 ;
        RECT 2269.730 1016.800 2270.010 1017.080 ;
        RECT 2280.310 1016.800 2280.590 1017.080 ;
        RECT 2283.530 1016.800 2283.810 1017.080 ;
        RECT 2287.210 1016.120 2287.490 1016.400 ;
        RECT 2249.030 1014.760 2249.310 1015.040 ;
        RECT 2255.010 1014.760 2255.290 1015.040 ;
        RECT 2262.830 1014.760 2263.110 1015.040 ;
        RECT 2242.130 1006.600 2242.410 1006.880 ;
        RECT 2296.870 1016.120 2297.150 1016.400 ;
        RECT 2304.230 1016.800 2304.510 1017.080 ;
        RECT 2311.130 1016.120 2311.410 1016.400 ;
        RECT 2317.570 1016.800 2317.850 1017.080 ;
        RECT 2318.030 1016.120 2318.310 1016.400 ;
        RECT 2330.910 1020.880 2331.190 1021.160 ;
        RECT 2338.730 1020.880 2339.010 1021.160 ;
        RECT 2345.170 1020.880 2345.450 1021.160 ;
        RECT 2324.470 1016.120 2324.750 1016.400 ;
        RECT 2289.970 1014.760 2290.250 1015.040 ;
        RECT 2293.650 1014.760 2293.930 1015.040 ;
        RECT 2303.310 1014.760 2303.590 1015.040 ;
        RECT 2307.910 1014.760 2308.190 1015.040 ;
        RECT 2312.050 1014.760 2312.330 1015.040 ;
        RECT 2317.110 1014.760 2317.390 1015.040 ;
        RECT 2323.550 1014.760 2323.830 1015.040 ;
        RECT 2329.530 1014.760 2329.810 1015.040 ;
        RECT 2335.510 1014.760 2335.790 1015.040 ;
        RECT 2342.410 1014.760 2342.690 1015.040 ;
        RECT 2352.530 1020.880 2352.810 1021.160 ;
        RECT 2359.430 1020.880 2359.710 1021.160 ;
        RECT 2351.610 1020.200 2351.890 1020.480 ;
        RECT 2359.890 1020.200 2360.170 1020.480 ;
        RECT 2355.290 1016.120 2355.570 1016.400 ;
        RECT 2373.690 1020.880 2373.970 1021.160 ;
        RECT 2403.130 1020.880 2403.410 1021.160 ;
        RECT 2380.590 1020.200 2380.870 1020.480 ;
        RECT 2387.490 1020.200 2387.770 1020.480 ;
        RECT 2387.950 1016.800 2388.230 1017.080 ;
        RECT 2381.050 1016.120 2381.330 1016.400 ;
        RECT 2408.190 1018.160 2408.470 1018.440 ;
        RECT 2408.190 1017.480 2408.470 1017.760 ;
        RECT 2421.990 1020.880 2422.270 1021.160 ;
        RECT 2450.970 1020.200 2451.250 1020.480 ;
        RECT 2428.890 1018.160 2429.170 1018.440 ;
        RECT 2394.390 1016.800 2394.670 1017.080 ;
        RECT 2415.090 1016.800 2415.370 1017.080 ;
        RECT 2421.990 1016.800 2422.270 1017.080 ;
        RECT 2388.410 1016.120 2388.690 1016.400 ;
        RECT 2347.010 1014.760 2347.290 1015.040 ;
        RECT 2355.750 1014.760 2356.030 1015.040 ;
        RECT 2363.570 1014.760 2363.850 1015.040 ;
        RECT 2366.790 1014.760 2367.070 1015.040 ;
        RECT 2373.230 1014.760 2373.510 1015.040 ;
        RECT 2377.830 1014.760 2378.110 1015.040 ;
        RECT 2380.590 1014.760 2380.870 1015.040 ;
        RECT 2387.490 1014.760 2387.770 1015.040 ;
        RECT 2394.390 1014.760 2394.670 1015.040 ;
        RECT 2402.210 1014.760 2402.490 1015.040 ;
        RECT 2415.090 1014.760 2415.370 1015.040 ;
        RECT 1900.810 573.440 1901.090 573.720 ;
        RECT 2083.890 556.440 2084.170 556.720 ;
        RECT 2482.250 906.640 2482.530 906.920 ;
        RECT 2504.330 915.480 2504.610 915.760 ;
        RECT 2500.650 618.320 2500.930 618.600 ;
        RECT 2500.190 610.160 2500.470 610.440 ;
        RECT 2499.730 604.040 2500.010 604.320 ;
        RECT 2499.270 593.160 2499.550 593.440 ;
        RECT 2498.810 590.440 2499.090 590.720 ;
        RECT 2498.350 578.880 2498.630 579.160 ;
        RECT 2497.890 576.160 2498.170 576.440 ;
      LAYER met3 ;
        RECT 1868.125 3063.900 1868.455 3063.905 ;
        RECT 1867.870 3063.890 1868.455 3063.900 ;
        RECT 2442.665 3063.900 2442.995 3063.905 ;
        RECT 2469.805 3063.900 2470.135 3063.905 ;
        RECT 2442.665 3063.890 2443.250 3063.900 ;
        RECT 2469.550 3063.890 2470.135 3063.900 ;
        RECT 1867.870 3063.590 1868.680 3063.890 ;
        RECT 2442.665 3063.590 2443.450 3063.890 ;
        RECT 2469.350 3063.590 2470.135 3063.890 ;
        RECT 1867.870 3063.580 1868.455 3063.590 ;
        RECT 1868.125 3063.575 1868.455 3063.580 ;
        RECT 2442.665 3063.580 2443.250 3063.590 ;
        RECT 2469.550 3063.580 2470.135 3063.590 ;
        RECT 2442.665 3063.575 2442.995 3063.580 ;
        RECT 2469.805 3063.575 2470.135 3063.580 ;
        RECT 1845.790 3055.050 1846.170 3055.060 ;
        RECT 1865.110 3055.050 1865.490 3055.060 ;
        RECT 1845.790 3054.750 1865.490 3055.050 ;
        RECT 1845.790 3054.740 1846.170 3054.750 ;
        RECT 1865.110 3054.740 1865.490 3054.750 ;
        RECT 1859.280 3051.235 1861.020 3052.140 ;
        RECT 2459.280 3051.235 2461.020 3052.140 ;
        RECT 1490.005 3033.290 1490.335 3033.305 ;
        RECT 1490.005 3033.085 1497.450 3033.290 ;
        RECT 1490.005 3032.990 1504.600 3033.085 ;
        RECT 1490.005 3032.975 1490.335 3032.990 ;
        RECT 1497.150 3032.785 1504.600 3032.990 ;
        RECT 1489.545 3027.170 1489.875 3027.185 ;
        RECT 1497.150 3027.170 1504.600 3027.445 ;
        RECT 1489.545 3027.145 1504.600 3027.170 ;
        RECT 1489.545 3026.870 1497.450 3027.145 ;
        RECT 1489.545 3026.855 1489.875 3026.870 ;
        RECT 1489.085 3019.010 1489.415 3019.025 ;
        RECT 1489.085 3018.945 1497.450 3019.010 ;
        RECT 1489.085 3018.710 1504.600 3018.945 ;
        RECT 1489.085 3018.695 1489.415 3018.710 ;
        RECT 1497.150 3018.645 1504.600 3018.710 ;
        RECT 1497.150 3013.005 1504.600 3013.305 ;
        RECT 1488.625 3012.890 1488.955 3012.905 ;
        RECT 1497.150 3012.890 1497.450 3013.005 ;
        RECT 1488.625 3012.590 1497.450 3012.890 ;
        RECT 1488.625 3012.575 1488.955 3012.590 ;
        RECT 1488.165 3004.730 1488.495 3004.745 ;
        RECT 1497.150 3004.730 1504.600 3004.805 ;
        RECT 1488.165 3004.505 1504.600 3004.730 ;
        RECT 1488.165 3004.430 1497.450 3004.505 ;
        RECT 1488.165 3004.415 1488.495 3004.430 ;
        RECT 1487.705 2999.290 1488.035 2999.305 ;
        RECT 1487.705 2999.165 1497.450 2999.290 ;
        RECT 1487.705 2998.990 1504.600 2999.165 ;
        RECT 1487.705 2998.975 1488.035 2998.990 ;
        RECT 1497.150 2998.865 1504.600 2998.990 ;
        RECT 1487.245 2990.450 1487.575 2990.465 ;
        RECT 1497.150 2990.450 1504.600 2990.665 ;
        RECT 1487.245 2990.365 1504.600 2990.450 ;
        RECT 1487.245 2990.150 1497.450 2990.365 ;
        RECT 1487.245 2990.135 1487.575 2990.150 ;
        RECT 1486.785 2701.450 1487.115 2701.465 ;
        RECT 1486.785 2701.425 1497.450 2701.450 ;
        RECT 1486.785 2701.150 1504.600 2701.425 ;
        RECT 1486.785 2701.135 1487.115 2701.150 ;
        RECT 1497.150 2701.125 1504.600 2701.150 ;
        RECT 1497.150 2692.625 1504.600 2692.925 ;
        RECT 1486.325 2692.610 1486.655 2692.625 ;
        RECT 1497.150 2692.610 1497.450 2692.625 ;
        RECT 1486.325 2692.310 1497.450 2692.610 ;
        RECT 1486.325 2692.295 1486.655 2692.310 ;
      LAYER met3 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
      LAYER met3 ;
        RECT 1881.880 3048.265 1889.370 3048.565 ;
        RECT 1889.070 3048.250 1889.370 3048.265 ;
        RECT 1898.485 3048.250 1898.815 3048.265 ;
        RECT 1899.865 3048.250 1900.195 3048.265 ;
        RECT 1889.070 3047.950 1900.195 3048.250 ;
        RECT 1898.485 3047.935 1898.815 3047.950 ;
        RECT 1899.865 3047.935 1900.195 3047.950 ;
        RECT 2100.000 3032.785 2104.600 3033.085 ;
        RECT 2087.085 3031.250 2087.415 3031.265 ;
        RECT 2100.670 3031.250 2100.970 3032.785 ;
        RECT 2087.085 3030.950 2100.970 3031.250 ;
        RECT 2087.085 3030.935 2087.415 3030.950 ;
        RECT 2100.000 3027.145 2104.600 3027.445 ;
        RECT 2087.545 3024.450 2087.875 3024.465 ;
        RECT 2100.670 3024.450 2100.970 3027.145 ;
        RECT 2087.545 3024.150 2100.970 3024.450 ;
        RECT 2087.545 3024.135 2087.875 3024.150 ;
        RECT 2100.000 3018.645 2104.600 3018.945 ;
        RECT 2088.005 3016.290 2088.335 3016.305 ;
        RECT 2100.670 3016.290 2100.970 3018.645 ;
        RECT 2088.005 3015.990 2100.970 3016.290 ;
        RECT 2088.005 3015.975 2088.335 3015.990 ;
        RECT 2100.000 3013.005 2104.600 3013.305 ;
        RECT 2088.465 3010.170 2088.795 3010.185 ;
        RECT 2100.670 3010.170 2100.970 3013.005 ;
        RECT 2088.465 3009.870 2100.970 3010.170 ;
        RECT 2088.465 3009.855 2088.795 3009.870 ;
        RECT 2100.000 3004.505 2104.600 3004.805 ;
        RECT 2088.925 3002.010 2089.255 3002.025 ;
        RECT 2100.670 3002.010 2100.970 3004.505 ;
        RECT 2088.925 3001.710 2100.970 3002.010 ;
        RECT 2088.925 3001.695 2089.255 3001.710 ;
        RECT 2100.000 2998.865 2104.600 2999.165 ;
        RECT 2089.385 2996.570 2089.715 2996.585 ;
        RECT 2100.670 2996.570 2100.970 2998.865 ;
        RECT 2089.385 2996.270 2100.970 2996.570 ;
        RECT 2089.385 2996.255 2089.715 2996.270 ;
        RECT 2100.000 2990.365 2104.600 2990.665 ;
        RECT 2089.845 2988.410 2090.175 2988.425 ;
        RECT 2100.670 2988.410 2100.970 2990.365 ;
        RECT 2089.845 2988.110 2100.970 2988.410 ;
        RECT 2089.845 2988.095 2090.175 2988.110 ;
        RECT 1881.880 2747.010 1889.370 2747.210 ;
        RECT 1898.025 2747.010 1898.355 2747.025 ;
        RECT 1881.880 2746.910 1898.355 2747.010 ;
        RECT 1885.390 2738.710 1885.690 2746.910 ;
        RECT 1889.070 2746.710 1898.355 2746.910 ;
        RECT 1898.025 2746.695 1898.355 2746.710 ;
        RECT 1881.880 2738.410 1886.480 2738.710 ;
        RECT 1885.390 2733.070 1885.690 2738.410 ;
        RECT 1881.880 2732.770 1886.480 2733.070 ;
        RECT 1885.390 2724.570 1885.690 2732.770 ;
        RECT 1881.880 2724.270 1886.480 2724.570 ;
        RECT 1885.390 2718.930 1885.690 2724.270 ;
        RECT 1881.880 2718.630 1886.480 2718.930 ;
        RECT 1885.390 2710.430 1885.690 2718.630 ;
        RECT 1881.880 2710.130 1886.480 2710.430 ;
        RECT 1885.390 2704.790 1885.690 2710.130 ;
        RECT 1898.025 2704.850 1898.355 2704.865 ;
        RECT 1887.230 2704.790 1898.355 2704.850 ;
        RECT 1881.880 2704.550 1898.355 2704.790 ;
        RECT 1881.880 2704.490 1887.530 2704.550 ;
        RECT 1898.025 2704.535 1898.355 2704.550 ;
        RECT 2100.000 2701.125 2104.600 2701.425 ;
        RECT 2083.865 2699.410 2084.195 2699.425 ;
        RECT 2100.670 2699.410 2100.970 2701.125 ;
        RECT 2083.865 2699.110 2100.970 2699.410 ;
        RECT 2083.865 2699.095 2084.195 2699.110 ;
        RECT 2100.000 2692.625 2104.600 2692.925 ;
        RECT 2090.305 2691.930 2090.635 2691.945 ;
        RECT 2100.670 2691.930 2100.970 2692.625 ;
        RECT 2090.305 2691.630 2100.970 2691.930 ;
        RECT 2090.305 2691.615 2090.635 2691.630 ;
      LAYER met3 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
      LAYER met3 ;
        RECT 2482.225 3049.610 2482.555 3049.625 ;
        RECT 2482.225 3049.295 2482.770 3049.610 ;
        RECT 2482.470 3048.565 2482.770 3049.295 ;
        RECT 2481.880 3048.265 2486.480 3048.565 ;
        RECT 2497.865 2747.690 2498.195 2747.705 ;
        RECT 2488.910 2747.390 2498.195 2747.690 ;
        RECT 2488.910 2747.210 2489.210 2747.390 ;
        RECT 2497.865 2747.375 2498.195 2747.390 ;
        RECT 2481.880 2746.910 2489.210 2747.210 ;
        RECT 2485.230 2739.530 2485.530 2746.910 ;
        RECT 2485.230 2739.230 2486.450 2739.530 ;
        RECT 2486.150 2738.710 2486.450 2739.230 ;
        RECT 2481.880 2738.410 2486.480 2738.710 ;
        RECT 2486.150 2733.070 2486.450 2738.410 ;
        RECT 2481.880 2732.770 2486.480 2733.070 ;
        RECT 2486.150 2724.570 2486.450 2732.770 ;
        RECT 2481.880 2724.270 2486.480 2724.570 ;
        RECT 2486.150 2718.930 2486.450 2724.270 ;
        RECT 2481.880 2718.630 2486.480 2718.930 ;
        RECT 2486.150 2710.430 2486.450 2718.630 ;
        RECT 2481.880 2710.290 2486.480 2710.430 ;
        RECT 2497.865 2710.290 2498.195 2710.305 ;
        RECT 2481.880 2710.130 2498.195 2710.290 ;
        RECT 2486.150 2709.990 2498.195 2710.130 ;
        RECT 2497.865 2709.975 2498.195 2709.990 ;
        RECT 2497.865 2704.850 2498.195 2704.865 ;
        RECT 2486.150 2704.790 2498.195 2704.850 ;
        RECT 2481.880 2704.550 2498.195 2704.790 ;
        RECT 2481.880 2704.490 2486.480 2704.550 ;
        RECT 2497.865 2704.535 2498.195 2704.550 ;
        RECT 2126.645 2598.770 2126.975 2598.785 ;
        RECT 2139.810 2598.770 2140.190 2598.780 ;
        RECT 2126.645 2598.470 2140.190 2598.770 ;
        RECT 2126.645 2598.455 2126.975 2598.470 ;
        RECT 2139.810 2598.460 2140.190 2598.470 ;
        RECT 1568.870 2594.010 1569.250 2594.020 ;
        RECT 1569.585 2594.010 1569.915 2594.025 ;
        RECT 1573.725 2594.020 1574.055 2594.025 ;
        RECT 1573.470 2594.010 1574.055 2594.020 ;
        RECT 1568.870 2593.710 1569.915 2594.010 ;
        RECT 1573.270 2593.710 1574.055 2594.010 ;
        RECT 1568.870 2593.700 1569.250 2593.710 ;
        RECT 1569.585 2593.695 1569.915 2593.710 ;
        RECT 1573.470 2593.700 1574.055 2593.710 ;
        RECT 1580.830 2594.010 1581.210 2594.020 ;
        RECT 1586.605 2594.010 1586.935 2594.025 ;
        RECT 1591.205 2594.020 1591.535 2594.025 ;
        RECT 1598.565 2594.020 1598.895 2594.025 ;
        RECT 1604.085 2594.020 1604.415 2594.025 ;
        RECT 1590.950 2594.010 1591.535 2594.020 ;
        RECT 1598.310 2594.010 1598.895 2594.020 ;
        RECT 1603.830 2594.010 1604.415 2594.020 ;
        RECT 1580.830 2593.710 1586.935 2594.010 ;
        RECT 1590.750 2593.710 1591.535 2594.010 ;
        RECT 1598.110 2593.710 1598.895 2594.010 ;
        RECT 1603.630 2593.710 1604.415 2594.010 ;
        RECT 1580.830 2593.700 1581.210 2593.710 ;
        RECT 1573.725 2593.695 1574.055 2593.700 ;
        RECT 1586.605 2593.695 1586.935 2593.710 ;
        RECT 1590.950 2593.700 1591.535 2593.710 ;
        RECT 1598.310 2593.700 1598.895 2593.710 ;
        RECT 1603.830 2593.700 1604.415 2593.710 ;
        RECT 1591.205 2593.695 1591.535 2593.700 ;
        RECT 1598.565 2593.695 1598.895 2593.700 ;
        RECT 1604.085 2593.695 1604.415 2593.700 ;
        RECT 1614.665 2594.020 1614.995 2594.025 ;
        RECT 1614.665 2594.010 1615.250 2594.020 ;
        RECT 1621.565 2594.010 1621.895 2594.025 ;
        RECT 1626.625 2594.020 1626.955 2594.025 ;
        RECT 1651.005 2594.020 1651.335 2594.025 ;
        RECT 1622.230 2594.010 1622.610 2594.020 ;
        RECT 1614.665 2593.710 1615.450 2594.010 ;
        RECT 1621.565 2593.710 1622.610 2594.010 ;
        RECT 1614.665 2593.700 1615.250 2593.710 ;
        RECT 1614.665 2593.695 1614.995 2593.700 ;
        RECT 1621.565 2593.695 1621.895 2593.710 ;
        RECT 1622.230 2593.700 1622.610 2593.710 ;
        RECT 1626.625 2594.010 1627.210 2594.020 ;
        RECT 1650.750 2594.010 1651.335 2594.020 ;
        RECT 1626.625 2593.710 1627.410 2594.010 ;
        RECT 1650.550 2593.710 1651.335 2594.010 ;
        RECT 1626.625 2593.700 1627.210 2593.710 ;
        RECT 1650.750 2593.700 1651.335 2593.710 ;
        RECT 1626.625 2593.695 1626.955 2593.700 ;
        RECT 1651.005 2593.695 1651.335 2593.700 ;
        RECT 1661.585 2594.020 1661.915 2594.025 ;
        RECT 1661.585 2594.010 1662.170 2594.020 ;
        RECT 1669.865 2594.010 1670.195 2594.025 ;
        RECT 1690.565 2594.020 1690.895 2594.025 ;
        RECT 1670.990 2594.010 1671.370 2594.020 ;
        RECT 1690.310 2594.010 1690.895 2594.020 ;
        RECT 1661.585 2593.710 1662.370 2594.010 ;
        RECT 1669.865 2593.710 1671.370 2594.010 ;
        RECT 1690.110 2593.710 1690.895 2594.010 ;
        RECT 1661.585 2593.700 1662.170 2593.710 ;
        RECT 1661.585 2593.695 1661.915 2593.700 ;
        RECT 1669.865 2593.695 1670.195 2593.710 ;
        RECT 1670.990 2593.700 1671.370 2593.710 ;
        RECT 1690.310 2593.700 1690.895 2593.710 ;
        RECT 1696.750 2594.010 1697.130 2594.020 ;
        RECT 1697.925 2594.010 1698.255 2594.025 ;
        RECT 1738.405 2594.020 1738.735 2594.025 ;
        RECT 2215.885 2594.020 2216.215 2594.025 ;
        RECT 2256.365 2594.020 2256.695 2594.025 ;
        RECT 2262.805 2594.020 2263.135 2594.025 ;
        RECT 2268.325 2594.020 2268.655 2594.025 ;
        RECT 1738.150 2594.010 1738.735 2594.020 ;
        RECT 2215.630 2594.010 2216.215 2594.020 ;
        RECT 1696.750 2593.710 1698.255 2594.010 ;
        RECT 1737.950 2593.710 1738.735 2594.010 ;
        RECT 2215.430 2593.710 2216.215 2594.010 ;
        RECT 1696.750 2593.700 1697.130 2593.710 ;
        RECT 1690.565 2593.695 1690.895 2593.700 ;
        RECT 1697.925 2593.695 1698.255 2593.710 ;
        RECT 1738.150 2593.700 1738.735 2593.710 ;
        RECT 2215.630 2593.700 2216.215 2593.710 ;
        RECT 2256.110 2594.010 2256.695 2594.020 ;
        RECT 2262.550 2594.010 2263.135 2594.020 ;
        RECT 2268.070 2594.010 2268.655 2594.020 ;
        RECT 2256.110 2593.710 2256.920 2594.010 ;
        RECT 2262.350 2593.710 2263.135 2594.010 ;
        RECT 2267.870 2593.710 2268.655 2594.010 ;
        RECT 2256.110 2593.700 2256.695 2593.710 ;
        RECT 2262.550 2593.700 2263.135 2593.710 ;
        RECT 2268.070 2593.700 2268.655 2593.710 ;
        RECT 1738.405 2593.695 1738.735 2593.700 ;
        RECT 2215.885 2593.695 2216.215 2593.700 ;
        RECT 2256.365 2593.695 2256.695 2593.700 ;
        RECT 2262.805 2593.695 2263.135 2593.700 ;
        RECT 2268.325 2593.695 2268.655 2593.700 ;
        RECT 2297.765 2594.010 2298.095 2594.025 ;
        RECT 2302.110 2594.010 2302.490 2594.020 ;
        RECT 2297.765 2593.710 2302.490 2594.010 ;
        RECT 2297.765 2593.695 2298.095 2593.710 ;
        RECT 2302.110 2593.700 2302.490 2593.710 ;
        RECT 2305.125 2594.010 2305.455 2594.025 ;
        RECT 2305.790 2594.010 2306.170 2594.020 ;
        RECT 2305.125 2593.710 2306.170 2594.010 ;
        RECT 2305.125 2593.695 2305.455 2593.710 ;
        RECT 2305.790 2593.700 2306.170 2593.710 ;
        RECT 1581.085 2593.330 1581.415 2593.345 ;
        RECT 1587.065 2593.340 1587.395 2593.345 ;
        RECT 1639.045 2593.340 1639.375 2593.345 ;
        RECT 1644.565 2593.340 1644.895 2593.345 ;
        RECT 1582.670 2593.330 1583.050 2593.340 ;
        RECT 1587.065 2593.330 1587.650 2593.340 ;
        RECT 1638.790 2593.330 1639.375 2593.340 ;
        RECT 1644.310 2593.330 1644.895 2593.340 ;
        RECT 1581.085 2593.030 1583.050 2593.330 ;
        RECT 1586.840 2593.030 1587.650 2593.330 ;
        RECT 1638.590 2593.030 1639.375 2593.330 ;
        RECT 1644.110 2593.030 1644.895 2593.330 ;
        RECT 1581.085 2593.015 1581.415 2593.030 ;
        RECT 1582.670 2593.020 1583.050 2593.030 ;
        RECT 1587.065 2593.020 1587.650 2593.030 ;
        RECT 1638.790 2593.020 1639.375 2593.030 ;
        RECT 1644.310 2593.020 1644.895 2593.030 ;
        RECT 1587.065 2593.015 1587.395 2593.020 ;
        RECT 1639.045 2593.015 1639.375 2593.020 ;
        RECT 1644.565 2593.015 1644.895 2593.020 ;
        RECT 1656.065 2593.340 1656.395 2593.345 ;
        RECT 1679.525 2593.340 1679.855 2593.345 ;
        RECT 1656.065 2593.330 1656.650 2593.340 ;
        RECT 1679.270 2593.330 1679.855 2593.340 ;
        RECT 1656.065 2593.030 1656.850 2593.330 ;
        RECT 1679.070 2593.030 1679.855 2593.330 ;
        RECT 1656.065 2593.020 1656.650 2593.030 ;
        RECT 1679.270 2593.020 1679.855 2593.030 ;
        RECT 1656.065 2593.015 1656.395 2593.020 ;
        RECT 1679.525 2593.015 1679.855 2593.020 ;
        RECT 1707.585 2593.340 1707.915 2593.345 ;
        RECT 1732.885 2593.340 1733.215 2593.345 ;
        RECT 1743.925 2593.340 1744.255 2593.345 ;
        RECT 1707.585 2593.330 1708.170 2593.340 ;
        RECT 1732.630 2593.330 1733.215 2593.340 ;
        RECT 1743.670 2593.330 1744.255 2593.340 ;
        RECT 1707.585 2593.030 1708.370 2593.330 ;
        RECT 1732.430 2593.030 1733.215 2593.330 ;
        RECT 1743.470 2593.030 1744.255 2593.330 ;
        RECT 1707.585 2593.020 1708.170 2593.030 ;
        RECT 1732.630 2593.020 1733.215 2593.030 ;
        RECT 1743.670 2593.020 1744.255 2593.030 ;
        RECT 1707.585 2593.015 1707.915 2593.020 ;
        RECT 1732.885 2593.015 1733.215 2593.020 ;
        RECT 1743.925 2593.015 1744.255 2593.020 ;
        RECT 2146.425 2593.330 2146.755 2593.345 ;
        RECT 2220.485 2593.340 2220.815 2593.345 ;
        RECT 2148.470 2593.330 2148.850 2593.340 ;
        RECT 2220.230 2593.330 2220.815 2593.340 ;
        RECT 2146.425 2593.030 2148.850 2593.330 ;
        RECT 2220.030 2593.030 2220.815 2593.330 ;
        RECT 2146.425 2593.015 2146.755 2593.030 ;
        RECT 2148.470 2593.020 2148.850 2593.030 ;
        RECT 2220.230 2593.020 2220.815 2593.030 ;
        RECT 2220.485 2593.015 2220.815 2593.020 ;
        RECT 2291.785 2593.340 2292.115 2593.345 ;
        RECT 2297.765 2593.340 2298.095 2593.345 ;
        RECT 2291.785 2593.330 2292.370 2593.340 ;
        RECT 2297.510 2593.330 2298.095 2593.340 ;
        RECT 2291.785 2593.030 2292.570 2593.330 ;
        RECT 2297.310 2593.030 2298.095 2593.330 ;
        RECT 2291.785 2593.020 2292.370 2593.030 ;
        RECT 2297.510 2593.020 2298.095 2593.030 ;
        RECT 2291.785 2593.015 2292.115 2593.020 ;
        RECT 2297.765 2593.015 2298.095 2593.020 ;
        RECT 2311.565 2593.330 2311.895 2593.345 ;
        RECT 2312.230 2593.330 2312.610 2593.340 ;
        RECT 2311.565 2593.030 2312.610 2593.330 ;
        RECT 2311.565 2593.015 2311.895 2593.030 ;
        RECT 2312.230 2593.020 2312.610 2593.030 ;
        RECT 2332.265 2593.330 2332.595 2593.345 ;
        RECT 2337.070 2593.330 2337.450 2593.340 ;
        RECT 2332.265 2593.030 2337.450 2593.330 ;
        RECT 2332.265 2593.015 2332.595 2593.030 ;
        RECT 2337.070 2593.020 2337.450 2593.030 ;
        RECT 1562.430 2592.650 1562.810 2592.660 ;
        RECT 1565.445 2592.650 1565.775 2592.665 ;
        RECT 1562.430 2592.350 1565.775 2592.650 ;
        RECT 1562.430 2592.340 1562.810 2592.350 ;
        RECT 1565.445 2592.335 1565.775 2592.350 ;
        RECT 1573.265 2592.650 1573.595 2592.665 ;
        RECT 1608.225 2592.660 1608.555 2592.665 ;
        RECT 1621.565 2592.660 1621.895 2592.665 ;
        RECT 1633.525 2592.660 1633.855 2592.665 ;
        RECT 1575.310 2592.650 1575.690 2592.660 ;
        RECT 1573.265 2592.350 1575.690 2592.650 ;
        RECT 1573.265 2592.335 1573.595 2592.350 ;
        RECT 1575.310 2592.340 1575.690 2592.350 ;
        RECT 1608.225 2592.650 1608.810 2592.660 ;
        RECT 1621.310 2592.650 1621.895 2592.660 ;
        RECT 1633.270 2592.650 1633.855 2592.660 ;
        RECT 1608.225 2592.350 1609.010 2592.650 ;
        RECT 1621.110 2592.350 1621.895 2592.650 ;
        RECT 1633.070 2592.350 1633.855 2592.650 ;
        RECT 1608.225 2592.340 1608.810 2592.350 ;
        RECT 1621.310 2592.340 1621.895 2592.350 ;
        RECT 1633.270 2592.340 1633.855 2592.350 ;
        RECT 1608.225 2592.335 1608.555 2592.340 ;
        RECT 1621.565 2592.335 1621.895 2592.340 ;
        RECT 1633.525 2592.335 1633.855 2592.340 ;
        RECT 1667.105 2592.660 1667.435 2592.665 ;
        RECT 1685.505 2592.660 1685.835 2592.665 ;
        RECT 1702.525 2592.660 1702.855 2592.665 ;
        RECT 1725.525 2592.660 1725.855 2592.665 ;
        RECT 1667.105 2592.650 1667.690 2592.660 ;
        RECT 1685.505 2592.650 1686.090 2592.660 ;
        RECT 1702.270 2592.650 1702.855 2592.660 ;
        RECT 1725.270 2592.650 1725.855 2592.660 ;
        RECT 1667.105 2592.350 1667.890 2592.650 ;
        RECT 1685.505 2592.350 1686.290 2592.650 ;
        RECT 1702.070 2592.350 1702.855 2592.650 ;
        RECT 1725.070 2592.350 1725.855 2592.650 ;
        RECT 1667.105 2592.340 1667.690 2592.350 ;
        RECT 1685.505 2592.340 1686.090 2592.350 ;
        RECT 1702.270 2592.340 1702.855 2592.350 ;
        RECT 1725.270 2592.340 1725.855 2592.350 ;
        RECT 1667.105 2592.335 1667.435 2592.340 ;
        RECT 1685.505 2592.335 1685.835 2592.340 ;
        RECT 1702.525 2592.335 1702.855 2592.340 ;
        RECT 1725.525 2592.335 1725.855 2592.340 ;
        RECT 2152.865 2592.650 2153.195 2592.665 ;
        RECT 2153.990 2592.650 2154.370 2592.660 ;
        RECT 2152.865 2592.350 2154.370 2592.650 ;
        RECT 2152.865 2592.335 2153.195 2592.350 ;
        RECT 2153.990 2592.340 2154.370 2592.350 ;
        RECT 2235.665 2592.650 2235.995 2592.665 ;
        RECT 2249.465 2592.660 2249.795 2592.665 ;
        RECT 2280.285 2592.660 2280.615 2592.665 ;
        RECT 2238.630 2592.650 2239.010 2592.660 ;
        RECT 2235.665 2592.350 2239.010 2592.650 ;
        RECT 2235.665 2592.335 2235.995 2592.350 ;
        RECT 2238.630 2592.340 2239.010 2592.350 ;
        RECT 2249.465 2592.650 2250.050 2592.660 ;
        RECT 2280.030 2592.650 2280.615 2592.660 ;
        RECT 2249.465 2592.350 2250.250 2592.650 ;
        RECT 2279.830 2592.350 2280.615 2592.650 ;
        RECT 2249.465 2592.340 2250.050 2592.350 ;
        RECT 2280.030 2592.340 2280.615 2592.350 ;
        RECT 2249.465 2592.335 2249.795 2592.340 ;
        RECT 2280.285 2592.335 2280.615 2592.340 ;
        RECT 2285.345 2592.660 2285.675 2592.665 ;
        RECT 2285.345 2592.650 2285.930 2592.660 ;
        RECT 2339.165 2592.650 2339.495 2592.665 ;
        RECT 2342.590 2592.650 2342.970 2592.660 ;
        RECT 2285.345 2592.350 2286.130 2592.650 ;
        RECT 2339.165 2592.350 2342.970 2592.650 ;
        RECT 2285.345 2592.340 2285.930 2592.350 ;
        RECT 2285.345 2592.335 2285.675 2592.340 ;
        RECT 2339.165 2592.335 2339.495 2592.350 ;
        RECT 2342.590 2592.340 2342.970 2592.350 ;
        RECT 1607.765 2591.970 1608.095 2591.985 ;
        RECT 1610.270 2591.970 1610.650 2591.980 ;
        RECT 1607.765 2591.670 1610.650 2591.970 ;
        RECT 1607.765 2591.655 1608.095 2591.670 ;
        RECT 1610.270 2591.660 1610.650 2591.670 ;
        RECT 1713.105 2591.970 1713.435 2591.985 ;
        RECT 1715.150 2591.970 1715.530 2591.980 ;
        RECT 1713.105 2591.670 1715.530 2591.970 ;
        RECT 1713.105 2591.655 1713.435 2591.670 ;
        RECT 1715.150 2591.660 1715.530 2591.670 ;
        RECT 1718.165 2591.970 1718.495 2591.985 ;
        RECT 2145.965 2591.980 2146.295 2591.985 ;
        RECT 1718.830 2591.970 1719.210 2591.980 ;
        RECT 1718.165 2591.670 1719.210 2591.970 ;
        RECT 1718.165 2591.655 1718.495 2591.670 ;
        RECT 1718.830 2591.660 1719.210 2591.670 ;
        RECT 2145.710 2591.970 2146.295 2591.980 ;
        RECT 2232.905 2591.980 2233.235 2591.985 ;
        RECT 2243.945 2591.980 2244.275 2591.985 ;
        RECT 2232.905 2591.970 2233.490 2591.980 ;
        RECT 2243.945 2591.970 2244.530 2591.980 ;
        RECT 2273.590 2591.970 2273.970 2591.980 ;
        RECT 2276.145 2591.970 2276.475 2591.985 ;
        RECT 2145.710 2591.670 2146.520 2591.970 ;
        RECT 2232.905 2591.670 2233.690 2591.970 ;
        RECT 2243.945 2591.670 2244.730 2591.970 ;
        RECT 2273.590 2591.670 2276.475 2591.970 ;
        RECT 2145.710 2591.660 2146.295 2591.670 ;
        RECT 2145.965 2591.655 2146.295 2591.660 ;
        RECT 2232.905 2591.660 2233.490 2591.670 ;
        RECT 2243.945 2591.660 2244.530 2591.670 ;
        RECT 2273.590 2591.660 2273.970 2591.670 ;
        RECT 2232.905 2591.655 2233.235 2591.660 ;
        RECT 2243.945 2591.655 2244.275 2591.660 ;
        RECT 2276.145 2591.655 2276.475 2591.670 ;
        RECT 2318.465 2591.970 2318.795 2591.985 ;
        RECT 2332.265 2591.980 2332.595 2591.985 ;
        RECT 2319.590 2591.970 2319.970 2591.980 ;
        RECT 2332.265 2591.970 2332.850 2591.980 ;
        RECT 2318.465 2591.670 2319.970 2591.970 ;
        RECT 2332.040 2591.670 2332.850 2591.970 ;
        RECT 2318.465 2591.655 2318.795 2591.670 ;
        RECT 2319.590 2591.660 2319.970 2591.670 ;
        RECT 2332.265 2591.660 2332.850 2591.670 ;
        RECT 2332.265 2591.655 2332.595 2591.660 ;
        RECT 1586.145 2591.300 1586.475 2591.305 ;
        RECT 1586.145 2591.290 1586.730 2591.300 ;
        RECT 1614.665 2591.290 1614.995 2591.305 ;
        RECT 2209.445 2591.300 2209.775 2591.305 ;
        RECT 1616.710 2591.290 1617.090 2591.300 ;
        RECT 2209.190 2591.290 2209.775 2591.300 ;
        RECT 1586.145 2590.990 1586.930 2591.290 ;
        RECT 1614.665 2590.990 1617.090 2591.290 ;
        RECT 2208.990 2590.990 2209.775 2591.290 ;
        RECT 1586.145 2590.980 1586.730 2590.990 ;
        RECT 1586.145 2590.975 1586.475 2590.980 ;
        RECT 1614.665 2590.975 1614.995 2590.990 ;
        RECT 1616.710 2590.980 1617.090 2590.990 ;
        RECT 2209.190 2590.980 2209.775 2590.990 ;
        RECT 2226.670 2591.290 2227.050 2591.300 ;
        RECT 2227.845 2591.290 2228.175 2591.305 ;
        RECT 2226.670 2590.990 2228.175 2591.290 ;
        RECT 2226.670 2590.980 2227.050 2590.990 ;
        RECT 2209.445 2590.975 2209.775 2590.980 ;
        RECT 2227.845 2590.975 2228.175 2590.990 ;
        RECT 2325.365 2591.290 2325.695 2591.305 ;
        RECT 2326.030 2591.290 2326.410 2591.300 ;
        RECT 2325.365 2590.990 2326.410 2591.290 ;
        RECT 2325.365 2590.975 2325.695 2590.990 ;
        RECT 2326.030 2590.980 2326.410 2590.990 ;
        RECT 1593.965 2590.610 1594.295 2590.625 ;
        RECT 1599.230 2590.610 1599.610 2590.620 ;
        RECT 1593.965 2590.310 1599.610 2590.610 ;
        RECT 1593.965 2590.295 1594.295 2590.310 ;
        RECT 1599.230 2590.300 1599.610 2590.310 ;
        RECT 1656.065 2590.610 1656.395 2590.625 ;
        RECT 1657.190 2590.610 1657.570 2590.620 ;
        RECT 1656.065 2590.310 1657.570 2590.610 ;
        RECT 1656.065 2590.295 1656.395 2590.310 ;
        RECT 1657.190 2590.300 1657.570 2590.310 ;
        RECT 1678.605 2590.610 1678.935 2590.625 ;
        RECT 1680.190 2590.610 1680.570 2590.620 ;
        RECT 1678.605 2590.310 1680.570 2590.610 ;
        RECT 1678.605 2590.295 1678.935 2590.310 ;
        RECT 1680.190 2590.300 1680.570 2590.310 ;
        RECT 2132.165 2590.610 2132.495 2590.625 ;
        RECT 2132.830 2590.610 2133.210 2590.620 ;
        RECT 2132.165 2590.310 2133.210 2590.610 ;
        RECT 2132.165 2590.295 2132.495 2590.310 ;
        RECT 2132.830 2590.300 2133.210 2590.310 ;
        RECT 2175.150 2590.610 2175.530 2590.620 ;
        RECT 2176.785 2590.610 2177.115 2590.625 ;
        RECT 2179.545 2590.610 2179.875 2590.625 ;
        RECT 2175.150 2590.310 2179.875 2590.610 ;
        RECT 2175.150 2590.300 2175.530 2590.310 ;
        RECT 2176.785 2590.295 2177.115 2590.310 ;
        RECT 2179.545 2590.295 2179.875 2590.310 ;
        RECT 2180.670 2590.610 2181.050 2590.620 ;
        RECT 2183.685 2590.610 2184.015 2590.625 ;
        RECT 2180.670 2590.310 2184.015 2590.610 ;
        RECT 2180.670 2590.300 2181.050 2590.310 ;
        RECT 2183.685 2590.295 2184.015 2590.310 ;
        RECT 1566.365 2589.930 1566.695 2589.945 ;
        RECT 1569.790 2589.930 1570.170 2589.940 ;
        RECT 1566.365 2589.630 1570.170 2589.930 ;
        RECT 1566.365 2589.615 1566.695 2589.630 ;
        RECT 1569.790 2589.620 1570.170 2589.630 ;
        RECT 1587.065 2589.930 1587.395 2589.945 ;
        RECT 1592.790 2589.930 1593.170 2589.940 ;
        RECT 1587.065 2589.630 1593.170 2589.930 ;
        RECT 1587.065 2589.615 1587.395 2589.630 ;
        RECT 1592.790 2589.620 1593.170 2589.630 ;
        RECT 1600.865 2589.930 1601.195 2589.945 ;
        RECT 1604.750 2589.930 1605.130 2589.940 ;
        RECT 1600.865 2589.630 1605.130 2589.930 ;
        RECT 1600.865 2589.615 1601.195 2589.630 ;
        RECT 1604.750 2589.620 1605.130 2589.630 ;
        RECT 1642.265 2589.930 1642.595 2589.945 ;
        RECT 1645.230 2589.930 1645.610 2589.940 ;
        RECT 1642.265 2589.630 1645.610 2589.930 ;
        RECT 1642.265 2589.615 1642.595 2589.630 ;
        RECT 1645.230 2589.620 1645.610 2589.630 ;
        RECT 1662.965 2589.930 1663.295 2589.945 ;
        RECT 2186.445 2589.940 2186.775 2589.945 ;
        RECT 1663.630 2589.930 1664.010 2589.940 ;
        RECT 1662.965 2589.630 1664.010 2589.930 ;
        RECT 1662.965 2589.615 1663.295 2589.630 ;
        RECT 1663.630 2589.620 1664.010 2589.630 ;
        RECT 2186.190 2589.930 2186.775 2589.940 ;
        RECT 2186.190 2589.630 2187.000 2589.930 ;
        RECT 2186.190 2589.620 2186.775 2589.630 ;
        RECT 2186.445 2589.615 2186.775 2589.620 ;
        RECT 1631.225 2589.250 1631.555 2589.265 ;
        RECT 1634.190 2589.250 1634.570 2589.260 ;
        RECT 1631.225 2588.950 1634.570 2589.250 ;
        RECT 1631.225 2588.935 1631.555 2588.950 ;
        RECT 1634.190 2588.940 1634.570 2588.950 ;
        RECT 1683.665 2589.250 1683.995 2589.265 ;
        RECT 1686.630 2589.250 1687.010 2589.260 ;
        RECT 1683.665 2588.950 1687.010 2589.250 ;
        RECT 1683.665 2588.935 1683.995 2588.950 ;
        RECT 1686.630 2588.940 1687.010 2588.950 ;
        RECT 1690.565 2589.250 1690.895 2589.265 ;
        RECT 1692.150 2589.250 1692.530 2589.260 ;
        RECT 1690.565 2588.950 1692.530 2589.250 ;
        RECT 1690.565 2588.935 1690.895 2588.950 ;
        RECT 1692.150 2588.940 1692.530 2588.950 ;
        RECT 2168.710 2589.250 2169.090 2589.260 ;
        RECT 2170.345 2589.250 2170.675 2589.265 ;
        RECT 2168.710 2588.950 2170.675 2589.250 ;
        RECT 2168.710 2588.940 2169.090 2588.950 ;
        RECT 2170.345 2588.935 2170.675 2588.950 ;
        RECT 1551.390 2588.570 1551.770 2588.580 ;
        RECT 1552.105 2588.570 1552.435 2588.585 ;
        RECT 1551.390 2588.270 1552.435 2588.570 ;
        RECT 1551.390 2588.260 1551.770 2588.270 ;
        RECT 1552.105 2588.255 1552.435 2588.270 ;
        RECT 1559.465 2588.570 1559.795 2588.585 ;
        RECT 1563.350 2588.570 1563.730 2588.580 ;
        RECT 1559.465 2588.270 1563.730 2588.570 ;
        RECT 1559.465 2588.255 1559.795 2588.270 ;
        RECT 1563.350 2588.260 1563.730 2588.270 ;
        RECT 1621.565 2588.570 1621.895 2588.585 ;
        RECT 1627.750 2588.570 1628.130 2588.580 ;
        RECT 1621.565 2588.270 1628.130 2588.570 ;
        RECT 1621.565 2588.255 1621.895 2588.270 ;
        RECT 1627.750 2588.260 1628.130 2588.270 ;
        RECT 1635.365 2588.570 1635.695 2588.585 ;
        RECT 1639.710 2588.570 1640.090 2588.580 ;
        RECT 1635.365 2588.270 1640.090 2588.570 ;
        RECT 1635.365 2588.255 1635.695 2588.270 ;
        RECT 1639.710 2588.260 1640.090 2588.270 ;
        RECT 1662.965 2588.570 1663.295 2588.585 ;
        RECT 1669.150 2588.570 1669.530 2588.580 ;
        RECT 1662.965 2588.270 1669.530 2588.570 ;
        RECT 1662.965 2588.255 1663.295 2588.270 ;
        RECT 1669.150 2588.260 1669.530 2588.270 ;
        RECT 1669.865 2588.570 1670.195 2588.585 ;
        RECT 1697.465 2588.580 1697.795 2588.585 ;
        RECT 1674.670 2588.570 1675.050 2588.580 ;
        RECT 1697.465 2588.570 1698.050 2588.580 ;
        RECT 1669.865 2588.270 1675.050 2588.570 ;
        RECT 1697.240 2588.270 1698.050 2588.570 ;
        RECT 1669.865 2588.255 1670.195 2588.270 ;
        RECT 1674.670 2588.260 1675.050 2588.270 ;
        RECT 1697.465 2588.260 1698.050 2588.270 ;
        RECT 1741.830 2588.570 1742.210 2588.580 ;
        RECT 1745.305 2588.570 1745.635 2588.585 ;
        RECT 2162.985 2588.580 2163.315 2588.585 ;
        RECT 2162.985 2588.570 2163.570 2588.580 ;
        RECT 1741.830 2588.270 1745.635 2588.570 ;
        RECT 2162.760 2588.270 2163.570 2588.570 ;
        RECT 1741.830 2588.260 1742.210 2588.270 ;
        RECT 1697.465 2588.255 1697.795 2588.260 ;
        RECT 1745.305 2588.255 1745.635 2588.270 ;
        RECT 2162.985 2588.260 2163.570 2588.270 ;
        RECT 2165.030 2588.570 2165.410 2588.580 ;
        RECT 2166.205 2588.570 2166.535 2588.585 ;
        RECT 2165.030 2588.270 2166.535 2588.570 ;
        RECT 2165.030 2588.260 2165.410 2588.270 ;
        RECT 2162.985 2588.255 2163.315 2588.260 ;
        RECT 2166.205 2588.255 2166.535 2588.270 ;
        RECT 2169.630 2588.570 2170.010 2588.580 ;
        RECT 2173.105 2588.570 2173.435 2588.585 ;
        RECT 2169.630 2588.270 2173.435 2588.570 ;
        RECT 2169.630 2588.260 2170.010 2588.270 ;
        RECT 2173.105 2588.255 2173.435 2588.270 ;
        RECT 2178.830 2588.570 2179.210 2588.580 ;
        RECT 2180.005 2588.570 2180.335 2588.585 ;
        RECT 2178.830 2588.270 2180.335 2588.570 ;
        RECT 2178.830 2588.260 2179.210 2588.270 ;
        RECT 2180.005 2588.255 2180.335 2588.270 ;
        RECT 2184.350 2588.570 2184.730 2588.580 ;
        RECT 2186.905 2588.570 2187.235 2588.585 ;
        RECT 2184.350 2588.270 2187.235 2588.570 ;
        RECT 2184.350 2588.260 2184.730 2588.270 ;
        RECT 2186.905 2588.255 2187.235 2588.270 ;
        RECT 2189.870 2588.570 2190.250 2588.580 ;
        RECT 2193.805 2588.570 2194.135 2588.585 ;
        RECT 2189.870 2588.270 2194.135 2588.570 ;
        RECT 2189.870 2588.260 2190.250 2588.270 ;
        RECT 2193.805 2588.255 2194.135 2588.270 ;
        RECT 2197.485 2588.570 2197.815 2588.585 ;
        RECT 2198.150 2588.570 2198.530 2588.580 ;
        RECT 2197.485 2588.270 2198.530 2588.570 ;
        RECT 2197.485 2588.255 2197.815 2588.270 ;
        RECT 2198.150 2588.260 2198.530 2588.270 ;
        RECT 2203.670 2588.570 2204.050 2588.580 ;
        RECT 2204.385 2588.570 2204.715 2588.585 ;
        RECT 2203.670 2588.270 2204.715 2588.570 ;
        RECT 2203.670 2588.260 2204.050 2588.270 ;
        RECT 2204.385 2588.255 2204.715 2588.270 ;
        RECT 2224.830 2588.570 2225.210 2588.580 ;
        RECT 2228.305 2588.570 2228.635 2588.585 ;
        RECT 2224.830 2588.270 2228.635 2588.570 ;
        RECT 2224.830 2588.260 2225.210 2588.270 ;
        RECT 2228.305 2588.255 2228.635 2588.270 ;
        RECT 2266.230 2588.570 2266.610 2588.580 ;
        RECT 2269.245 2588.570 2269.575 2588.585 ;
        RECT 2266.230 2588.270 2269.575 2588.570 ;
        RECT 2266.230 2588.260 2266.610 2588.270 ;
        RECT 2269.245 2588.255 2269.575 2588.270 ;
        RECT 2301.190 2588.570 2301.570 2588.580 ;
        RECT 2303.745 2588.570 2304.075 2588.585 ;
        RECT 2301.190 2588.270 2304.075 2588.570 ;
        RECT 2301.190 2588.260 2301.570 2588.270 ;
        RECT 2303.745 2588.255 2304.075 2588.270 ;
        RECT 2341.670 2588.570 2342.050 2588.580 ;
        RECT 2345.145 2588.570 2345.475 2588.585 ;
        RECT 2341.670 2588.270 2345.475 2588.570 ;
        RECT 2341.670 2588.260 2342.050 2588.270 ;
        RECT 2345.145 2588.255 2345.475 2588.270 ;
        RECT 1536.670 2587.890 1537.050 2587.900 ;
        RECT 1538.305 2587.890 1538.635 2587.905 ;
        RECT 1536.670 2587.590 1538.635 2587.890 ;
        RECT 1536.670 2587.580 1537.050 2587.590 ;
        RECT 1538.305 2587.575 1538.635 2587.590 ;
        RECT 1543.110 2587.890 1543.490 2587.900 ;
        RECT 1545.205 2587.890 1545.535 2587.905 ;
        RECT 1543.110 2587.590 1545.535 2587.890 ;
        RECT 1543.110 2587.580 1543.490 2587.590 ;
        RECT 1545.205 2587.575 1545.535 2587.590 ;
        RECT 1548.630 2587.890 1549.010 2587.900 ;
        RECT 1551.185 2587.890 1551.515 2587.905 ;
        RECT 1559.005 2587.900 1559.335 2587.905 ;
        RECT 1558.750 2587.890 1559.335 2587.900 ;
        RECT 1548.630 2587.590 1551.515 2587.890 ;
        RECT 1558.550 2587.590 1559.335 2587.890 ;
        RECT 1548.630 2587.580 1549.010 2587.590 ;
        RECT 1551.185 2587.575 1551.515 2587.590 ;
        RECT 1558.750 2587.580 1559.335 2587.590 ;
        RECT 1559.005 2587.575 1559.335 2587.580 ;
        RECT 1649.165 2587.890 1649.495 2587.905 ;
        RECT 1651.670 2587.890 1652.050 2587.900 ;
        RECT 1649.165 2587.590 1652.050 2587.890 ;
        RECT 1649.165 2587.575 1649.495 2587.590 ;
        RECT 1651.670 2587.580 1652.050 2587.590 ;
        RECT 1697.005 2587.890 1697.335 2587.905 ;
        RECT 1703.190 2587.890 1703.570 2587.900 ;
        RECT 1697.005 2587.590 1703.570 2587.890 ;
        RECT 1697.005 2587.575 1697.335 2587.590 ;
        RECT 1703.190 2587.580 1703.570 2587.590 ;
        RECT 1703.905 2587.890 1704.235 2587.905 ;
        RECT 1709.630 2587.890 1710.010 2587.900 ;
        RECT 1703.905 2587.590 1710.010 2587.890 ;
        RECT 1703.905 2587.575 1704.235 2587.590 ;
        RECT 1709.630 2587.580 1710.010 2587.590 ;
        RECT 1714.485 2587.890 1714.815 2587.905 ;
        RECT 1721.385 2587.900 1721.715 2587.905 ;
        RECT 1716.990 2587.890 1717.370 2587.900 ;
        RECT 1721.385 2587.890 1721.970 2587.900 ;
        RECT 1714.485 2587.590 1717.370 2587.890 ;
        RECT 1721.160 2587.590 1721.970 2587.890 ;
        RECT 1714.485 2587.575 1714.815 2587.590 ;
        RECT 1716.990 2587.580 1717.370 2587.590 ;
        RECT 1721.385 2587.580 1721.970 2587.590 ;
        RECT 1729.870 2587.890 1730.250 2587.900 ;
        RECT 1731.505 2587.890 1731.835 2587.905 ;
        RECT 1736.565 2587.900 1736.895 2587.905 ;
        RECT 1744.845 2587.900 1745.175 2587.905 ;
        RECT 1736.310 2587.890 1736.895 2587.900 ;
        RECT 1744.590 2587.890 1745.175 2587.900 ;
        RECT 1729.870 2587.590 1731.835 2587.890 ;
        RECT 1736.110 2587.590 1736.895 2587.890 ;
        RECT 1744.390 2587.590 1745.175 2587.890 ;
        RECT 1729.870 2587.580 1730.250 2587.590 ;
        RECT 1721.385 2587.575 1721.715 2587.580 ;
        RECT 1731.505 2587.575 1731.835 2587.590 ;
        RECT 1736.310 2587.580 1736.895 2587.590 ;
        RECT 1744.590 2587.580 1745.175 2587.590 ;
        RECT 1736.565 2587.575 1736.895 2587.580 ;
        RECT 1744.845 2587.575 1745.175 2587.580 ;
        RECT 2190.585 2587.890 2190.915 2587.905 ;
        RECT 2193.345 2587.900 2193.675 2587.905 ;
        RECT 2191.710 2587.890 2192.090 2587.900 ;
        RECT 2193.345 2587.890 2193.930 2587.900 ;
        RECT 2190.585 2587.590 2192.090 2587.890 ;
        RECT 2193.120 2587.590 2193.930 2587.890 ;
        RECT 2190.585 2587.575 2190.915 2587.590 ;
        RECT 2191.710 2587.580 2192.090 2587.590 ;
        RECT 2193.345 2587.580 2193.930 2587.590 ;
        RECT 2199.990 2587.890 2200.370 2587.900 ;
        RECT 2200.705 2587.890 2201.035 2587.905 ;
        RECT 2207.605 2587.900 2207.935 2587.905 ;
        RECT 2207.350 2587.890 2207.935 2587.900 ;
        RECT 2199.990 2587.590 2201.035 2587.890 ;
        RECT 2207.150 2587.590 2207.935 2587.890 ;
        RECT 2199.990 2587.580 2200.370 2587.590 ;
        RECT 2193.345 2587.575 2193.675 2587.580 ;
        RECT 2200.705 2587.575 2201.035 2587.590 ;
        RECT 2207.350 2587.580 2207.935 2587.590 ;
        RECT 2213.790 2587.890 2214.170 2587.900 ;
        RECT 2214.505 2587.890 2214.835 2587.905 ;
        RECT 2213.790 2587.590 2214.835 2587.890 ;
        RECT 2213.790 2587.580 2214.170 2587.590 ;
        RECT 2207.605 2587.575 2207.935 2587.580 ;
        RECT 2214.505 2587.575 2214.835 2587.590 ;
        RECT 2219.310 2587.890 2219.690 2587.900 ;
        RECT 2221.405 2587.890 2221.735 2587.905 ;
        RECT 2227.845 2587.900 2228.175 2587.905 ;
        RECT 2235.205 2587.900 2235.535 2587.905 ;
        RECT 2227.590 2587.890 2228.175 2587.900 ;
        RECT 2234.950 2587.890 2235.535 2587.900 ;
        RECT 2219.310 2587.590 2221.735 2587.890 ;
        RECT 2227.390 2587.590 2228.175 2587.890 ;
        RECT 2234.750 2587.590 2235.535 2587.890 ;
        RECT 2219.310 2587.580 2219.690 2587.590 ;
        RECT 2221.405 2587.575 2221.735 2587.590 ;
        RECT 2227.590 2587.580 2228.175 2587.590 ;
        RECT 2234.950 2587.580 2235.535 2587.590 ;
        RECT 2241.390 2587.890 2241.770 2587.900 ;
        RECT 2242.105 2587.890 2242.435 2587.905 ;
        RECT 2249.005 2587.900 2249.335 2587.905 ;
        RECT 2248.750 2587.890 2249.335 2587.900 ;
        RECT 2241.390 2587.590 2242.435 2587.890 ;
        RECT 2248.550 2587.590 2249.335 2587.890 ;
        RECT 2241.390 2587.580 2241.770 2587.590 ;
        RECT 2227.845 2587.575 2228.175 2587.580 ;
        RECT 2235.205 2587.575 2235.535 2587.580 ;
        RECT 2242.105 2587.575 2242.435 2587.590 ;
        RECT 2248.750 2587.580 2249.335 2587.590 ;
        RECT 2254.270 2587.890 2254.650 2587.900 ;
        RECT 2255.905 2587.890 2256.235 2587.905 ;
        RECT 2254.270 2587.590 2256.235 2587.890 ;
        RECT 2254.270 2587.580 2254.650 2587.590 ;
        RECT 2249.005 2587.575 2249.335 2587.580 ;
        RECT 2255.905 2587.575 2256.235 2587.590 ;
        RECT 2259.790 2587.890 2260.170 2587.900 ;
        RECT 2262.805 2587.890 2263.135 2587.905 ;
        RECT 2259.790 2587.590 2263.135 2587.890 ;
        RECT 2259.790 2587.580 2260.170 2587.590 ;
        RECT 2262.805 2587.575 2263.135 2587.590 ;
        RECT 2268.990 2587.890 2269.370 2587.900 ;
        RECT 2269.705 2587.890 2270.035 2587.905 ;
        RECT 2276.605 2587.900 2276.935 2587.905 ;
        RECT 2276.350 2587.890 2276.935 2587.900 ;
        RECT 2268.990 2587.590 2270.035 2587.890 ;
        RECT 2276.150 2587.590 2276.935 2587.890 ;
        RECT 2268.990 2587.580 2269.370 2587.590 ;
        RECT 2269.705 2587.575 2270.035 2587.590 ;
        RECT 2276.350 2587.580 2276.935 2587.590 ;
        RECT 2281.870 2587.890 2282.250 2587.900 ;
        RECT 2283.505 2587.890 2283.835 2587.905 ;
        RECT 2281.870 2587.590 2283.835 2587.890 ;
        RECT 2281.870 2587.580 2282.250 2587.590 ;
        RECT 2276.605 2587.575 2276.935 2587.580 ;
        RECT 2283.505 2587.575 2283.835 2587.590 ;
        RECT 2289.230 2587.890 2289.610 2587.900 ;
        RECT 2290.405 2587.890 2290.735 2587.905 ;
        RECT 2289.230 2587.590 2290.735 2587.890 ;
        RECT 2289.230 2587.580 2289.610 2587.590 ;
        RECT 2290.405 2587.575 2290.735 2587.590 ;
        RECT 2295.670 2587.890 2296.050 2587.900 ;
        RECT 2297.305 2587.890 2297.635 2587.905 ;
        RECT 2304.205 2587.900 2304.535 2587.905 ;
        RECT 2303.950 2587.890 2304.535 2587.900 ;
        RECT 2295.670 2587.590 2297.635 2587.890 ;
        RECT 2303.750 2587.590 2304.535 2587.890 ;
        RECT 2295.670 2587.580 2296.050 2587.590 ;
        RECT 2297.305 2587.575 2297.635 2587.590 ;
        RECT 2303.950 2587.580 2304.535 2587.590 ;
        RECT 2310.390 2587.890 2310.770 2587.900 ;
        RECT 2311.105 2587.890 2311.435 2587.905 ;
        RECT 2318.005 2587.900 2318.335 2587.905 ;
        RECT 2317.750 2587.890 2318.335 2587.900 ;
        RECT 2310.390 2587.590 2311.435 2587.890 ;
        RECT 2317.550 2587.590 2318.335 2587.890 ;
        RECT 2310.390 2587.580 2310.770 2587.590 ;
        RECT 2304.205 2587.575 2304.535 2587.580 ;
        RECT 2311.105 2587.575 2311.435 2587.590 ;
        RECT 2317.750 2587.580 2318.335 2587.590 ;
        RECT 2324.190 2587.890 2324.570 2587.900 ;
        RECT 2324.905 2587.890 2325.235 2587.905 ;
        RECT 2324.190 2587.590 2325.235 2587.890 ;
        RECT 2324.190 2587.580 2324.570 2587.590 ;
        RECT 2318.005 2587.575 2318.335 2587.580 ;
        RECT 2324.905 2587.575 2325.235 2587.590 ;
        RECT 2330.630 2587.890 2331.010 2587.900 ;
        RECT 2331.805 2587.890 2332.135 2587.905 ;
        RECT 2330.630 2587.590 2332.135 2587.890 ;
        RECT 2330.630 2587.580 2331.010 2587.590 ;
        RECT 2331.805 2587.575 2332.135 2587.590 ;
        RECT 2336.150 2587.890 2336.530 2587.900 ;
        RECT 2338.705 2587.890 2339.035 2587.905 ;
        RECT 2345.605 2587.900 2345.935 2587.905 ;
        RECT 2345.350 2587.890 2345.935 2587.900 ;
        RECT 2336.150 2587.590 2339.035 2587.890 ;
        RECT 2345.150 2587.590 2345.935 2587.890 ;
        RECT 2336.150 2587.580 2336.530 2587.590 ;
        RECT 2338.705 2587.575 2339.035 2587.590 ;
        RECT 2345.350 2587.580 2345.935 2587.590 ;
        RECT 2345.605 2587.575 2345.935 2587.580 ;
        RECT 2168.965 2560.010 2169.295 2560.025 ;
        RECT 2169.885 2560.010 2170.215 2560.025 ;
        RECT 2168.965 2559.710 2170.215 2560.010 ;
        RECT 2168.965 2559.695 2169.295 2559.710 ;
        RECT 2169.885 2559.695 2170.215 2559.710 ;
        RECT 2168.045 2415.170 2168.375 2415.185 ;
        RECT 2168.965 2415.170 2169.295 2415.185 ;
        RECT 2168.045 2414.870 2169.295 2415.170 ;
        RECT 2168.045 2414.855 2168.375 2414.870 ;
        RECT 2168.965 2414.855 2169.295 2414.870 ;
        RECT 1835.925 2412.450 1836.255 2412.465 ;
        RECT 1877.325 2412.450 1877.655 2412.465 ;
        RECT 1835.925 2412.150 1877.655 2412.450 ;
        RECT 1835.925 2412.135 1836.255 2412.150 ;
        RECT 1877.325 2412.135 1877.655 2412.150 ;
        RECT 2338.705 2412.450 2339.035 2412.465 ;
        RECT 2559.965 2412.450 2560.295 2412.465 ;
        RECT 2338.705 2412.150 2560.295 2412.450 ;
        RECT 2338.705 2412.135 2339.035 2412.150 ;
        RECT 2559.965 2412.135 2560.295 2412.150 ;
        RECT 1490.005 2411.770 1490.335 2411.785 ;
        RECT 1942.645 2411.770 1942.975 2411.785 ;
        RECT 1490.005 2411.470 1942.975 2411.770 ;
        RECT 1490.005 2411.455 1490.335 2411.470 ;
        RECT 1942.645 2411.455 1942.975 2411.470 ;
        RECT 2345.605 2411.770 2345.935 2411.785 ;
        RECT 2581.585 2411.770 2581.915 2411.785 ;
        RECT 2345.605 2411.470 2581.915 2411.770 ;
        RECT 2345.605 2411.455 2345.935 2411.470 ;
        RECT 2581.585 2411.455 2581.915 2411.470 ;
        RECT 1417.325 2411.090 1417.655 2411.105 ;
        RECT 1898.485 2411.090 1898.815 2411.105 ;
        RECT 1417.325 2410.790 1898.815 2411.090 ;
        RECT 1417.325 2410.775 1417.655 2410.790 ;
        RECT 1898.485 2410.775 1898.815 2410.790 ;
        RECT 1932.525 2411.090 1932.855 2411.105 ;
        RECT 1945.865 2411.090 1946.195 2411.105 ;
        RECT 1932.525 2410.790 1946.195 2411.090 ;
        RECT 1932.525 2410.775 1932.855 2410.790 ;
        RECT 1945.865 2410.775 1946.195 2410.790 ;
        RECT 2090.305 2411.090 2090.635 2411.105 ;
        RECT 2592.625 2411.090 2592.955 2411.105 ;
        RECT 2090.305 2410.790 2592.955 2411.090 ;
        RECT 2090.305 2410.775 2090.635 2410.790 ;
        RECT 2592.625 2410.775 2592.955 2410.790 ;
        RECT 1593.965 2410.410 1594.295 2410.425 ;
        RECT 1609.605 2410.410 1609.935 2410.425 ;
        RECT 1593.965 2410.110 1609.935 2410.410 ;
        RECT 1593.965 2410.095 1594.295 2410.110 ;
        RECT 1609.605 2410.095 1609.935 2410.110 ;
      LAYER met3 ;
        RECT 1403.990 2395.120 2596.000 2395.945 ;
        RECT 1404.400 2393.720 2595.600 2395.120 ;
        RECT 1403.990 2384.920 2596.000 2393.720 ;
        RECT 1403.990 2384.240 2595.600 2384.920 ;
        RECT 1404.400 2383.520 2595.600 2384.240 ;
        RECT 1404.400 2382.840 2596.000 2383.520 ;
        RECT 1403.990 2374.040 2596.000 2382.840 ;
        RECT 1404.400 2372.640 2595.600 2374.040 ;
        RECT 1403.990 2363.840 2596.000 2372.640 ;
        RECT 1403.990 2363.160 2595.600 2363.840 ;
        RECT 1404.400 2362.440 2595.600 2363.160 ;
        RECT 1404.400 2361.760 2596.000 2362.440 ;
        RECT 1403.990 2352.960 2596.000 2361.760 ;
        RECT 1403.990 2352.280 2595.600 2352.960 ;
        RECT 1404.400 2351.560 2595.600 2352.280 ;
        RECT 1404.400 2350.880 2596.000 2351.560 ;
        RECT 1403.990 2342.760 2596.000 2350.880 ;
        RECT 1403.990 2342.080 2595.600 2342.760 ;
        RECT 1404.400 2341.360 2595.600 2342.080 ;
        RECT 1404.400 2340.680 2596.000 2341.360 ;
        RECT 1403.990 2331.880 2596.000 2340.680 ;
        RECT 1403.990 2331.200 2595.600 2331.880 ;
        RECT 1404.400 2330.480 2595.600 2331.200 ;
        RECT 1404.400 2329.800 2596.000 2330.480 ;
        RECT 1403.990 2321.680 2596.000 2329.800 ;
        RECT 1403.990 2321.000 2595.600 2321.680 ;
        RECT 1404.400 2320.280 2595.600 2321.000 ;
        RECT 1404.400 2319.600 2596.000 2320.280 ;
        RECT 1403.990 2310.800 2596.000 2319.600 ;
        RECT 1403.990 2310.120 2595.600 2310.800 ;
        RECT 1404.400 2309.400 2595.600 2310.120 ;
        RECT 1404.400 2308.720 2596.000 2309.400 ;
        RECT 1403.990 2300.600 2596.000 2308.720 ;
        RECT 1403.990 2299.240 2595.600 2300.600 ;
        RECT 1404.400 2299.200 2595.600 2299.240 ;
        RECT 1404.400 2297.840 2596.000 2299.200 ;
        RECT 1403.990 2289.720 2596.000 2297.840 ;
        RECT 1403.990 2289.040 2595.600 2289.720 ;
        RECT 1404.400 2288.320 2595.600 2289.040 ;
        RECT 1404.400 2287.640 2596.000 2288.320 ;
        RECT 1403.990 2279.520 2596.000 2287.640 ;
        RECT 1403.990 2278.160 2595.600 2279.520 ;
        RECT 1404.400 2278.120 2595.600 2278.160 ;
        RECT 1404.400 2276.760 2596.000 2278.120 ;
        RECT 1403.990 2268.640 2596.000 2276.760 ;
        RECT 1403.990 2267.280 2595.600 2268.640 ;
        RECT 1404.400 2267.240 2595.600 2267.280 ;
        RECT 1404.400 2265.880 2596.000 2267.240 ;
        RECT 1403.990 2258.440 2596.000 2265.880 ;
        RECT 1403.990 2257.080 2595.600 2258.440 ;
        RECT 1404.400 2257.040 2595.600 2257.080 ;
        RECT 1404.400 2255.680 2596.000 2257.040 ;
        RECT 1403.990 2247.560 2596.000 2255.680 ;
        RECT 1403.990 2246.200 2595.600 2247.560 ;
        RECT 1404.400 2246.160 2595.600 2246.200 ;
        RECT 1404.400 2244.800 2596.000 2246.160 ;
        RECT 1403.990 2237.360 2596.000 2244.800 ;
        RECT 1403.990 2236.000 2595.600 2237.360 ;
        RECT 1404.400 2235.960 2595.600 2236.000 ;
        RECT 1404.400 2234.600 2596.000 2235.960 ;
        RECT 1403.990 2226.480 2596.000 2234.600 ;
        RECT 1403.990 2225.120 2595.600 2226.480 ;
        RECT 1404.400 2225.080 2595.600 2225.120 ;
        RECT 1404.400 2223.720 2596.000 2225.080 ;
        RECT 1403.990 2216.280 2596.000 2223.720 ;
        RECT 1403.990 2214.880 2595.600 2216.280 ;
        RECT 1403.990 2214.240 2596.000 2214.880 ;
        RECT 1404.400 2212.840 2596.000 2214.240 ;
        RECT 1403.990 2205.400 2596.000 2212.840 ;
        RECT 1403.990 2204.040 2595.600 2205.400 ;
        RECT 1404.400 2204.000 2595.600 2204.040 ;
        RECT 1404.400 2202.640 2596.000 2204.000 ;
        RECT 1403.990 2195.200 2596.000 2202.640 ;
        RECT 1403.990 2193.800 2595.600 2195.200 ;
        RECT 1403.990 2193.160 2596.000 2193.800 ;
        RECT 1404.400 2191.760 2596.000 2193.160 ;
        RECT 1403.990 2184.320 2596.000 2191.760 ;
        RECT 1403.990 2182.920 2595.600 2184.320 ;
        RECT 1403.990 2182.280 2596.000 2182.920 ;
        RECT 1404.400 2180.880 2596.000 2182.280 ;
        RECT 1403.990 2174.120 2596.000 2180.880 ;
        RECT 1403.990 2172.720 2595.600 2174.120 ;
        RECT 1403.990 2172.080 2596.000 2172.720 ;
        RECT 1404.400 2170.680 2596.000 2172.080 ;
        RECT 1403.990 2163.240 2596.000 2170.680 ;
        RECT 1403.990 2161.840 2595.600 2163.240 ;
        RECT 1403.990 2161.200 2596.000 2161.840 ;
        RECT 1404.400 2159.800 2596.000 2161.200 ;
        RECT 1403.990 2153.040 2596.000 2159.800 ;
        RECT 1403.990 2151.640 2595.600 2153.040 ;
        RECT 1403.990 2151.000 2596.000 2151.640 ;
        RECT 1404.400 2149.600 2596.000 2151.000 ;
        RECT 1403.990 2142.160 2596.000 2149.600 ;
        RECT 1403.990 2140.760 2595.600 2142.160 ;
        RECT 1403.990 2140.120 2596.000 2140.760 ;
        RECT 1404.400 2138.720 2596.000 2140.120 ;
        RECT 1403.990 2131.960 2596.000 2138.720 ;
        RECT 1403.990 2130.560 2595.600 2131.960 ;
        RECT 1403.990 2129.240 2596.000 2130.560 ;
        RECT 1404.400 2127.840 2596.000 2129.240 ;
        RECT 1403.990 2121.080 2596.000 2127.840 ;
        RECT 1403.990 2119.680 2595.600 2121.080 ;
        RECT 1403.990 2119.040 2596.000 2119.680 ;
        RECT 1404.400 2117.640 2596.000 2119.040 ;
        RECT 1403.990 2110.880 2596.000 2117.640 ;
        RECT 1403.990 2109.480 2595.600 2110.880 ;
        RECT 1403.990 2108.160 2596.000 2109.480 ;
        RECT 1404.400 2106.760 2596.000 2108.160 ;
        RECT 1403.990 2100.680 2596.000 2106.760 ;
        RECT 1403.990 2099.280 2595.600 2100.680 ;
        RECT 1403.990 2097.960 2596.000 2099.280 ;
        RECT 1404.400 2096.560 2596.000 2097.960 ;
        RECT 1403.990 2089.800 2596.000 2096.560 ;
        RECT 1403.990 2088.400 2595.600 2089.800 ;
        RECT 1403.990 2087.080 2596.000 2088.400 ;
        RECT 1404.400 2085.680 2596.000 2087.080 ;
        RECT 1403.990 2079.600 2596.000 2085.680 ;
        RECT 1403.990 2078.200 2595.600 2079.600 ;
        RECT 1403.990 2076.200 2596.000 2078.200 ;
        RECT 1404.400 2074.800 2596.000 2076.200 ;
        RECT 1403.990 2068.720 2596.000 2074.800 ;
        RECT 1403.990 2067.320 2595.600 2068.720 ;
        RECT 1403.990 2066.000 2596.000 2067.320 ;
        RECT 1404.400 2064.600 2596.000 2066.000 ;
        RECT 1403.990 2058.520 2596.000 2064.600 ;
        RECT 1403.990 2057.120 2595.600 2058.520 ;
        RECT 1403.990 2055.120 2596.000 2057.120 ;
        RECT 1404.400 2053.720 2596.000 2055.120 ;
        RECT 1403.990 2047.640 2596.000 2053.720 ;
        RECT 1403.990 2046.240 2595.600 2047.640 ;
        RECT 1403.990 2044.240 2596.000 2046.240 ;
        RECT 1404.400 2042.840 2596.000 2044.240 ;
        RECT 1403.990 2037.440 2596.000 2042.840 ;
        RECT 1403.990 2036.040 2595.600 2037.440 ;
        RECT 1403.990 2034.040 2596.000 2036.040 ;
        RECT 1404.400 2032.640 2596.000 2034.040 ;
        RECT 1403.990 2026.560 2596.000 2032.640 ;
        RECT 1403.990 2025.160 2595.600 2026.560 ;
        RECT 1403.990 2023.160 2596.000 2025.160 ;
        RECT 1404.400 2021.760 2596.000 2023.160 ;
        RECT 1403.990 2016.360 2596.000 2021.760 ;
        RECT 1403.990 2014.960 2595.600 2016.360 ;
        RECT 1403.990 2012.960 2596.000 2014.960 ;
        RECT 1404.400 2011.560 2596.000 2012.960 ;
        RECT 1403.990 2005.480 2596.000 2011.560 ;
        RECT 1403.990 2004.080 2595.600 2005.480 ;
        RECT 1403.990 2002.080 2596.000 2004.080 ;
        RECT 1404.400 2000.680 2596.000 2002.080 ;
        RECT 1403.990 1995.280 2596.000 2000.680 ;
        RECT 1403.990 1993.880 2595.600 1995.280 ;
        RECT 1403.990 1991.200 2596.000 1993.880 ;
        RECT 1404.400 1989.800 2596.000 1991.200 ;
        RECT 1403.990 1984.400 2596.000 1989.800 ;
        RECT 1403.990 1983.000 2595.600 1984.400 ;
        RECT 1403.990 1981.000 2596.000 1983.000 ;
        RECT 1404.400 1979.600 2596.000 1981.000 ;
        RECT 1403.990 1974.200 2596.000 1979.600 ;
        RECT 1403.990 1972.800 2595.600 1974.200 ;
        RECT 1403.990 1970.120 2596.000 1972.800 ;
        RECT 1404.400 1968.720 2596.000 1970.120 ;
        RECT 1403.990 1963.320 2596.000 1968.720 ;
        RECT 1403.990 1961.920 2595.600 1963.320 ;
        RECT 1403.990 1959.240 2596.000 1961.920 ;
        RECT 1404.400 1957.840 2596.000 1959.240 ;
        RECT 1403.990 1953.120 2596.000 1957.840 ;
        RECT 1403.990 1951.720 2595.600 1953.120 ;
        RECT 1403.990 1949.040 2596.000 1951.720 ;
        RECT 1404.400 1947.640 2596.000 1949.040 ;
        RECT 1403.990 1942.240 2596.000 1947.640 ;
        RECT 1403.990 1940.840 2595.600 1942.240 ;
        RECT 1403.990 1938.160 2596.000 1940.840 ;
        RECT 1404.400 1936.760 2596.000 1938.160 ;
        RECT 1403.990 1932.040 2596.000 1936.760 ;
        RECT 1403.990 1930.640 2595.600 1932.040 ;
        RECT 1403.990 1927.960 2596.000 1930.640 ;
        RECT 1404.400 1926.560 2596.000 1927.960 ;
        RECT 1403.990 1921.160 2596.000 1926.560 ;
        RECT 1403.990 1919.760 2595.600 1921.160 ;
        RECT 1403.990 1917.080 2596.000 1919.760 ;
        RECT 1404.400 1915.680 2596.000 1917.080 ;
        RECT 1403.990 1910.960 2596.000 1915.680 ;
        RECT 1403.990 1909.560 2595.600 1910.960 ;
        RECT 1403.990 1906.200 2596.000 1909.560 ;
        RECT 1404.400 1904.800 2596.000 1906.200 ;
        RECT 1403.990 1900.080 2596.000 1904.800 ;
        RECT 1403.990 1898.680 2595.600 1900.080 ;
        RECT 1403.990 1896.000 2596.000 1898.680 ;
        RECT 1404.400 1894.600 2596.000 1896.000 ;
        RECT 1403.990 1889.880 2596.000 1894.600 ;
        RECT 1403.990 1888.480 2595.600 1889.880 ;
        RECT 1403.990 1885.120 2596.000 1888.480 ;
        RECT 1404.400 1883.720 2596.000 1885.120 ;
        RECT 1403.990 1879.000 2596.000 1883.720 ;
        RECT 1403.990 1877.600 2595.600 1879.000 ;
        RECT 1403.990 1874.920 2596.000 1877.600 ;
        RECT 1404.400 1873.520 2596.000 1874.920 ;
        RECT 1403.990 1868.800 2596.000 1873.520 ;
        RECT 1403.990 1867.400 2595.600 1868.800 ;
        RECT 1403.990 1864.040 2596.000 1867.400 ;
        RECT 1404.400 1862.640 2596.000 1864.040 ;
        RECT 1403.990 1857.920 2596.000 1862.640 ;
        RECT 1403.990 1856.520 2595.600 1857.920 ;
        RECT 1403.990 1853.160 2596.000 1856.520 ;
        RECT 1404.400 1851.760 2596.000 1853.160 ;
        RECT 1403.990 1847.720 2596.000 1851.760 ;
        RECT 1403.990 1846.320 2595.600 1847.720 ;
        RECT 1403.990 1842.960 2596.000 1846.320 ;
        RECT 1404.400 1841.560 2596.000 1842.960 ;
        RECT 1403.990 1836.840 2596.000 1841.560 ;
        RECT 1403.990 1835.440 2595.600 1836.840 ;
        RECT 1403.990 1832.080 2596.000 1835.440 ;
        RECT 1404.400 1830.680 2596.000 1832.080 ;
        RECT 1403.990 1826.640 2596.000 1830.680 ;
        RECT 1403.990 1825.240 2595.600 1826.640 ;
        RECT 1403.990 1821.200 2596.000 1825.240 ;
        RECT 1404.400 1819.800 2596.000 1821.200 ;
        RECT 1403.990 1815.760 2596.000 1819.800 ;
        RECT 1403.990 1814.360 2595.600 1815.760 ;
        RECT 1403.990 1811.000 2596.000 1814.360 ;
        RECT 1404.400 1809.600 2596.000 1811.000 ;
        RECT 1403.990 1805.560 2596.000 1809.600 ;
        RECT 1403.990 1804.160 2595.600 1805.560 ;
        RECT 1403.990 1800.120 2596.000 1804.160 ;
        RECT 1404.400 1798.720 2596.000 1800.120 ;
        RECT 1403.990 1795.360 2596.000 1798.720 ;
        RECT 1403.990 1793.960 2595.600 1795.360 ;
        RECT 1403.990 1789.920 2596.000 1793.960 ;
        RECT 1404.400 1788.520 2596.000 1789.920 ;
        RECT 1403.990 1784.480 2596.000 1788.520 ;
        RECT 1403.990 1783.080 2595.600 1784.480 ;
        RECT 1403.990 1779.040 2596.000 1783.080 ;
        RECT 1404.400 1777.640 2596.000 1779.040 ;
        RECT 1403.990 1774.280 2596.000 1777.640 ;
        RECT 1403.990 1772.880 2595.600 1774.280 ;
        RECT 1403.990 1768.160 2596.000 1772.880 ;
        RECT 1404.400 1766.760 2596.000 1768.160 ;
        RECT 1403.990 1763.400 2596.000 1766.760 ;
        RECT 1403.990 1762.000 2595.600 1763.400 ;
        RECT 1403.990 1757.960 2596.000 1762.000 ;
        RECT 1404.400 1756.560 2596.000 1757.960 ;
        RECT 1403.990 1753.200 2596.000 1756.560 ;
        RECT 1403.990 1751.800 2595.600 1753.200 ;
        RECT 1403.990 1747.080 2596.000 1751.800 ;
        RECT 1404.400 1745.680 2596.000 1747.080 ;
        RECT 1403.990 1742.320 2596.000 1745.680 ;
        RECT 1403.990 1740.920 2595.600 1742.320 ;
        RECT 1403.990 1736.200 2596.000 1740.920 ;
        RECT 1404.400 1734.800 2596.000 1736.200 ;
        RECT 1403.990 1732.120 2596.000 1734.800 ;
        RECT 1403.990 1730.720 2595.600 1732.120 ;
        RECT 1403.990 1726.000 2596.000 1730.720 ;
        RECT 1404.400 1724.600 2596.000 1726.000 ;
        RECT 1403.990 1721.240 2596.000 1724.600 ;
        RECT 1403.990 1719.840 2595.600 1721.240 ;
        RECT 1403.990 1715.120 2596.000 1719.840 ;
        RECT 1404.400 1713.720 2596.000 1715.120 ;
        RECT 1403.990 1711.040 2596.000 1713.720 ;
        RECT 1403.990 1709.640 2595.600 1711.040 ;
        RECT 1403.990 1704.920 2596.000 1709.640 ;
        RECT 1404.400 1703.520 2596.000 1704.920 ;
        RECT 1403.990 1700.160 2596.000 1703.520 ;
        RECT 1403.990 1698.760 2595.600 1700.160 ;
        RECT 1403.990 1694.040 2596.000 1698.760 ;
        RECT 1404.400 1692.640 2596.000 1694.040 ;
        RECT 1403.990 1689.960 2596.000 1692.640 ;
        RECT 1403.990 1688.560 2595.600 1689.960 ;
        RECT 1403.990 1683.160 2596.000 1688.560 ;
        RECT 1404.400 1681.760 2596.000 1683.160 ;
        RECT 1403.990 1679.080 2596.000 1681.760 ;
        RECT 1403.990 1677.680 2595.600 1679.080 ;
        RECT 1403.990 1672.960 2596.000 1677.680 ;
        RECT 1404.400 1671.560 2596.000 1672.960 ;
        RECT 1403.990 1668.880 2596.000 1671.560 ;
        RECT 1403.990 1667.480 2595.600 1668.880 ;
        RECT 1403.990 1662.080 2596.000 1667.480 ;
        RECT 1404.400 1660.680 2596.000 1662.080 ;
        RECT 1403.990 1658.000 2596.000 1660.680 ;
        RECT 1403.990 1656.600 2595.600 1658.000 ;
        RECT 1403.990 1651.880 2596.000 1656.600 ;
        RECT 1404.400 1650.480 2596.000 1651.880 ;
        RECT 1403.990 1647.800 2596.000 1650.480 ;
        RECT 1403.990 1646.400 2595.600 1647.800 ;
        RECT 1403.990 1641.000 2596.000 1646.400 ;
        RECT 1404.400 1639.600 2596.000 1641.000 ;
        RECT 1403.990 1636.920 2596.000 1639.600 ;
        RECT 1403.990 1635.520 2595.600 1636.920 ;
        RECT 1403.990 1630.120 2596.000 1635.520 ;
        RECT 1404.400 1628.720 2596.000 1630.120 ;
        RECT 1403.990 1626.720 2596.000 1628.720 ;
        RECT 1403.990 1625.320 2595.600 1626.720 ;
        RECT 1403.990 1619.920 2596.000 1625.320 ;
        RECT 1404.400 1618.520 2596.000 1619.920 ;
        RECT 1403.990 1615.840 2596.000 1618.520 ;
        RECT 1403.990 1614.440 2595.600 1615.840 ;
        RECT 1403.990 1609.040 2596.000 1614.440 ;
        RECT 1404.400 1607.640 2596.000 1609.040 ;
        RECT 1403.990 1605.640 2596.000 1607.640 ;
        RECT 1403.990 1604.240 2595.600 1605.640 ;
        RECT 1403.990 1598.160 2596.000 1604.240 ;
        RECT 1404.400 1596.760 2596.000 1598.160 ;
        RECT 1403.990 1594.760 2596.000 1596.760 ;
        RECT 1403.990 1593.360 2595.600 1594.760 ;
        RECT 1403.990 1587.960 2596.000 1593.360 ;
        RECT 1404.400 1586.560 2596.000 1587.960 ;
        RECT 1403.990 1584.560 2596.000 1586.560 ;
        RECT 1403.990 1583.160 2595.600 1584.560 ;
        RECT 1403.990 1577.080 2596.000 1583.160 ;
        RECT 1404.400 1575.680 2596.000 1577.080 ;
        RECT 1403.990 1573.680 2596.000 1575.680 ;
        RECT 1403.990 1572.280 2595.600 1573.680 ;
        RECT 1403.990 1566.880 2596.000 1572.280 ;
        RECT 1404.400 1565.480 2596.000 1566.880 ;
        RECT 1403.990 1563.480 2596.000 1565.480 ;
        RECT 1403.990 1562.080 2595.600 1563.480 ;
        RECT 1403.990 1556.000 2596.000 1562.080 ;
        RECT 1404.400 1554.600 2596.000 1556.000 ;
        RECT 1403.990 1552.600 2596.000 1554.600 ;
        RECT 1403.990 1551.200 2595.600 1552.600 ;
        RECT 1403.990 1545.120 2596.000 1551.200 ;
        RECT 1404.400 1543.720 2596.000 1545.120 ;
        RECT 1403.990 1542.400 2596.000 1543.720 ;
        RECT 1403.990 1541.000 2595.600 1542.400 ;
        RECT 1403.990 1534.920 2596.000 1541.000 ;
        RECT 1404.400 1533.520 2596.000 1534.920 ;
        RECT 1403.990 1531.520 2596.000 1533.520 ;
        RECT 1403.990 1530.120 2595.600 1531.520 ;
        RECT 1403.990 1524.040 2596.000 1530.120 ;
        RECT 1404.400 1522.640 2596.000 1524.040 ;
        RECT 1403.990 1521.320 2596.000 1522.640 ;
        RECT 1403.990 1519.920 2595.600 1521.320 ;
        RECT 1403.990 1513.160 2596.000 1519.920 ;
        RECT 1404.400 1511.760 2596.000 1513.160 ;
        RECT 1403.990 1510.440 2596.000 1511.760 ;
        RECT 1403.990 1509.040 2595.600 1510.440 ;
        RECT 1403.990 1502.960 2596.000 1509.040 ;
        RECT 1404.400 1501.560 2596.000 1502.960 ;
        RECT 1403.990 1500.240 2596.000 1501.560 ;
        RECT 1403.990 1498.840 2595.600 1500.240 ;
        RECT 1403.990 1492.080 2596.000 1498.840 ;
        RECT 1404.400 1490.680 2596.000 1492.080 ;
        RECT 1403.990 1490.040 2596.000 1490.680 ;
        RECT 1403.990 1488.640 2595.600 1490.040 ;
        RECT 1403.990 1481.880 2596.000 1488.640 ;
        RECT 1404.400 1480.480 2596.000 1481.880 ;
        RECT 1403.990 1479.160 2596.000 1480.480 ;
        RECT 1403.990 1477.760 2595.600 1479.160 ;
        RECT 1403.990 1471.000 2596.000 1477.760 ;
        RECT 1404.400 1469.600 2596.000 1471.000 ;
        RECT 1403.990 1468.960 2596.000 1469.600 ;
        RECT 1403.990 1467.560 2595.600 1468.960 ;
        RECT 1403.990 1460.120 2596.000 1467.560 ;
        RECT 1404.400 1458.720 2596.000 1460.120 ;
        RECT 1403.990 1458.080 2596.000 1458.720 ;
        RECT 1403.990 1456.680 2595.600 1458.080 ;
        RECT 1403.990 1449.920 2596.000 1456.680 ;
        RECT 1404.400 1448.520 2596.000 1449.920 ;
        RECT 1403.990 1447.880 2596.000 1448.520 ;
        RECT 1403.990 1446.480 2595.600 1447.880 ;
        RECT 1403.990 1439.040 2596.000 1446.480 ;
        RECT 1404.400 1437.640 2596.000 1439.040 ;
        RECT 1403.990 1437.000 2596.000 1437.640 ;
        RECT 1403.990 1435.600 2595.600 1437.000 ;
        RECT 1403.990 1428.840 2596.000 1435.600 ;
        RECT 1404.400 1427.440 2596.000 1428.840 ;
        RECT 1403.990 1426.800 2596.000 1427.440 ;
        RECT 1403.990 1425.400 2595.600 1426.800 ;
        RECT 1403.990 1417.960 2596.000 1425.400 ;
        RECT 1404.400 1416.560 2596.000 1417.960 ;
        RECT 1403.990 1415.920 2596.000 1416.560 ;
        RECT 1403.990 1414.520 2595.600 1415.920 ;
        RECT 1403.990 1407.080 2596.000 1414.520 ;
        RECT 1404.400 1405.720 2596.000 1407.080 ;
        RECT 1404.400 1405.680 2595.600 1405.720 ;
        RECT 1403.990 1404.320 2595.600 1405.680 ;
        RECT 1403.990 1396.880 2596.000 1404.320 ;
        RECT 1404.400 1395.480 2596.000 1396.880 ;
        RECT 1403.990 1394.840 2596.000 1395.480 ;
        RECT 1403.990 1393.440 2595.600 1394.840 ;
        RECT 1403.990 1386.000 2596.000 1393.440 ;
        RECT 1404.400 1384.640 2596.000 1386.000 ;
        RECT 1404.400 1384.600 2595.600 1384.640 ;
        RECT 1403.990 1383.240 2595.600 1384.600 ;
        RECT 1403.990 1375.120 2596.000 1383.240 ;
        RECT 1404.400 1373.760 2596.000 1375.120 ;
        RECT 1404.400 1373.720 2595.600 1373.760 ;
        RECT 1403.990 1372.360 2595.600 1373.720 ;
        RECT 1403.990 1364.920 2596.000 1372.360 ;
        RECT 1404.400 1363.560 2596.000 1364.920 ;
        RECT 1404.400 1363.520 2595.600 1363.560 ;
        RECT 1403.990 1362.160 2595.600 1363.520 ;
        RECT 1403.990 1354.040 2596.000 1362.160 ;
        RECT 1404.400 1352.680 2596.000 1354.040 ;
        RECT 1404.400 1352.640 2595.600 1352.680 ;
        RECT 1403.990 1351.280 2595.600 1352.640 ;
        RECT 1403.990 1343.840 2596.000 1351.280 ;
        RECT 1404.400 1342.480 2596.000 1343.840 ;
        RECT 1404.400 1342.440 2595.600 1342.480 ;
        RECT 1403.990 1341.080 2595.600 1342.440 ;
        RECT 1403.990 1332.960 2596.000 1341.080 ;
        RECT 1404.400 1331.600 2596.000 1332.960 ;
        RECT 1404.400 1331.560 2595.600 1331.600 ;
        RECT 1403.990 1330.200 2595.600 1331.560 ;
        RECT 1403.990 1322.080 2596.000 1330.200 ;
        RECT 1404.400 1321.400 2596.000 1322.080 ;
        RECT 1404.400 1320.680 2595.600 1321.400 ;
        RECT 1403.990 1320.000 2595.600 1320.680 ;
        RECT 1403.990 1311.880 2596.000 1320.000 ;
        RECT 1404.400 1310.520 2596.000 1311.880 ;
        RECT 1404.400 1310.480 2595.600 1310.520 ;
        RECT 1403.990 1309.120 2595.600 1310.480 ;
        RECT 1403.990 1301.000 2596.000 1309.120 ;
        RECT 1404.400 1300.320 2596.000 1301.000 ;
        RECT 1404.400 1299.600 2595.600 1300.320 ;
        RECT 1403.990 1298.920 2595.600 1299.600 ;
        RECT 1403.990 1290.120 2596.000 1298.920 ;
        RECT 1404.400 1289.440 2596.000 1290.120 ;
        RECT 1404.400 1288.720 2595.600 1289.440 ;
        RECT 1403.990 1288.040 2595.600 1288.720 ;
        RECT 1403.990 1279.920 2596.000 1288.040 ;
        RECT 1404.400 1279.240 2596.000 1279.920 ;
        RECT 1404.400 1278.520 2595.600 1279.240 ;
        RECT 1403.990 1277.840 2595.600 1278.520 ;
        RECT 1403.990 1269.040 2596.000 1277.840 ;
        RECT 1404.400 1268.360 2596.000 1269.040 ;
        RECT 1404.400 1267.640 2595.600 1268.360 ;
        RECT 1403.990 1266.960 2595.600 1267.640 ;
        RECT 1403.990 1258.840 2596.000 1266.960 ;
        RECT 1404.400 1258.160 2596.000 1258.840 ;
        RECT 1404.400 1257.440 2595.600 1258.160 ;
        RECT 1403.990 1256.760 2595.600 1257.440 ;
        RECT 1403.990 1247.960 2596.000 1256.760 ;
        RECT 1404.400 1247.280 2596.000 1247.960 ;
        RECT 1404.400 1246.560 2595.600 1247.280 ;
        RECT 1403.990 1245.880 2595.600 1246.560 ;
        RECT 1403.990 1237.080 2596.000 1245.880 ;
        RECT 1404.400 1235.680 2595.600 1237.080 ;
        RECT 1403.990 1226.880 2596.000 1235.680 ;
        RECT 1404.400 1226.200 2596.000 1226.880 ;
        RECT 1404.400 1225.480 2595.600 1226.200 ;
        RECT 1403.990 1224.800 2595.600 1225.480 ;
        RECT 1403.990 1216.000 2596.000 1224.800 ;
        RECT 1404.400 1214.600 2595.600 1216.000 ;
        RECT 1403.990 1205.800 2596.000 1214.600 ;
        RECT 1404.400 1204.935 2595.600 1205.800 ;
      LAYER met3 ;
        RECT 1646.865 1062.660 1647.195 1062.665 ;
        RECT 1646.865 1062.650 1647.450 1062.660 ;
        RECT 1646.640 1062.350 1647.450 1062.650 ;
        RECT 1646.865 1062.340 1647.450 1062.350 ;
        RECT 1646.865 1062.335 1647.195 1062.340 ;
        RECT 1682.030 1038.850 1682.410 1038.860 ;
        RECT 1683.205 1038.850 1683.535 1038.865 ;
        RECT 1682.030 1038.550 1683.535 1038.850 ;
        RECT 1682.030 1038.540 1682.410 1038.550 ;
        RECT 1683.205 1038.535 1683.535 1038.550 ;
        RECT 1704.365 1021.180 1704.695 1021.185 ;
        RECT 1704.110 1021.170 1704.695 1021.180 ;
        RECT 1752.205 1021.170 1752.535 1021.185 ;
        RECT 1704.110 1020.870 1704.920 1021.170 ;
        RECT 1738.880 1020.870 1752.535 1021.170 ;
        RECT 1704.110 1020.860 1704.695 1020.870 ;
        RECT 1704.365 1020.855 1704.695 1020.860 ;
        RECT 1496.905 1020.490 1497.235 1020.505 ;
        RECT 1738.880 1020.490 1739.180 1020.870 ;
        RECT 1752.205 1020.855 1752.535 1020.870 ;
        RECT 1786.705 1021.170 1787.035 1021.185 ;
        RECT 1834.085 1021.170 1834.415 1021.185 ;
        RECT 1834.750 1021.170 1835.130 1021.180 ;
        RECT 1786.705 1020.870 1789.090 1021.170 ;
        RECT 1786.705 1020.855 1787.035 1020.870 ;
        RECT 1496.905 1020.190 1739.180 1020.490 ;
        RECT 1496.905 1020.175 1497.235 1020.190 ;
        RECT 1441.705 1019.810 1442.035 1019.825 ;
        RECT 1776.585 1019.810 1776.915 1019.825 ;
        RECT 1787.165 1019.820 1787.495 1019.825 ;
        RECT 1441.705 1019.510 1776.915 1019.810 ;
        RECT 1441.705 1019.495 1442.035 1019.510 ;
        RECT 1776.585 1019.495 1776.915 1019.510 ;
        RECT 1786.910 1019.810 1787.495 1019.820 ;
        RECT 1788.790 1019.810 1789.090 1020.870 ;
        RECT 1834.085 1020.870 1835.130 1021.170 ;
        RECT 1834.085 1020.855 1834.415 1020.870 ;
        RECT 1834.750 1020.860 1835.130 1020.870 ;
        RECT 1842.365 1021.170 1842.695 1021.185 ;
        RECT 1843.950 1021.170 1844.330 1021.180 ;
        RECT 1842.365 1020.870 1844.330 1021.170 ;
        RECT 1842.365 1020.855 1842.695 1020.870 ;
        RECT 1843.950 1020.860 1844.330 1020.870 ;
        RECT 1854.990 1021.170 1855.370 1021.180 ;
        RECT 1855.705 1021.170 1856.035 1021.185 ;
        RECT 1854.990 1020.870 1856.035 1021.170 ;
        RECT 1854.990 1020.860 1855.370 1020.870 ;
        RECT 1855.705 1020.855 1856.035 1020.870 ;
        RECT 2241.390 1021.170 2241.770 1021.180 ;
        RECT 2242.105 1021.170 2242.435 1021.185 ;
        RECT 2241.390 1020.870 2242.435 1021.170 ;
        RECT 2241.390 1020.860 2241.770 1020.870 ;
        RECT 2242.105 1020.855 2242.435 1020.870 ;
        RECT 2259.585 1021.170 2259.915 1021.185 ;
        RECT 2266.485 1021.180 2266.815 1021.185 ;
        RECT 2260.710 1021.170 2261.090 1021.180 ;
        RECT 2259.585 1020.870 2261.090 1021.170 ;
        RECT 2259.585 1020.855 2259.915 1020.870 ;
        RECT 2260.710 1020.860 2261.090 1020.870 ;
        RECT 2266.230 1021.170 2266.815 1021.180 ;
        RECT 2270.830 1021.170 2271.210 1021.180 ;
        RECT 2276.605 1021.170 2276.935 1021.185 ;
        RECT 2266.230 1020.870 2267.040 1021.170 ;
        RECT 2270.830 1020.870 2276.935 1021.170 ;
        RECT 2266.230 1020.860 2266.815 1020.870 ;
        RECT 2270.830 1020.860 2271.210 1020.870 ;
        RECT 2266.485 1020.855 2266.815 1020.860 ;
        RECT 2276.605 1020.855 2276.935 1020.870 ;
        RECT 2281.870 1021.170 2282.250 1021.180 ;
        RECT 2283.505 1021.170 2283.835 1021.185 ;
        RECT 2281.870 1020.870 2283.835 1021.170 ;
        RECT 2281.870 1020.860 2282.250 1020.870 ;
        RECT 2283.505 1020.855 2283.835 1020.870 ;
        RECT 2328.790 1021.170 2329.170 1021.180 ;
        RECT 2330.885 1021.170 2331.215 1021.185 ;
        RECT 2328.790 1020.870 2331.215 1021.170 ;
        RECT 2328.790 1020.860 2329.170 1020.870 ;
        RECT 2330.885 1020.855 2331.215 1020.870 ;
        RECT 2333.390 1021.170 2333.770 1021.180 ;
        RECT 2338.705 1021.170 2339.035 1021.185 ;
        RECT 2333.390 1020.870 2339.035 1021.170 ;
        RECT 2333.390 1020.860 2333.770 1020.870 ;
        RECT 2338.705 1020.855 2339.035 1020.870 ;
        RECT 2340.750 1021.170 2341.130 1021.180 ;
        RECT 2345.145 1021.170 2345.475 1021.185 ;
        RECT 2340.750 1020.870 2345.475 1021.170 ;
        RECT 2340.750 1020.860 2341.130 1020.870 ;
        RECT 2345.145 1020.855 2345.475 1020.870 ;
        RECT 2351.790 1021.170 2352.170 1021.180 ;
        RECT 2352.505 1021.170 2352.835 1021.185 ;
        RECT 2351.790 1020.870 2352.835 1021.170 ;
        RECT 2351.790 1020.860 2352.170 1020.870 ;
        RECT 2352.505 1020.855 2352.835 1020.870 ;
        RECT 2358.230 1021.170 2358.610 1021.180 ;
        RECT 2359.405 1021.170 2359.735 1021.185 ;
        RECT 2373.665 1021.180 2373.995 1021.185 ;
        RECT 2403.105 1021.180 2403.435 1021.185 ;
        RECT 2421.965 1021.180 2422.295 1021.185 ;
        RECT 2373.665 1021.170 2374.250 1021.180 ;
        RECT 2403.105 1021.170 2403.690 1021.180 ;
        RECT 2358.230 1020.870 2359.735 1021.170 ;
        RECT 2373.440 1020.870 2374.250 1021.170 ;
        RECT 2402.880 1020.870 2403.690 1021.170 ;
        RECT 2358.230 1020.860 2358.610 1020.870 ;
        RECT 2359.405 1020.855 2359.735 1020.870 ;
        RECT 2373.665 1020.860 2374.250 1020.870 ;
        RECT 2403.105 1020.860 2403.690 1020.870 ;
        RECT 2421.710 1021.170 2422.295 1021.180 ;
        RECT 2421.710 1020.870 2422.520 1021.170 ;
        RECT 2421.710 1020.860 2422.295 1020.870 ;
        RECT 2373.665 1020.855 2373.995 1020.860 ;
        RECT 2403.105 1020.855 2403.435 1020.860 ;
        RECT 2421.965 1020.855 2422.295 1020.860 ;
        RECT 1834.545 1020.490 1834.875 1020.505 ;
        RECT 1837.510 1020.490 1837.890 1020.500 ;
        RECT 1834.545 1020.190 1837.890 1020.490 ;
        RECT 1834.545 1020.175 1834.875 1020.190 ;
        RECT 1837.510 1020.180 1837.890 1020.190 ;
        RECT 2245.785 1020.490 2246.115 1020.505 ;
        RECT 2254.525 1020.500 2254.855 1020.505 ;
        RECT 2247.830 1020.490 2248.210 1020.500 ;
        RECT 2245.785 1020.190 2248.210 1020.490 ;
        RECT 2245.785 1020.175 2246.115 1020.190 ;
        RECT 2247.830 1020.180 2248.210 1020.190 ;
        RECT 2254.270 1020.490 2254.855 1020.500 ;
        RECT 2281.205 1020.490 2281.535 1020.505 ;
        RECT 2282.790 1020.490 2283.170 1020.500 ;
        RECT 2254.270 1020.190 2255.080 1020.490 ;
        RECT 2281.205 1020.190 2283.170 1020.490 ;
        RECT 2254.270 1020.180 2254.855 1020.190 ;
        RECT 2254.525 1020.175 2254.855 1020.180 ;
        RECT 2281.205 1020.175 2281.535 1020.190 ;
        RECT 2282.790 1020.180 2283.170 1020.190 ;
        RECT 2346.270 1020.490 2346.650 1020.500 ;
        RECT 2351.585 1020.490 2351.915 1020.505 ;
        RECT 2346.270 1020.190 2351.915 1020.490 ;
        RECT 2346.270 1020.180 2346.650 1020.190 ;
        RECT 2351.585 1020.175 2351.915 1020.190 ;
        RECT 2359.865 1020.490 2360.195 1020.505 ;
        RECT 2360.990 1020.490 2361.370 1020.500 ;
        RECT 2359.865 1020.190 2361.370 1020.490 ;
        RECT 2359.865 1020.175 2360.195 1020.190 ;
        RECT 2360.990 1020.180 2361.370 1020.190 ;
        RECT 2380.565 1020.490 2380.895 1020.505 ;
        RECT 2387.465 1020.500 2387.795 1020.505 ;
        RECT 2450.945 1020.500 2451.275 1020.505 ;
        RECT 2381.230 1020.490 2381.610 1020.500 ;
        RECT 2387.465 1020.490 2388.050 1020.500 ;
        RECT 2450.945 1020.490 2451.530 1020.500 ;
        RECT 2380.565 1020.190 2381.610 1020.490 ;
        RECT 2387.240 1020.190 2388.050 1020.490 ;
        RECT 2450.720 1020.190 2451.530 1020.490 ;
        RECT 2380.565 1020.175 2380.895 1020.190 ;
        RECT 2381.230 1020.180 2381.610 1020.190 ;
        RECT 2387.465 1020.180 2388.050 1020.190 ;
        RECT 2450.945 1020.180 2451.530 1020.190 ;
        RECT 2387.465 1020.175 2387.795 1020.180 ;
        RECT 2450.945 1020.175 2451.275 1020.180 ;
        RECT 1801.630 1019.810 1802.010 1019.820 ;
        RECT 1786.910 1019.510 1787.720 1019.810 ;
        RECT 1788.790 1019.510 1802.010 1019.810 ;
        RECT 1786.910 1019.500 1787.495 1019.510 ;
        RECT 1801.630 1019.500 1802.010 1019.510 ;
        RECT 1831.990 1019.810 1832.370 1019.820 ;
        RECT 1835.005 1019.810 1835.335 1019.825 ;
        RECT 1831.990 1019.510 1835.335 1019.810 ;
        RECT 1831.990 1019.500 1832.370 1019.510 ;
        RECT 1787.165 1019.495 1787.495 1019.500 ;
        RECT 1835.005 1019.495 1835.335 1019.510 ;
        RECT 2272.670 1019.810 2273.050 1019.820 ;
        RECT 2273.385 1019.810 2273.715 1019.825 ;
        RECT 2276.605 1019.820 2276.935 1019.825 ;
        RECT 2272.670 1019.510 2273.715 1019.810 ;
        RECT 2272.670 1019.500 2273.050 1019.510 ;
        RECT 2273.385 1019.495 2273.715 1019.510 ;
        RECT 2276.350 1019.810 2276.935 1019.820 ;
        RECT 2276.350 1019.510 2277.160 1019.810 ;
        RECT 2276.350 1019.500 2276.935 1019.510 ;
        RECT 2276.605 1019.495 2276.935 1019.500 ;
        RECT 1448.605 1019.130 1448.935 1019.145 ;
        RECT 1808.070 1019.130 1808.450 1019.140 ;
        RECT 1448.605 1018.830 1808.450 1019.130 ;
        RECT 1448.605 1018.815 1448.935 1018.830 ;
        RECT 1808.070 1018.820 1808.450 1018.830 ;
        RECT 1814.305 1019.130 1814.635 1019.145 ;
        RECT 2429.070 1019.130 2429.450 1019.140 ;
        RECT 1814.305 1018.830 2429.450 1019.130 ;
        RECT 1814.305 1018.815 1814.635 1018.830 ;
        RECT 2429.070 1018.820 2429.450 1018.830 ;
        RECT 1711.265 1018.460 1711.595 1018.465 ;
        RECT 1711.265 1018.450 1711.850 1018.460 ;
        RECT 1711.040 1018.150 1711.850 1018.450 ;
        RECT 1711.265 1018.140 1711.850 1018.150 ;
        RECT 1718.165 1018.450 1718.495 1018.465 ;
        RECT 1745.765 1018.460 1746.095 1018.465 ;
        RECT 1719.750 1018.450 1720.130 1018.460 ;
        RECT 1718.165 1018.150 1720.130 1018.450 ;
        RECT 1711.265 1018.135 1711.595 1018.140 ;
        RECT 1718.165 1018.135 1718.495 1018.150 ;
        RECT 1719.750 1018.140 1720.130 1018.150 ;
        RECT 1745.510 1018.450 1746.095 1018.460 ;
        RECT 1759.565 1018.450 1759.895 1018.465 ;
        RECT 1763.910 1018.450 1764.290 1018.460 ;
        RECT 1745.510 1018.150 1746.320 1018.450 ;
        RECT 1759.565 1018.150 1764.290 1018.450 ;
        RECT 1745.510 1018.140 1746.095 1018.150 ;
        RECT 1745.765 1018.135 1746.095 1018.140 ;
        RECT 1759.565 1018.135 1759.895 1018.150 ;
        RECT 1763.910 1018.140 1764.290 1018.150 ;
        RECT 1773.365 1018.450 1773.695 1018.465 ;
        RECT 1774.030 1018.450 1774.410 1018.460 ;
        RECT 1773.365 1018.150 1774.410 1018.450 ;
        RECT 1773.365 1018.135 1773.695 1018.150 ;
        RECT 1774.030 1018.140 1774.410 1018.150 ;
        RECT 1793.605 1018.450 1793.935 1018.465 ;
        RECT 2408.165 1018.450 2408.495 1018.465 ;
        RECT 2408.830 1018.450 2409.210 1018.460 ;
        RECT 1793.605 1018.150 2407.330 1018.450 ;
        RECT 1793.605 1018.135 1793.935 1018.150 ;
        RECT 1711.265 1017.770 1711.595 1017.785 ;
        RECT 1714.230 1017.770 1714.610 1017.780 ;
        RECT 1711.265 1017.470 1714.610 1017.770 ;
        RECT 1711.265 1017.455 1711.595 1017.470 ;
        RECT 1714.230 1017.460 1714.610 1017.470 ;
        RECT 1779.805 1017.770 1780.135 1017.785 ;
        RECT 1779.805 1017.470 2406.410 1017.770 ;
        RECT 1779.805 1017.455 1780.135 1017.470 ;
        RECT 1641.805 1017.100 1642.135 1017.105 ;
        RECT 1654.685 1017.100 1655.015 1017.105 ;
        RECT 1641.550 1017.090 1642.135 1017.100 ;
        RECT 1654.430 1017.090 1655.015 1017.100 ;
        RECT 1670.990 1017.090 1671.370 1017.100 ;
        RECT 1675.845 1017.090 1676.175 1017.105 ;
        RECT 1641.550 1016.790 1642.360 1017.090 ;
        RECT 1654.430 1016.790 1655.240 1017.090 ;
        RECT 1670.990 1016.790 1676.175 1017.090 ;
        RECT 1641.550 1016.780 1642.135 1016.790 ;
        RECT 1654.430 1016.780 1655.015 1016.790 ;
        RECT 1670.990 1016.780 1671.370 1016.790 ;
        RECT 1641.805 1016.775 1642.135 1016.780 ;
        RECT 1654.685 1016.775 1655.015 1016.780 ;
        RECT 1675.845 1016.775 1676.175 1016.790 ;
        RECT 1683.665 1017.090 1683.995 1017.105 ;
        RECT 1684.790 1017.090 1685.170 1017.100 ;
        RECT 1683.665 1016.790 1685.170 1017.090 ;
        RECT 1683.665 1016.775 1683.995 1016.790 ;
        RECT 1684.790 1016.780 1685.170 1016.790 ;
        RECT 1776.585 1017.090 1776.915 1017.105 ;
        RECT 1821.665 1017.100 1821.995 1017.105 ;
        RECT 1814.510 1017.090 1814.890 1017.100 ;
        RECT 1776.585 1016.790 1814.890 1017.090 ;
        RECT 1776.585 1016.775 1776.915 1016.790 ;
        RECT 1814.510 1016.780 1814.890 1016.790 ;
        RECT 1821.665 1017.090 1822.250 1017.100 ;
        RECT 2264.390 1017.090 2264.770 1017.100 ;
        RECT 2269.705 1017.090 2270.035 1017.105 ;
        RECT 2280.285 1017.100 2280.615 1017.105 ;
        RECT 2280.030 1017.090 2280.615 1017.100 ;
        RECT 2283.505 1017.090 2283.835 1017.105 ;
        RECT 1821.665 1016.790 1822.450 1017.090 ;
        RECT 2264.390 1016.790 2270.035 1017.090 ;
        RECT 2279.650 1016.790 2283.835 1017.090 ;
        RECT 1821.665 1016.780 1822.250 1016.790 ;
        RECT 2264.390 1016.780 2264.770 1016.790 ;
        RECT 1821.665 1016.775 1821.995 1016.780 ;
        RECT 2269.705 1016.775 2270.035 1016.790 ;
        RECT 2280.030 1016.780 2280.615 1016.790 ;
        RECT 2280.285 1016.775 2280.615 1016.780 ;
        RECT 2283.505 1016.775 2283.835 1016.790 ;
        RECT 2300.270 1017.090 2300.650 1017.100 ;
        RECT 2304.205 1017.090 2304.535 1017.105 ;
        RECT 2300.270 1016.790 2304.535 1017.090 ;
        RECT 2300.270 1016.780 2300.650 1016.790 ;
        RECT 2304.205 1016.775 2304.535 1016.790 ;
        RECT 2311.310 1017.090 2311.690 1017.100 ;
        RECT 2317.545 1017.090 2317.875 1017.105 ;
        RECT 2311.310 1016.790 2317.875 1017.090 ;
        RECT 2311.310 1016.780 2311.690 1016.790 ;
        RECT 2317.545 1016.775 2317.875 1016.790 ;
        RECT 2387.925 1017.090 2388.255 1017.105 ;
        RECT 2393.190 1017.090 2393.570 1017.100 ;
        RECT 2387.925 1016.790 2393.570 1017.090 ;
        RECT 2387.925 1016.775 2388.255 1016.790 ;
        RECT 2393.190 1016.780 2393.570 1016.790 ;
        RECT 2394.365 1017.090 2394.695 1017.105 ;
        RECT 2395.950 1017.090 2396.330 1017.100 ;
        RECT 2394.365 1016.790 2396.330 1017.090 ;
        RECT 2394.365 1016.775 2394.695 1016.790 ;
        RECT 2395.950 1016.780 2396.330 1016.790 ;
        RECT 1640.630 1016.410 1641.010 1016.420 ;
        RECT 1641.345 1016.410 1641.675 1016.425 ;
        RECT 1640.630 1016.110 1641.675 1016.410 ;
        RECT 1640.630 1016.100 1641.010 1016.110 ;
        RECT 1641.345 1016.095 1641.675 1016.110 ;
        RECT 1653.510 1016.410 1653.890 1016.420 ;
        RECT 1655.605 1016.410 1655.935 1016.425 ;
        RECT 1653.510 1016.110 1655.935 1016.410 ;
        RECT 1653.510 1016.100 1653.890 1016.110 ;
        RECT 1655.605 1016.095 1655.935 1016.110 ;
        RECT 1658.110 1016.410 1658.490 1016.420 ;
        RECT 1662.505 1016.410 1662.835 1016.425 ;
        RECT 1658.110 1016.110 1662.835 1016.410 ;
        RECT 1658.110 1016.100 1658.490 1016.110 ;
        RECT 1662.505 1016.095 1662.835 1016.110 ;
        RECT 1664.550 1016.410 1664.930 1016.420 ;
        RECT 1669.405 1016.410 1669.735 1016.425 ;
        RECT 1664.550 1016.110 1669.735 1016.410 ;
        RECT 1664.550 1016.100 1664.930 1016.110 ;
        RECT 1669.405 1016.095 1669.735 1016.110 ;
        RECT 1675.590 1016.410 1675.970 1016.420 ;
        RECT 1676.305 1016.410 1676.635 1016.425 ;
        RECT 1675.590 1016.110 1676.635 1016.410 ;
        RECT 1675.590 1016.100 1675.970 1016.110 ;
        RECT 1676.305 1016.095 1676.635 1016.110 ;
        RECT 1691.025 1016.410 1691.355 1016.425 ;
        RECT 1692.150 1016.410 1692.530 1016.420 ;
        RECT 1691.025 1016.110 1692.530 1016.410 ;
        RECT 1691.025 1016.095 1691.355 1016.110 ;
        RECT 1692.150 1016.100 1692.530 1016.110 ;
        RECT 1697.925 1016.410 1698.255 1016.425 ;
        RECT 1698.590 1016.410 1698.970 1016.420 ;
        RECT 1697.925 1016.110 1698.970 1016.410 ;
        RECT 1697.925 1016.095 1698.255 1016.110 ;
        RECT 1698.590 1016.100 1698.970 1016.110 ;
        RECT 1725.065 1016.410 1725.395 1016.425 ;
        RECT 1726.190 1016.410 1726.570 1016.420 ;
        RECT 1725.065 1016.110 1726.570 1016.410 ;
        RECT 1725.065 1016.095 1725.395 1016.110 ;
        RECT 1726.190 1016.100 1726.570 1016.110 ;
        RECT 1731.965 1016.410 1732.295 1016.425 ;
        RECT 1732.630 1016.410 1733.010 1016.420 ;
        RECT 1731.965 1016.110 1733.010 1016.410 ;
        RECT 1731.965 1016.095 1732.295 1016.110 ;
        RECT 1732.630 1016.100 1733.010 1016.110 ;
        RECT 1745.765 1016.410 1746.095 1016.425 ;
        RECT 1780.265 1016.420 1780.595 1016.425 ;
        RECT 1749.190 1016.410 1749.570 1016.420 ;
        RECT 1780.265 1016.410 1780.850 1016.420 ;
        RECT 1745.765 1016.110 1749.570 1016.410 ;
        RECT 1780.040 1016.110 1780.850 1016.410 ;
        RECT 1745.765 1016.095 1746.095 1016.110 ;
        RECT 1749.190 1016.100 1749.570 1016.110 ;
        RECT 1780.265 1016.100 1780.850 1016.110 ;
        RECT 2287.185 1016.410 2287.515 1016.425 ;
        RECT 2289.230 1016.410 2289.610 1016.420 ;
        RECT 2287.185 1016.110 2289.610 1016.410 ;
        RECT 1780.265 1016.095 1780.595 1016.100 ;
        RECT 2287.185 1016.095 2287.515 1016.110 ;
        RECT 2289.230 1016.100 2289.610 1016.110 ;
        RECT 2293.830 1016.410 2294.210 1016.420 ;
        RECT 2296.845 1016.410 2297.175 1016.425 ;
        RECT 2293.830 1016.110 2297.175 1016.410 ;
        RECT 2293.830 1016.100 2294.210 1016.110 ;
        RECT 2296.845 1016.095 2297.175 1016.110 ;
        RECT 2304.870 1016.410 2305.250 1016.420 ;
        RECT 2311.105 1016.410 2311.435 1016.425 ;
        RECT 2304.870 1016.110 2311.435 1016.410 ;
        RECT 2304.870 1016.100 2305.250 1016.110 ;
        RECT 2311.105 1016.095 2311.435 1016.110 ;
        RECT 2315.910 1016.410 2316.290 1016.420 ;
        RECT 2318.005 1016.410 2318.335 1016.425 ;
        RECT 2315.910 1016.110 2318.335 1016.410 ;
        RECT 2315.910 1016.100 2316.290 1016.110 ;
        RECT 2318.005 1016.095 2318.335 1016.110 ;
        RECT 2322.350 1016.410 2322.730 1016.420 ;
        RECT 2324.445 1016.410 2324.775 1016.425 ;
        RECT 2322.350 1016.110 2324.775 1016.410 ;
        RECT 2322.350 1016.100 2322.730 1016.110 ;
        RECT 2324.445 1016.095 2324.775 1016.110 ;
        RECT 2355.265 1016.410 2355.595 1016.425 ;
        RECT 2359.150 1016.410 2359.530 1016.420 ;
        RECT 2381.025 1016.410 2381.355 1016.425 ;
        RECT 2355.265 1016.110 2381.355 1016.410 ;
        RECT 2355.265 1016.095 2355.595 1016.110 ;
        RECT 2359.150 1016.100 2359.530 1016.110 ;
        RECT 2381.025 1016.095 2381.355 1016.110 ;
        RECT 2388.385 1016.410 2388.715 1016.425 ;
        RECT 2390.430 1016.410 2390.810 1016.420 ;
        RECT 2388.385 1016.110 2390.810 1016.410 ;
        RECT 2406.110 1016.410 2406.410 1017.470 ;
        RECT 2407.030 1017.090 2407.330 1018.150 ;
        RECT 2408.165 1018.150 2409.210 1018.450 ;
        RECT 2408.165 1018.135 2408.495 1018.150 ;
        RECT 2408.830 1018.140 2409.210 1018.150 ;
        RECT 2428.865 1018.450 2429.195 1018.465 ;
        RECT 2431.830 1018.450 2432.210 1018.460 ;
        RECT 2428.865 1018.150 2432.210 1018.450 ;
        RECT 2428.865 1018.135 2429.195 1018.150 ;
        RECT 2431.830 1018.140 2432.210 1018.150 ;
        RECT 2408.165 1017.770 2408.495 1017.785 ;
        RECT 2410.670 1017.770 2411.050 1017.780 ;
        RECT 2437.350 1017.770 2437.730 1017.780 ;
        RECT 2408.165 1017.470 2411.050 1017.770 ;
        RECT 2408.165 1017.455 2408.495 1017.470 ;
        RECT 2410.670 1017.460 2411.050 1017.470 ;
        RECT 2412.550 1017.470 2437.730 1017.770 ;
        RECT 2412.550 1017.090 2412.850 1017.470 ;
        RECT 2437.350 1017.460 2437.730 1017.470 ;
        RECT 2415.065 1017.100 2415.395 1017.105 ;
        RECT 2415.065 1017.090 2415.650 1017.100 ;
        RECT 2407.030 1016.790 2412.850 1017.090 ;
        RECT 2414.840 1016.790 2415.650 1017.090 ;
        RECT 2415.065 1016.780 2415.650 1016.790 ;
        RECT 2421.965 1017.090 2422.295 1017.105 ;
        RECT 2423.550 1017.090 2423.930 1017.100 ;
        RECT 2421.965 1016.790 2423.930 1017.090 ;
        RECT 2415.065 1016.775 2415.395 1016.780 ;
        RECT 2421.965 1016.775 2422.295 1016.790 ;
        RECT 2423.550 1016.780 2423.930 1016.790 ;
        RECT 2442.870 1016.410 2443.250 1016.420 ;
        RECT 2406.110 1016.110 2443.250 1016.410 ;
        RECT 2388.385 1016.095 2388.715 1016.110 ;
        RECT 2390.430 1016.100 2390.810 1016.110 ;
        RECT 2442.870 1016.100 2443.250 1016.110 ;
        RECT 1662.045 1015.740 1662.375 1015.745 ;
        RECT 1661.790 1015.730 1662.375 1015.740 ;
        RECT 1668.230 1015.730 1668.610 1015.740 ;
        RECT 1668.945 1015.730 1669.275 1015.745 ;
        RECT 1661.790 1015.430 1662.600 1015.730 ;
        RECT 1668.230 1015.430 1669.275 1015.730 ;
        RECT 1661.790 1015.420 1662.375 1015.430 ;
        RECT 1668.230 1015.420 1668.610 1015.430 ;
        RECT 1662.045 1015.415 1662.375 1015.420 ;
        RECT 1668.945 1015.415 1669.275 1015.430 ;
        RECT 1673.750 1015.730 1674.130 1015.740 ;
        RECT 1675.385 1015.730 1675.715 1015.745 ;
        RECT 1683.205 1015.740 1683.535 1015.745 ;
        RECT 1673.750 1015.430 1675.715 1015.730 ;
        RECT 1673.750 1015.420 1674.130 1015.430 ;
        RECT 1675.385 1015.415 1675.715 1015.430 ;
        RECT 1682.950 1015.730 1683.535 1015.740 ;
        RECT 1738.865 1015.740 1739.195 1015.745 ;
        RECT 1755.425 1015.740 1755.755 1015.745 ;
        RECT 1766.465 1015.740 1766.795 1015.745 ;
        RECT 1738.865 1015.730 1739.450 1015.740 ;
        RECT 1755.425 1015.730 1756.010 1015.740 ;
        RECT 1766.465 1015.730 1767.050 1015.740 ;
        RECT 1682.950 1015.430 1683.760 1015.730 ;
        RECT 1738.640 1015.430 1739.450 1015.730 ;
        RECT 1755.200 1015.430 1756.010 1015.730 ;
        RECT 1766.240 1015.430 1767.050 1015.730 ;
        RECT 1682.950 1015.420 1683.535 1015.430 ;
        RECT 1683.205 1015.415 1683.535 1015.420 ;
        RECT 1738.865 1015.420 1739.450 1015.430 ;
        RECT 1755.425 1015.420 1756.010 1015.430 ;
        RECT 1766.465 1015.420 1767.050 1015.430 ;
        RECT 1787.625 1015.730 1787.955 1015.745 ;
        RECT 1788.750 1015.730 1789.130 1015.740 ;
        RECT 1787.625 1015.430 1789.130 1015.730 ;
        RECT 1738.865 1015.415 1739.195 1015.420 ;
        RECT 1755.425 1015.415 1755.755 1015.420 ;
        RECT 1766.465 1015.415 1766.795 1015.420 ;
        RECT 1787.625 1015.415 1787.955 1015.430 ;
        RECT 1788.750 1015.420 1789.130 1015.430 ;
        RECT 1647.990 1015.050 1648.370 1015.060 ;
        RECT 1648.705 1015.050 1649.035 1015.065 ;
        RECT 1647.990 1014.750 1649.035 1015.050 ;
        RECT 1647.990 1014.740 1648.370 1014.750 ;
        RECT 1648.705 1014.735 1649.035 1014.750 ;
        RECT 1680.190 1015.050 1680.570 1015.060 ;
        RECT 1683.205 1015.050 1683.535 1015.065 ;
        RECT 1689.645 1015.060 1689.975 1015.065 ;
        RECT 1696.085 1015.060 1696.415 1015.065 ;
        RECT 1700.685 1015.060 1701.015 1015.065 ;
        RECT 1707.125 1015.060 1707.455 1015.065 ;
        RECT 1713.565 1015.060 1713.895 1015.065 ;
        RECT 1718.165 1015.060 1718.495 1015.065 ;
        RECT 1724.605 1015.060 1724.935 1015.065 ;
        RECT 1689.390 1015.050 1689.975 1015.060 ;
        RECT 1695.830 1015.050 1696.415 1015.060 ;
        RECT 1700.430 1015.050 1701.015 1015.060 ;
        RECT 1706.870 1015.050 1707.455 1015.060 ;
        RECT 1713.310 1015.050 1713.895 1015.060 ;
        RECT 1717.910 1015.050 1718.495 1015.060 ;
        RECT 1724.350 1015.050 1724.935 1015.060 ;
        RECT 1680.190 1014.750 1683.535 1015.050 ;
        RECT 1689.190 1014.750 1689.975 1015.050 ;
        RECT 1695.630 1014.750 1696.415 1015.050 ;
        RECT 1700.230 1014.750 1701.015 1015.050 ;
        RECT 1706.670 1014.750 1707.455 1015.050 ;
        RECT 1713.110 1014.750 1713.895 1015.050 ;
        RECT 1717.710 1014.750 1718.495 1015.050 ;
        RECT 1724.150 1014.750 1724.935 1015.050 ;
        RECT 1680.190 1014.740 1680.570 1014.750 ;
        RECT 1683.205 1014.735 1683.535 1014.750 ;
        RECT 1689.390 1014.740 1689.975 1014.750 ;
        RECT 1695.830 1014.740 1696.415 1014.750 ;
        RECT 1700.430 1014.740 1701.015 1014.750 ;
        RECT 1706.870 1014.740 1707.455 1014.750 ;
        RECT 1713.310 1014.740 1713.895 1014.750 ;
        RECT 1717.910 1014.740 1718.495 1014.750 ;
        RECT 1724.350 1014.740 1724.935 1014.750 ;
        RECT 1689.645 1014.735 1689.975 1014.740 ;
        RECT 1696.085 1014.735 1696.415 1014.740 ;
        RECT 1700.685 1014.735 1701.015 1014.740 ;
        RECT 1707.125 1014.735 1707.455 1014.740 ;
        RECT 1713.565 1014.735 1713.895 1014.740 ;
        RECT 1718.165 1014.735 1718.495 1014.740 ;
        RECT 1724.605 1014.735 1724.935 1014.740 ;
        RECT 1729.665 1015.050 1729.995 1015.065 ;
        RECT 1735.645 1015.060 1735.975 1015.065 ;
        RECT 1730.790 1015.050 1731.170 1015.060 ;
        RECT 1735.390 1015.050 1735.975 1015.060 ;
        RECT 1729.665 1014.750 1731.170 1015.050 ;
        RECT 1735.190 1014.750 1735.975 1015.050 ;
        RECT 1729.665 1014.735 1729.995 1014.750 ;
        RECT 1730.790 1014.740 1731.170 1014.750 ;
        RECT 1735.390 1014.740 1735.975 1014.750 ;
        RECT 1735.645 1014.735 1735.975 1014.740 ;
        RECT 1741.625 1015.060 1741.955 1015.065 ;
        RECT 1748.065 1015.060 1748.395 1015.065 ;
        RECT 1741.625 1015.050 1742.210 1015.060 ;
        RECT 1748.065 1015.050 1748.650 1015.060 ;
        RECT 1754.710 1015.050 1755.090 1015.060 ;
        RECT 1755.885 1015.050 1756.215 1015.065 ;
        RECT 1741.625 1014.750 1742.410 1015.050 ;
        RECT 1748.065 1014.750 1748.850 1015.050 ;
        RECT 1754.710 1014.750 1756.215 1015.050 ;
        RECT 1741.625 1014.740 1742.210 1014.750 ;
        RECT 1748.065 1014.740 1748.650 1014.750 ;
        RECT 1754.710 1014.740 1755.090 1014.750 ;
        RECT 1741.625 1014.735 1741.955 1014.740 ;
        RECT 1748.065 1014.735 1748.395 1014.740 ;
        RECT 1755.885 1014.735 1756.215 1014.750 ;
        RECT 1758.390 1015.050 1758.770 1015.060 ;
        RECT 1759.105 1015.050 1759.435 1015.065 ;
        RECT 1766.005 1015.060 1766.335 1015.065 ;
        RECT 1765.750 1015.050 1766.335 1015.060 ;
        RECT 1758.390 1014.750 1759.435 1015.050 ;
        RECT 1765.550 1014.750 1766.335 1015.050 ;
        RECT 1758.390 1014.740 1758.770 1014.750 ;
        RECT 1759.105 1014.735 1759.435 1014.750 ;
        RECT 1765.750 1014.740 1766.335 1014.750 ;
        RECT 1772.190 1015.050 1772.570 1015.060 ;
        RECT 1772.905 1015.050 1773.235 1015.065 ;
        RECT 1777.965 1015.060 1778.295 1015.065 ;
        RECT 1777.710 1015.050 1778.295 1015.060 ;
        RECT 1772.190 1014.750 1773.235 1015.050 ;
        RECT 1777.510 1014.750 1778.295 1015.050 ;
        RECT 1772.190 1014.740 1772.570 1014.750 ;
        RECT 1766.005 1014.735 1766.335 1014.740 ;
        RECT 1772.905 1014.735 1773.235 1014.750 ;
        RECT 1777.710 1014.740 1778.295 1014.750 ;
        RECT 1777.965 1014.735 1778.295 1014.740 ;
        RECT 1782.105 1015.060 1782.435 1015.065 ;
        RECT 1782.105 1015.050 1782.690 1015.060 ;
        RECT 1787.165 1015.050 1787.495 1015.065 ;
        RECT 1789.670 1015.050 1790.050 1015.060 ;
        RECT 1782.105 1014.750 1782.890 1015.050 ;
        RECT 1787.165 1014.750 1790.050 1015.050 ;
        RECT 1782.105 1014.740 1782.690 1014.750 ;
        RECT 1782.105 1014.735 1782.435 1014.740 ;
        RECT 1787.165 1014.735 1787.495 1014.750 ;
        RECT 1789.670 1014.740 1790.050 1014.750 ;
        RECT 1790.385 1015.050 1790.715 1015.065 ;
        RECT 1793.350 1015.050 1793.730 1015.060 ;
        RECT 1790.385 1014.750 1793.730 1015.050 ;
        RECT 1790.385 1014.735 1790.715 1014.750 ;
        RECT 1793.350 1014.740 1793.730 1014.750 ;
        RECT 1794.065 1015.050 1794.395 1015.065 ;
        RECT 1800.045 1015.060 1800.375 1015.065 ;
        RECT 1796.110 1015.050 1796.490 1015.060 ;
        RECT 1799.790 1015.050 1800.375 1015.060 ;
        RECT 1794.065 1014.750 1796.490 1015.050 ;
        RECT 1799.590 1014.750 1800.375 1015.050 ;
        RECT 1794.065 1014.735 1794.395 1014.750 ;
        RECT 1796.110 1014.740 1796.490 1014.750 ;
        RECT 1799.790 1014.740 1800.375 1014.750 ;
        RECT 1800.045 1014.735 1800.375 1014.740 ;
        RECT 1806.025 1015.060 1806.355 1015.065 ;
        RECT 1812.925 1015.060 1813.255 1015.065 ;
        RECT 1817.525 1015.060 1817.855 1015.065 ;
        RECT 1823.965 1015.060 1824.295 1015.065 ;
        RECT 1806.025 1015.050 1806.610 1015.060 ;
        RECT 1812.670 1015.050 1813.255 1015.060 ;
        RECT 1817.270 1015.050 1817.855 1015.060 ;
        RECT 1823.710 1015.050 1824.295 1015.060 ;
        RECT 1806.025 1014.750 1806.810 1015.050 ;
        RECT 1812.470 1014.750 1813.255 1015.050 ;
        RECT 1817.070 1014.750 1817.855 1015.050 ;
        RECT 1823.510 1014.750 1824.295 1015.050 ;
        RECT 1806.025 1014.740 1806.610 1014.750 ;
        RECT 1812.670 1014.740 1813.255 1014.750 ;
        RECT 1817.270 1014.740 1817.855 1014.750 ;
        RECT 1823.710 1014.740 1824.295 1014.750 ;
        RECT 2246.910 1015.050 2247.290 1015.060 ;
        RECT 2249.005 1015.050 2249.335 1015.065 ;
        RECT 2246.910 1014.750 2249.335 1015.050 ;
        RECT 2246.910 1014.740 2247.290 1014.750 ;
        RECT 1806.025 1014.735 1806.355 1014.740 ;
        RECT 1812.925 1014.735 1813.255 1014.740 ;
        RECT 1817.525 1014.735 1817.855 1014.740 ;
        RECT 1823.965 1014.735 1824.295 1014.740 ;
        RECT 2249.005 1014.735 2249.335 1014.750 ;
        RECT 2253.350 1015.050 2253.730 1015.060 ;
        RECT 2254.985 1015.050 2255.315 1015.065 ;
        RECT 2253.350 1014.750 2255.315 1015.050 ;
        RECT 2253.350 1014.740 2253.730 1014.750 ;
        RECT 2254.985 1014.735 2255.315 1014.750 ;
        RECT 2258.870 1015.050 2259.250 1015.060 ;
        RECT 2262.805 1015.050 2263.135 1015.065 ;
        RECT 2258.870 1014.750 2263.135 1015.050 ;
        RECT 2258.870 1014.740 2259.250 1014.750 ;
        RECT 2262.805 1014.735 2263.135 1014.750 ;
        RECT 2287.390 1015.050 2287.770 1015.060 ;
        RECT 2289.945 1015.050 2290.275 1015.065 ;
        RECT 2287.390 1014.750 2290.275 1015.050 ;
        RECT 2287.390 1014.740 2287.770 1014.750 ;
        RECT 2289.945 1014.735 2290.275 1014.750 ;
        RECT 2293.625 1015.050 2293.955 1015.065 ;
        RECT 2303.285 1015.060 2303.615 1015.065 ;
        RECT 2307.885 1015.060 2308.215 1015.065 ;
        RECT 2294.750 1015.050 2295.130 1015.060 ;
        RECT 2303.030 1015.050 2303.615 1015.060 ;
        RECT 2307.630 1015.050 2308.215 1015.060 ;
        RECT 2293.625 1014.750 2295.130 1015.050 ;
        RECT 2302.830 1014.750 2303.615 1015.050 ;
        RECT 2307.430 1014.750 2308.215 1015.050 ;
        RECT 2293.625 1014.735 2293.955 1014.750 ;
        RECT 2294.750 1014.740 2295.130 1014.750 ;
        RECT 2303.030 1014.740 2303.615 1014.750 ;
        RECT 2307.630 1014.740 2308.215 1014.750 ;
        RECT 2303.285 1014.735 2303.615 1014.740 ;
        RECT 2307.885 1014.735 2308.215 1014.740 ;
        RECT 2312.025 1015.060 2312.355 1015.065 ;
        RECT 2312.025 1015.050 2312.610 1015.060 ;
        RECT 2317.085 1015.050 2317.415 1015.065 ;
        RECT 2323.525 1015.060 2323.855 1015.065 ;
        RECT 2317.750 1015.050 2318.130 1015.060 ;
        RECT 2323.270 1015.050 2323.855 1015.060 ;
        RECT 2312.025 1014.750 2312.810 1015.050 ;
        RECT 2317.085 1014.750 2318.130 1015.050 ;
        RECT 2323.070 1014.750 2323.855 1015.050 ;
        RECT 2312.025 1014.740 2312.610 1014.750 ;
        RECT 2312.025 1014.735 2312.355 1014.740 ;
        RECT 2317.085 1014.735 2317.415 1014.750 ;
        RECT 2317.750 1014.740 2318.130 1014.750 ;
        RECT 2323.270 1014.740 2323.855 1014.750 ;
        RECT 2323.525 1014.735 2323.855 1014.740 ;
        RECT 2329.505 1015.060 2329.835 1015.065 ;
        RECT 2335.485 1015.060 2335.815 1015.065 ;
        RECT 2329.505 1015.050 2330.090 1015.060 ;
        RECT 2335.230 1015.050 2335.815 1015.060 ;
        RECT 2329.505 1014.750 2330.290 1015.050 ;
        RECT 2335.030 1014.750 2335.815 1015.050 ;
        RECT 2329.505 1014.740 2330.090 1014.750 ;
        RECT 2335.230 1014.740 2335.815 1014.750 ;
        RECT 2329.505 1014.735 2329.835 1014.740 ;
        RECT 2335.485 1014.735 2335.815 1014.740 ;
        RECT 2342.385 1015.060 2342.715 1015.065 ;
        RECT 2346.985 1015.060 2347.315 1015.065 ;
        RECT 2355.725 1015.060 2356.055 1015.065 ;
        RECT 2342.385 1015.050 2342.970 1015.060 ;
        RECT 2346.985 1015.050 2347.570 1015.060 ;
        RECT 2355.470 1015.050 2356.055 1015.060 ;
        RECT 2342.385 1014.750 2343.170 1015.050 ;
        RECT 2346.985 1014.750 2347.770 1015.050 ;
        RECT 2355.270 1014.750 2356.055 1015.050 ;
        RECT 2342.385 1014.740 2342.970 1014.750 ;
        RECT 2346.985 1014.740 2347.570 1014.750 ;
        RECT 2355.470 1014.740 2356.055 1014.750 ;
        RECT 2342.385 1014.735 2342.715 1014.740 ;
        RECT 2346.985 1014.735 2347.315 1014.740 ;
        RECT 2355.725 1014.735 2356.055 1014.740 ;
        RECT 2363.545 1015.050 2363.875 1015.065 ;
        RECT 2364.670 1015.050 2365.050 1015.060 ;
        RECT 2363.545 1014.750 2365.050 1015.050 ;
        RECT 2363.545 1014.735 2363.875 1014.750 ;
        RECT 2364.670 1014.740 2365.050 1014.750 ;
        RECT 2366.765 1015.050 2367.095 1015.065 ;
        RECT 2373.205 1015.060 2373.535 1015.065 ;
        RECT 2377.805 1015.060 2378.135 1015.065 ;
        RECT 2367.430 1015.050 2367.810 1015.060 ;
        RECT 2372.950 1015.050 2373.535 1015.060 ;
        RECT 2377.550 1015.050 2378.135 1015.060 ;
        RECT 2366.765 1014.750 2367.810 1015.050 ;
        RECT 2372.750 1014.750 2373.535 1015.050 ;
        RECT 2377.350 1014.750 2378.135 1015.050 ;
        RECT 2366.765 1014.735 2367.095 1014.750 ;
        RECT 2367.430 1014.740 2367.810 1014.750 ;
        RECT 2372.950 1014.740 2373.535 1014.750 ;
        RECT 2377.550 1014.740 2378.135 1014.750 ;
        RECT 2373.205 1014.735 2373.535 1014.740 ;
        RECT 2377.805 1014.735 2378.135 1014.740 ;
        RECT 2380.565 1015.050 2380.895 1015.065 ;
        RECT 2382.150 1015.050 2382.530 1015.060 ;
        RECT 2380.565 1014.750 2382.530 1015.050 ;
        RECT 2380.565 1014.735 2380.895 1014.750 ;
        RECT 2382.150 1014.740 2382.530 1014.750 ;
        RECT 2387.465 1015.050 2387.795 1015.065 ;
        RECT 2388.590 1015.050 2388.970 1015.060 ;
        RECT 2387.465 1014.750 2388.970 1015.050 ;
        RECT 2387.465 1014.735 2387.795 1014.750 ;
        RECT 2388.590 1014.740 2388.970 1014.750 ;
        RECT 2394.365 1015.050 2394.695 1015.065 ;
        RECT 2399.630 1015.050 2400.010 1015.060 ;
        RECT 2394.365 1014.750 2400.010 1015.050 ;
        RECT 2394.365 1014.735 2394.695 1014.750 ;
        RECT 2399.630 1014.740 2400.010 1014.750 ;
        RECT 2402.185 1015.050 2402.515 1015.065 ;
        RECT 2406.070 1015.050 2406.450 1015.060 ;
        RECT 2402.185 1014.750 2406.450 1015.050 ;
        RECT 2402.185 1014.735 2402.515 1014.750 ;
        RECT 2406.070 1014.740 2406.450 1014.750 ;
        RECT 2415.065 1015.050 2415.395 1015.065 ;
        RECT 2417.110 1015.050 2417.490 1015.060 ;
        RECT 2415.065 1014.750 2417.490 1015.050 ;
        RECT 2415.065 1014.735 2415.395 1014.750 ;
        RECT 2417.110 1014.740 2417.490 1014.750 ;
        RECT 2242.105 1006.900 2242.435 1006.905 ;
        RECT 2241.890 1006.890 2242.435 1006.900 ;
        RECT 2241.650 1006.590 2242.435 1006.890 ;
        RECT 2241.890 1006.580 2242.435 1006.590 ;
        RECT 2242.105 1006.575 2242.435 1006.580 ;
        RECT 1490.005 558.770 1490.335 558.785 ;
        RECT 1490.005 558.470 1503.890 558.770 ;
        RECT 1490.005 558.455 1490.335 558.470 ;
        RECT 1503.590 557.970 1503.890 558.470 ;
        RECT 1500.000 557.670 1504.600 557.970 ;
        RECT 1503.590 556.745 1503.890 557.670 ;
        RECT 1503.590 556.430 1504.135 556.745 ;
        RECT 1503.805 556.415 1504.135 556.430 ;
      LAYER met3 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
      LAYER met3 ;
        RECT 1898.945 913.730 1899.275 913.745 ;
        RECT 1889.070 913.610 1899.275 913.730 ;
        RECT 1881.880 913.430 1899.275 913.610 ;
        RECT 1881.880 913.310 1889.370 913.430 ;
        RECT 1898.945 913.415 1899.275 913.430 ;
        RECT 1884.225 908.290 1884.555 908.305 ;
        RECT 1884.225 907.975 1884.770 908.290 ;
        RECT 1884.470 905.110 1884.770 907.975 ;
        RECT 1881.880 904.810 1886.480 905.110 ;
        RECT 1899.865 615.890 1900.195 615.905 ;
        RECT 1889.070 615.870 1900.195 615.890 ;
        RECT 1881.880 615.590 1900.195 615.870 ;
        RECT 1881.880 615.570 1889.370 615.590 ;
        RECT 1899.865 615.575 1900.195 615.590 ;
        RECT 1902.165 610.450 1902.495 610.465 ;
        RECT 1885.390 610.150 1902.495 610.450 ;
        RECT 1885.390 607.370 1885.690 610.150 ;
        RECT 1902.165 610.135 1902.495 610.150 ;
        RECT 1881.880 607.070 1886.480 607.370 ;
        RECT 1881.880 601.610 1889.370 601.730 ;
        RECT 1901.705 601.610 1902.035 601.625 ;
        RECT 1881.880 601.430 1902.035 601.610 ;
        RECT 1889.070 601.310 1902.035 601.430 ;
        RECT 1901.705 601.295 1902.035 601.310 ;
        RECT 1901.245 593.450 1901.575 593.465 ;
        RECT 1889.070 593.230 1901.575 593.450 ;
        RECT 1881.880 593.150 1901.575 593.230 ;
        RECT 1881.880 592.930 1889.370 593.150 ;
        RECT 1901.245 593.135 1901.575 593.150 ;
        RECT 1900.325 590.730 1900.655 590.745 ;
        RECT 1885.390 590.430 1900.655 590.730 ;
        RECT 1885.390 587.590 1885.690 590.430 ;
        RECT 1900.325 590.415 1900.655 590.430 ;
        RECT 1881.880 587.290 1886.480 587.590 ;
        RECT 1900.325 579.170 1900.655 579.185 ;
        RECT 1889.070 579.090 1900.655 579.170 ;
        RECT 1881.880 578.870 1900.655 579.090 ;
        RECT 1881.880 578.790 1889.370 578.870 ;
        RECT 1900.325 578.855 1900.655 578.870 ;
        RECT 1900.785 573.730 1901.115 573.745 ;
        RECT 1889.070 573.450 1901.115 573.730 ;
        RECT 1881.880 573.430 1901.115 573.450 ;
        RECT 1881.880 573.150 1889.370 573.430 ;
        RECT 1900.785 573.415 1901.115 573.430 ;
        RECT 2100.000 557.670 2104.600 557.970 ;
        RECT 2083.865 556.730 2084.195 556.745 ;
        RECT 2100.670 556.730 2100.970 557.670 ;
        RECT 2083.865 556.430 2100.970 556.730 ;
        RECT 2083.865 556.415 2084.195 556.430 ;
      LAYER met3 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met3 ;
        RECT 2504.305 915.770 2504.635 915.785 ;
        RECT 2486.150 915.470 2504.635 915.770 ;
        RECT 2486.150 913.610 2486.450 915.470 ;
        RECT 2504.305 915.455 2504.635 915.470 ;
        RECT 2481.880 913.310 2486.480 913.610 ;
        RECT 2482.225 906.930 2482.555 906.945 ;
        RECT 2482.225 906.615 2482.770 906.930 ;
        RECT 2482.470 905.110 2482.770 906.615 ;
        RECT 2481.880 904.810 2486.480 905.110 ;
        RECT 2500.625 618.610 2500.955 618.625 ;
        RECT 2486.150 618.310 2500.955 618.610 ;
        RECT 2486.150 615.870 2486.450 618.310 ;
        RECT 2500.625 618.295 2500.955 618.310 ;
        RECT 2481.880 615.570 2486.480 615.870 ;
        RECT 2500.165 610.450 2500.495 610.465 ;
        RECT 2486.150 610.150 2500.495 610.450 ;
        RECT 2486.150 607.370 2486.450 610.150 ;
        RECT 2500.165 610.135 2500.495 610.150 ;
        RECT 2481.880 607.070 2486.480 607.370 ;
        RECT 2499.705 604.330 2500.035 604.345 ;
        RECT 2486.150 604.030 2500.035 604.330 ;
        RECT 2486.150 601.730 2486.450 604.030 ;
        RECT 2499.705 604.015 2500.035 604.030 ;
        RECT 2481.880 601.430 2486.480 601.730 ;
        RECT 2499.245 593.450 2499.575 593.465 ;
        RECT 2486.150 593.230 2499.575 593.450 ;
        RECT 2481.880 593.150 2499.575 593.230 ;
        RECT 2481.880 592.930 2486.480 593.150 ;
        RECT 2499.245 593.135 2499.575 593.150 ;
        RECT 2498.785 590.730 2499.115 590.745 ;
        RECT 2486.150 590.430 2499.115 590.730 ;
        RECT 2486.150 587.590 2486.450 590.430 ;
        RECT 2498.785 590.415 2499.115 590.430 ;
        RECT 2481.880 587.290 2486.480 587.590 ;
        RECT 2498.325 579.170 2498.655 579.185 ;
        RECT 2486.150 579.090 2498.655 579.170 ;
        RECT 2481.880 578.870 2498.655 579.090 ;
        RECT 2481.880 578.790 2486.480 578.870 ;
        RECT 2498.325 578.855 2498.655 578.870 ;
        RECT 2497.865 576.450 2498.195 576.465 ;
        RECT 2486.150 576.150 2498.195 576.450 ;
        RECT 2486.150 573.450 2486.450 576.150 ;
        RECT 2497.865 576.135 2498.195 576.150 ;
        RECT 2481.880 573.150 2486.480 573.450 ;
        RECT 1525.460 554.095 1527.200 555.000 ;
        RECT 2125.460 554.095 2127.200 555.000 ;
      LAYER via3 ;
        RECT 1867.900 3063.580 1868.220 3063.900 ;
        RECT 2442.900 3063.580 2443.220 3063.900 ;
        RECT 2469.580 3063.580 2469.900 3063.900 ;
        RECT 1845.820 3054.740 1846.140 3055.060 ;
        RECT 1865.140 3054.740 1865.460 3055.060 ;
        RECT 2139.840 2598.460 2140.160 2598.780 ;
        RECT 1568.900 2593.700 1569.220 2594.020 ;
        RECT 1573.500 2593.700 1573.820 2594.020 ;
        RECT 1580.860 2593.700 1581.180 2594.020 ;
        RECT 1590.980 2593.700 1591.300 2594.020 ;
        RECT 1598.340 2593.700 1598.660 2594.020 ;
        RECT 1603.860 2593.700 1604.180 2594.020 ;
        RECT 1614.900 2593.700 1615.220 2594.020 ;
        RECT 1622.260 2593.700 1622.580 2594.020 ;
        RECT 1626.860 2593.700 1627.180 2594.020 ;
        RECT 1650.780 2593.700 1651.100 2594.020 ;
        RECT 1661.820 2593.700 1662.140 2594.020 ;
        RECT 1671.020 2593.700 1671.340 2594.020 ;
        RECT 1690.340 2593.700 1690.660 2594.020 ;
        RECT 1696.780 2593.700 1697.100 2594.020 ;
        RECT 1738.180 2593.700 1738.500 2594.020 ;
        RECT 2215.660 2593.700 2215.980 2594.020 ;
        RECT 2256.140 2593.700 2256.460 2594.020 ;
        RECT 2262.580 2593.700 2262.900 2594.020 ;
        RECT 2268.100 2593.700 2268.420 2594.020 ;
        RECT 2302.140 2593.700 2302.460 2594.020 ;
        RECT 2305.820 2593.700 2306.140 2594.020 ;
        RECT 1582.700 2593.020 1583.020 2593.340 ;
        RECT 1587.300 2593.020 1587.620 2593.340 ;
        RECT 1638.820 2593.020 1639.140 2593.340 ;
        RECT 1644.340 2593.020 1644.660 2593.340 ;
        RECT 1656.300 2593.020 1656.620 2593.340 ;
        RECT 1679.300 2593.020 1679.620 2593.340 ;
        RECT 1707.820 2593.020 1708.140 2593.340 ;
        RECT 1732.660 2593.020 1732.980 2593.340 ;
        RECT 1743.700 2593.020 1744.020 2593.340 ;
        RECT 2148.500 2593.020 2148.820 2593.340 ;
        RECT 2220.260 2593.020 2220.580 2593.340 ;
        RECT 2292.020 2593.020 2292.340 2593.340 ;
        RECT 2297.540 2593.020 2297.860 2593.340 ;
        RECT 2312.260 2593.020 2312.580 2593.340 ;
        RECT 2337.100 2593.020 2337.420 2593.340 ;
        RECT 1562.460 2592.340 1562.780 2592.660 ;
        RECT 1575.340 2592.340 1575.660 2592.660 ;
        RECT 1608.460 2592.340 1608.780 2592.660 ;
        RECT 1621.340 2592.340 1621.660 2592.660 ;
        RECT 1633.300 2592.340 1633.620 2592.660 ;
        RECT 1667.340 2592.340 1667.660 2592.660 ;
        RECT 1685.740 2592.340 1686.060 2592.660 ;
        RECT 1702.300 2592.340 1702.620 2592.660 ;
        RECT 1725.300 2592.340 1725.620 2592.660 ;
        RECT 2154.020 2592.340 2154.340 2592.660 ;
        RECT 2238.660 2592.340 2238.980 2592.660 ;
        RECT 2249.700 2592.340 2250.020 2592.660 ;
        RECT 2280.060 2592.340 2280.380 2592.660 ;
        RECT 2285.580 2592.340 2285.900 2592.660 ;
        RECT 2342.620 2592.340 2342.940 2592.660 ;
        RECT 1610.300 2591.660 1610.620 2591.980 ;
        RECT 1715.180 2591.660 1715.500 2591.980 ;
        RECT 1718.860 2591.660 1719.180 2591.980 ;
        RECT 2145.740 2591.660 2146.060 2591.980 ;
        RECT 2233.140 2591.660 2233.460 2591.980 ;
        RECT 2244.180 2591.660 2244.500 2591.980 ;
        RECT 2273.620 2591.660 2273.940 2591.980 ;
        RECT 2319.620 2591.660 2319.940 2591.980 ;
        RECT 2332.500 2591.660 2332.820 2591.980 ;
        RECT 1586.380 2590.980 1586.700 2591.300 ;
        RECT 1616.740 2590.980 1617.060 2591.300 ;
        RECT 2209.220 2590.980 2209.540 2591.300 ;
        RECT 2226.700 2590.980 2227.020 2591.300 ;
        RECT 2326.060 2590.980 2326.380 2591.300 ;
        RECT 1599.260 2590.300 1599.580 2590.620 ;
        RECT 1657.220 2590.300 1657.540 2590.620 ;
        RECT 1680.220 2590.300 1680.540 2590.620 ;
        RECT 2132.860 2590.300 2133.180 2590.620 ;
        RECT 2175.180 2590.300 2175.500 2590.620 ;
        RECT 2180.700 2590.300 2181.020 2590.620 ;
        RECT 1569.820 2589.620 1570.140 2589.940 ;
        RECT 1592.820 2589.620 1593.140 2589.940 ;
        RECT 1604.780 2589.620 1605.100 2589.940 ;
        RECT 1645.260 2589.620 1645.580 2589.940 ;
        RECT 1663.660 2589.620 1663.980 2589.940 ;
        RECT 2186.220 2589.620 2186.540 2589.940 ;
        RECT 1634.220 2588.940 1634.540 2589.260 ;
        RECT 1686.660 2588.940 1686.980 2589.260 ;
        RECT 1692.180 2588.940 1692.500 2589.260 ;
        RECT 2168.740 2588.940 2169.060 2589.260 ;
        RECT 1551.420 2588.260 1551.740 2588.580 ;
        RECT 1563.380 2588.260 1563.700 2588.580 ;
        RECT 1627.780 2588.260 1628.100 2588.580 ;
        RECT 1639.740 2588.260 1640.060 2588.580 ;
        RECT 1669.180 2588.260 1669.500 2588.580 ;
        RECT 1674.700 2588.260 1675.020 2588.580 ;
        RECT 1697.700 2588.260 1698.020 2588.580 ;
        RECT 1741.860 2588.260 1742.180 2588.580 ;
        RECT 2163.220 2588.260 2163.540 2588.580 ;
        RECT 2165.060 2588.260 2165.380 2588.580 ;
        RECT 2169.660 2588.260 2169.980 2588.580 ;
        RECT 2178.860 2588.260 2179.180 2588.580 ;
        RECT 2184.380 2588.260 2184.700 2588.580 ;
        RECT 2189.900 2588.260 2190.220 2588.580 ;
        RECT 2198.180 2588.260 2198.500 2588.580 ;
        RECT 2203.700 2588.260 2204.020 2588.580 ;
        RECT 2224.860 2588.260 2225.180 2588.580 ;
        RECT 2266.260 2588.260 2266.580 2588.580 ;
        RECT 2301.220 2588.260 2301.540 2588.580 ;
        RECT 2341.700 2588.260 2342.020 2588.580 ;
        RECT 1536.700 2587.580 1537.020 2587.900 ;
        RECT 1543.140 2587.580 1543.460 2587.900 ;
        RECT 1548.660 2587.580 1548.980 2587.900 ;
        RECT 1558.780 2587.580 1559.100 2587.900 ;
        RECT 1651.700 2587.580 1652.020 2587.900 ;
        RECT 1703.220 2587.580 1703.540 2587.900 ;
        RECT 1709.660 2587.580 1709.980 2587.900 ;
        RECT 1717.020 2587.580 1717.340 2587.900 ;
        RECT 1721.620 2587.580 1721.940 2587.900 ;
        RECT 1729.900 2587.580 1730.220 2587.900 ;
        RECT 1736.340 2587.580 1736.660 2587.900 ;
        RECT 1744.620 2587.580 1744.940 2587.900 ;
        RECT 2191.740 2587.580 2192.060 2587.900 ;
        RECT 2193.580 2587.580 2193.900 2587.900 ;
        RECT 2200.020 2587.580 2200.340 2587.900 ;
        RECT 2207.380 2587.580 2207.700 2587.900 ;
        RECT 2213.820 2587.580 2214.140 2587.900 ;
        RECT 2219.340 2587.580 2219.660 2587.900 ;
        RECT 2227.620 2587.580 2227.940 2587.900 ;
        RECT 2234.980 2587.580 2235.300 2587.900 ;
        RECT 2241.420 2587.580 2241.740 2587.900 ;
        RECT 2248.780 2587.580 2249.100 2587.900 ;
        RECT 2254.300 2587.580 2254.620 2587.900 ;
        RECT 2259.820 2587.580 2260.140 2587.900 ;
        RECT 2269.020 2587.580 2269.340 2587.900 ;
        RECT 2276.380 2587.580 2276.700 2587.900 ;
        RECT 2281.900 2587.580 2282.220 2587.900 ;
        RECT 2289.260 2587.580 2289.580 2587.900 ;
        RECT 2295.700 2587.580 2296.020 2587.900 ;
        RECT 2303.980 2587.580 2304.300 2587.900 ;
        RECT 2310.420 2587.580 2310.740 2587.900 ;
        RECT 2317.780 2587.580 2318.100 2587.900 ;
        RECT 2324.220 2587.580 2324.540 2587.900 ;
        RECT 2330.660 2587.580 2330.980 2587.900 ;
        RECT 2336.180 2587.580 2336.500 2587.900 ;
        RECT 2345.380 2587.580 2345.700 2587.900 ;
        RECT 1647.100 1062.340 1647.420 1062.660 ;
        RECT 1682.060 1038.540 1682.380 1038.860 ;
        RECT 1704.140 1020.860 1704.460 1021.180 ;
        RECT 1786.940 1019.500 1787.260 1019.820 ;
        RECT 1834.780 1020.860 1835.100 1021.180 ;
        RECT 1843.980 1020.860 1844.300 1021.180 ;
        RECT 1855.020 1020.860 1855.340 1021.180 ;
        RECT 2241.420 1020.860 2241.740 1021.180 ;
        RECT 2260.740 1020.860 2261.060 1021.180 ;
        RECT 2266.260 1020.860 2266.580 1021.180 ;
        RECT 2270.860 1020.860 2271.180 1021.180 ;
        RECT 2281.900 1020.860 2282.220 1021.180 ;
        RECT 2328.820 1020.860 2329.140 1021.180 ;
        RECT 2333.420 1020.860 2333.740 1021.180 ;
        RECT 2340.780 1020.860 2341.100 1021.180 ;
        RECT 2351.820 1020.860 2352.140 1021.180 ;
        RECT 2358.260 1020.860 2358.580 1021.180 ;
        RECT 2373.900 1020.860 2374.220 1021.180 ;
        RECT 2403.340 1020.860 2403.660 1021.180 ;
        RECT 2421.740 1020.860 2422.060 1021.180 ;
        RECT 1837.540 1020.180 1837.860 1020.500 ;
        RECT 2247.860 1020.180 2248.180 1020.500 ;
        RECT 2254.300 1020.180 2254.620 1020.500 ;
        RECT 2282.820 1020.180 2283.140 1020.500 ;
        RECT 2346.300 1020.180 2346.620 1020.500 ;
        RECT 2361.020 1020.180 2361.340 1020.500 ;
        RECT 2381.260 1020.180 2381.580 1020.500 ;
        RECT 2387.700 1020.180 2388.020 1020.500 ;
        RECT 2451.180 1020.180 2451.500 1020.500 ;
        RECT 1801.660 1019.500 1801.980 1019.820 ;
        RECT 1832.020 1019.500 1832.340 1019.820 ;
        RECT 2272.700 1019.500 2273.020 1019.820 ;
        RECT 2276.380 1019.500 2276.700 1019.820 ;
        RECT 1808.100 1018.820 1808.420 1019.140 ;
        RECT 2429.100 1018.820 2429.420 1019.140 ;
        RECT 1711.500 1018.140 1711.820 1018.460 ;
        RECT 1719.780 1018.140 1720.100 1018.460 ;
        RECT 1745.540 1018.140 1745.860 1018.460 ;
        RECT 1763.940 1018.140 1764.260 1018.460 ;
        RECT 1774.060 1018.140 1774.380 1018.460 ;
        RECT 1714.260 1017.460 1714.580 1017.780 ;
        RECT 1641.580 1016.780 1641.900 1017.100 ;
        RECT 1654.460 1016.780 1654.780 1017.100 ;
        RECT 1671.020 1016.780 1671.340 1017.100 ;
        RECT 1684.820 1016.780 1685.140 1017.100 ;
        RECT 1814.540 1016.780 1814.860 1017.100 ;
        RECT 1821.900 1016.780 1822.220 1017.100 ;
        RECT 2264.420 1016.780 2264.740 1017.100 ;
        RECT 2280.060 1016.780 2280.380 1017.100 ;
        RECT 2300.300 1016.780 2300.620 1017.100 ;
        RECT 2311.340 1016.780 2311.660 1017.100 ;
        RECT 2393.220 1016.780 2393.540 1017.100 ;
        RECT 2395.980 1016.780 2396.300 1017.100 ;
        RECT 1640.660 1016.100 1640.980 1016.420 ;
        RECT 1653.540 1016.100 1653.860 1016.420 ;
        RECT 1658.140 1016.100 1658.460 1016.420 ;
        RECT 1664.580 1016.100 1664.900 1016.420 ;
        RECT 1675.620 1016.100 1675.940 1016.420 ;
        RECT 1692.180 1016.100 1692.500 1016.420 ;
        RECT 1698.620 1016.100 1698.940 1016.420 ;
        RECT 1726.220 1016.100 1726.540 1016.420 ;
        RECT 1732.660 1016.100 1732.980 1016.420 ;
        RECT 1749.220 1016.100 1749.540 1016.420 ;
        RECT 1780.500 1016.100 1780.820 1016.420 ;
        RECT 2289.260 1016.100 2289.580 1016.420 ;
        RECT 2293.860 1016.100 2294.180 1016.420 ;
        RECT 2304.900 1016.100 2305.220 1016.420 ;
        RECT 2315.940 1016.100 2316.260 1016.420 ;
        RECT 2322.380 1016.100 2322.700 1016.420 ;
        RECT 2359.180 1016.100 2359.500 1016.420 ;
        RECT 2390.460 1016.100 2390.780 1016.420 ;
        RECT 2408.860 1018.140 2409.180 1018.460 ;
        RECT 2431.860 1018.140 2432.180 1018.460 ;
        RECT 2410.700 1017.460 2411.020 1017.780 ;
        RECT 2437.380 1017.460 2437.700 1017.780 ;
        RECT 2415.300 1016.780 2415.620 1017.100 ;
        RECT 2423.580 1016.780 2423.900 1017.100 ;
        RECT 2442.900 1016.100 2443.220 1016.420 ;
        RECT 1661.820 1015.420 1662.140 1015.740 ;
        RECT 1668.260 1015.420 1668.580 1015.740 ;
        RECT 1673.780 1015.420 1674.100 1015.740 ;
        RECT 1682.980 1015.420 1683.300 1015.740 ;
        RECT 1739.100 1015.420 1739.420 1015.740 ;
        RECT 1755.660 1015.420 1755.980 1015.740 ;
        RECT 1766.700 1015.420 1767.020 1015.740 ;
        RECT 1788.780 1015.420 1789.100 1015.740 ;
        RECT 1648.020 1014.740 1648.340 1015.060 ;
        RECT 1680.220 1014.740 1680.540 1015.060 ;
        RECT 1689.420 1014.740 1689.740 1015.060 ;
        RECT 1695.860 1014.740 1696.180 1015.060 ;
        RECT 1700.460 1014.740 1700.780 1015.060 ;
        RECT 1706.900 1014.740 1707.220 1015.060 ;
        RECT 1713.340 1014.740 1713.660 1015.060 ;
        RECT 1717.940 1014.740 1718.260 1015.060 ;
        RECT 1724.380 1014.740 1724.700 1015.060 ;
        RECT 1730.820 1014.740 1731.140 1015.060 ;
        RECT 1735.420 1014.740 1735.740 1015.060 ;
        RECT 1741.860 1014.740 1742.180 1015.060 ;
        RECT 1748.300 1014.740 1748.620 1015.060 ;
        RECT 1754.740 1014.740 1755.060 1015.060 ;
        RECT 1758.420 1014.740 1758.740 1015.060 ;
        RECT 1765.780 1014.740 1766.100 1015.060 ;
        RECT 1772.220 1014.740 1772.540 1015.060 ;
        RECT 1777.740 1014.740 1778.060 1015.060 ;
        RECT 1782.340 1014.740 1782.660 1015.060 ;
        RECT 1789.700 1014.740 1790.020 1015.060 ;
        RECT 1793.380 1014.740 1793.700 1015.060 ;
        RECT 1796.140 1014.740 1796.460 1015.060 ;
        RECT 1799.820 1014.740 1800.140 1015.060 ;
        RECT 1806.260 1014.740 1806.580 1015.060 ;
        RECT 1812.700 1014.740 1813.020 1015.060 ;
        RECT 1817.300 1014.740 1817.620 1015.060 ;
        RECT 1823.740 1014.740 1824.060 1015.060 ;
        RECT 2246.940 1014.740 2247.260 1015.060 ;
        RECT 2253.380 1014.740 2253.700 1015.060 ;
        RECT 2258.900 1014.740 2259.220 1015.060 ;
        RECT 2287.420 1014.740 2287.740 1015.060 ;
        RECT 2294.780 1014.740 2295.100 1015.060 ;
        RECT 2303.060 1014.740 2303.380 1015.060 ;
        RECT 2307.660 1014.740 2307.980 1015.060 ;
        RECT 2312.260 1014.740 2312.580 1015.060 ;
        RECT 2317.780 1014.740 2318.100 1015.060 ;
        RECT 2323.300 1014.740 2323.620 1015.060 ;
        RECT 2329.740 1014.740 2330.060 1015.060 ;
        RECT 2335.260 1014.740 2335.580 1015.060 ;
        RECT 2342.620 1014.740 2342.940 1015.060 ;
        RECT 2347.220 1014.740 2347.540 1015.060 ;
        RECT 2355.500 1014.740 2355.820 1015.060 ;
        RECT 2364.700 1014.740 2365.020 1015.060 ;
        RECT 2367.460 1014.740 2367.780 1015.060 ;
        RECT 2372.980 1014.740 2373.300 1015.060 ;
        RECT 2377.580 1014.740 2377.900 1015.060 ;
        RECT 2382.180 1014.740 2382.500 1015.060 ;
        RECT 2388.620 1014.740 2388.940 1015.060 ;
        RECT 2399.660 1014.740 2399.980 1015.060 ;
        RECT 2406.100 1014.740 2406.420 1015.060 ;
        RECT 2417.140 1014.740 2417.460 1015.060 ;
        RECT 2241.920 1006.580 2242.240 1006.900 ;
      LAYER met4 ;
        RECT 1867.895 3063.575 1868.225 3063.905 ;
        RECT 2442.895 3063.575 2443.225 3063.905 ;
        RECT 2469.575 3063.575 2469.905 3063.905 ;
        RECT 1867.910 3056.235 1868.210 3063.575 ;
        RECT 2442.910 3056.235 2443.210 3063.575 ;
        RECT 1594.025 3051.635 1594.325 3056.235 ;
        RECT 1600.265 3051.635 1600.565 3056.235 ;
        RECT 1606.505 3051.635 1606.805 3056.235 ;
        RECT 1612.745 3051.635 1613.045 3056.235 ;
        RECT 1618.985 3051.635 1619.285 3056.235 ;
        RECT 1625.225 3051.635 1625.525 3056.235 ;
        RECT 1631.465 3051.635 1631.765 3056.235 ;
        RECT 1637.705 3051.635 1638.005 3056.235 ;
        RECT 1643.945 3051.635 1644.245 3056.235 ;
        RECT 1650.185 3051.635 1650.485 3056.235 ;
        RECT 1656.425 3051.635 1656.725 3056.235 ;
        RECT 1662.665 3051.635 1662.965 3056.235 ;
        RECT 1668.905 3051.635 1669.205 3056.235 ;
        RECT 1675.145 3051.635 1675.445 3056.235 ;
        RECT 1681.385 3051.635 1681.685 3056.235 ;
        RECT 1687.625 3051.635 1687.925 3056.235 ;
        RECT 1693.865 3051.635 1694.165 3056.235 ;
        RECT 1700.105 3051.635 1700.405 3056.235 ;
        RECT 1706.345 3051.635 1706.645 3056.235 ;
        RECT 1712.585 3051.635 1712.885 3056.235 ;
        RECT 1718.825 3051.635 1719.125 3056.235 ;
        RECT 1725.065 3051.635 1725.365 3056.235 ;
        RECT 1731.305 3051.635 1731.605 3056.235 ;
        RECT 1737.545 3051.635 1737.845 3056.235 ;
        RECT 1743.785 3051.635 1744.085 3056.235 ;
        RECT 1750.025 3051.635 1750.325 3056.235 ;
        RECT 1756.265 3051.635 1756.565 3056.235 ;
        RECT 1762.505 3051.635 1762.805 3056.235 ;
        RECT 1768.745 3051.635 1769.045 3056.235 ;
        RECT 1774.985 3051.635 1775.285 3056.235 ;
        RECT 1781.225 3051.635 1781.525 3056.235 ;
        RECT 1787.465 3051.635 1787.765 3056.235 ;
        RECT 1842.890 3055.050 1843.190 3056.235 ;
        RECT 1845.815 3055.050 1846.145 3055.065 ;
        RECT 1842.890 3054.750 1846.145 3055.050 ;
        RECT 1842.890 3051.635 1843.190 3054.750 ;
        RECT 1845.815 3054.735 1846.145 3054.750 ;
        RECT 1865.135 3055.050 1865.465 3055.065 ;
        RECT 1867.865 3055.050 1868.210 3056.235 ;
        RECT 1865.135 3054.750 1868.210 3055.050 ;
        RECT 1865.135 3054.735 1865.465 3054.750 ;
        RECT 1867.865 3051.635 1868.165 3054.750 ;
        RECT 2194.025 3051.635 2194.325 3056.235 ;
        RECT 2200.265 3051.635 2200.565 3056.235 ;
        RECT 2206.505 3051.635 2206.805 3056.235 ;
        RECT 2212.745 3051.635 2213.045 3056.235 ;
        RECT 2218.985 3051.635 2219.285 3056.235 ;
        RECT 2225.225 3051.635 2225.525 3056.235 ;
        RECT 2231.465 3051.635 2231.765 3056.235 ;
        RECT 2237.705 3051.635 2238.005 3056.235 ;
        RECT 2243.945 3051.635 2244.245 3056.235 ;
        RECT 2250.185 3051.635 2250.485 3056.235 ;
        RECT 2256.425 3051.635 2256.725 3056.235 ;
        RECT 2262.665 3051.635 2262.965 3056.235 ;
        RECT 2268.905 3051.635 2269.205 3056.235 ;
        RECT 2275.145 3051.635 2275.445 3056.235 ;
        RECT 2281.385 3051.635 2281.685 3056.235 ;
        RECT 2287.625 3051.635 2287.925 3056.235 ;
        RECT 2293.865 3051.635 2294.165 3056.235 ;
        RECT 2300.105 3051.635 2300.405 3056.235 ;
        RECT 2306.345 3051.635 2306.645 3056.235 ;
        RECT 2312.585 3051.635 2312.885 3056.235 ;
        RECT 2318.825 3051.635 2319.125 3056.235 ;
        RECT 2325.065 3051.635 2325.365 3056.235 ;
        RECT 2331.305 3051.635 2331.605 3056.235 ;
        RECT 2337.545 3051.635 2337.845 3056.235 ;
        RECT 2343.785 3051.635 2344.085 3056.235 ;
        RECT 2350.025 3051.635 2350.325 3056.235 ;
        RECT 2356.265 3051.635 2356.565 3056.235 ;
        RECT 2362.505 3051.635 2362.805 3056.235 ;
        RECT 2368.745 3051.635 2369.045 3056.235 ;
        RECT 2374.985 3051.635 2375.285 3056.235 ;
        RECT 2381.225 3051.635 2381.525 3056.235 ;
        RECT 2387.465 3051.635 2387.765 3056.235 ;
        RECT 2442.890 3054.750 2443.210 3056.235 ;
        RECT 2467.865 3055.050 2468.165 3056.235 ;
        RECT 2469.590 3055.050 2469.890 3063.575 ;
        RECT 2467.865 3054.750 2469.890 3055.050 ;
        RECT 2442.890 3051.635 2443.190 3054.750 ;
        RECT 2467.865 3051.635 2468.165 3054.750 ;
      LAYER met4 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
      LAYER met4 ;
        RECT 1534.010 2601.150 1534.310 2604.600 ;
        RECT 1539.850 2601.150 1540.150 2604.600 ;
        RECT 1545.690 2601.150 1545.990 2604.600 ;
        RECT 1551.530 2601.150 1551.830 2604.600 ;
        RECT 1534.010 2600.850 1537.010 2601.150 ;
        RECT 1534.010 2600.000 1534.310 2600.850 ;
        RECT 1536.710 2587.905 1537.010 2600.850 ;
        RECT 1539.850 2600.850 1543.450 2601.150 ;
        RECT 1539.850 2600.000 1540.150 2600.850 ;
        RECT 1543.150 2587.905 1543.450 2600.850 ;
        RECT 1545.690 2600.850 1548.970 2601.150 ;
        RECT 1545.690 2600.000 1545.990 2600.850 ;
        RECT 1548.670 2587.905 1548.970 2600.850 ;
        RECT 1551.430 2600.000 1551.830 2601.150 ;
        RECT 1557.370 2601.150 1557.670 2604.600 ;
        RECT 1563.210 2601.150 1563.510 2604.600 ;
        RECT 1557.370 2600.850 1559.090 2601.150 ;
        RECT 1557.370 2600.000 1557.670 2600.850 ;
        RECT 1551.430 2588.585 1551.730 2600.000 ;
        RECT 1551.415 2588.255 1551.745 2588.585 ;
        RECT 1558.790 2587.905 1559.090 2600.850 ;
        RECT 1562.470 2600.850 1563.510 2601.150 ;
        RECT 1562.470 2592.665 1562.770 2600.850 ;
        RECT 1563.210 2600.000 1563.510 2600.850 ;
        RECT 1563.830 2599.450 1564.130 2604.600 ;
        RECT 1569.050 2601.150 1569.350 2604.600 ;
        RECT 1563.390 2599.150 1564.130 2599.450 ;
        RECT 1568.910 2600.000 1569.350 2601.150 ;
        RECT 1569.670 2601.150 1569.970 2604.600 ;
        RECT 1574.890 2602.850 1575.190 2604.600 ;
        RECT 1573.510 2602.550 1575.190 2602.850 ;
        RECT 1569.670 2600.000 1570.130 2601.150 ;
        RECT 1562.455 2592.335 1562.785 2592.665 ;
        RECT 1563.390 2588.585 1563.690 2599.150 ;
        RECT 1568.910 2594.025 1569.210 2600.000 ;
        RECT 1568.895 2593.695 1569.225 2594.025 ;
        RECT 1569.830 2589.945 1570.130 2600.000 ;
        RECT 1573.510 2594.025 1573.810 2602.550 ;
        RECT 1574.890 2600.000 1575.190 2602.550 ;
        RECT 1575.510 2599.450 1575.810 2604.600 ;
        RECT 1575.350 2599.150 1575.810 2599.450 ;
        RECT 1580.730 2599.450 1581.030 2604.600 ;
        RECT 1581.350 2602.850 1581.650 2604.600 ;
        RECT 1581.350 2602.550 1583.010 2602.850 ;
        RECT 1581.350 2600.000 1581.650 2602.550 ;
        RECT 1580.730 2599.150 1581.170 2599.450 ;
        RECT 1573.495 2593.695 1573.825 2594.025 ;
        RECT 1575.350 2592.665 1575.650 2599.150 ;
        RECT 1580.870 2594.025 1581.170 2599.150 ;
        RECT 1580.855 2593.695 1581.185 2594.025 ;
        RECT 1582.710 2593.345 1583.010 2602.550 ;
        RECT 1586.570 2601.150 1586.870 2604.600 ;
        RECT 1586.390 2600.000 1586.870 2601.150 ;
        RECT 1587.190 2601.150 1587.490 2604.600 ;
        RECT 1592.410 2602.850 1592.710 2604.600 ;
        RECT 1590.990 2602.550 1592.710 2602.850 ;
        RECT 1587.190 2600.000 1587.610 2601.150 ;
        RECT 1582.695 2593.015 1583.025 2593.345 ;
        RECT 1575.335 2592.335 1575.665 2592.665 ;
        RECT 1586.390 2591.305 1586.690 2600.000 ;
        RECT 1587.310 2593.345 1587.610 2600.000 ;
        RECT 1590.990 2594.025 1591.290 2602.550 ;
        RECT 1592.410 2600.000 1592.710 2602.550 ;
        RECT 1593.030 2599.450 1593.330 2604.600 ;
        RECT 1592.830 2599.150 1593.330 2599.450 ;
        RECT 1590.975 2593.695 1591.305 2594.025 ;
        RECT 1587.295 2593.015 1587.625 2593.345 ;
        RECT 1586.375 2590.975 1586.705 2591.305 ;
        RECT 1592.830 2589.945 1593.130 2599.150 ;
        RECT 1598.250 2596.050 1598.550 2604.600 ;
        RECT 1598.870 2599.450 1599.170 2604.600 ;
        RECT 1604.090 2601.150 1604.390 2604.600 ;
        RECT 1603.870 2600.000 1604.390 2601.150 ;
        RECT 1604.710 2601.150 1605.010 2604.600 ;
        RECT 1609.930 2602.850 1610.230 2604.600 ;
        RECT 1608.470 2602.550 1610.230 2602.850 ;
        RECT 1604.710 2600.000 1605.090 2601.150 ;
        RECT 1598.870 2599.150 1599.570 2599.450 ;
        RECT 1598.250 2595.750 1598.650 2596.050 ;
        RECT 1598.350 2594.025 1598.650 2595.750 ;
        RECT 1598.335 2593.695 1598.665 2594.025 ;
        RECT 1599.270 2590.625 1599.570 2599.150 ;
        RECT 1603.870 2594.025 1604.170 2600.000 ;
        RECT 1603.855 2593.695 1604.185 2594.025 ;
        RECT 1599.255 2590.295 1599.585 2590.625 ;
        RECT 1604.790 2589.945 1605.090 2600.000 ;
        RECT 1608.470 2592.665 1608.770 2602.550 ;
        RECT 1609.930 2600.000 1610.230 2602.550 ;
        RECT 1610.550 2599.450 1610.850 2604.600 ;
        RECT 1615.770 2601.150 1616.070 2604.600 ;
        RECT 1610.310 2599.150 1610.850 2599.450 ;
        RECT 1614.910 2600.850 1616.070 2601.150 ;
        RECT 1608.455 2592.335 1608.785 2592.665 ;
        RECT 1610.310 2591.985 1610.610 2599.150 ;
        RECT 1614.910 2594.025 1615.210 2600.850 ;
        RECT 1615.770 2600.000 1616.070 2600.850 ;
        RECT 1616.390 2599.450 1616.690 2604.600 ;
        RECT 1621.610 2601.150 1621.910 2604.600 ;
        RECT 1621.350 2600.000 1621.910 2601.150 ;
        RECT 1622.230 2601.150 1622.530 2604.600 ;
        RECT 1627.450 2602.850 1627.750 2604.600 ;
        RECT 1625.950 2602.550 1627.750 2602.850 ;
        RECT 1622.230 2600.000 1622.570 2601.150 ;
        RECT 1616.390 2599.150 1617.050 2599.450 ;
        RECT 1614.895 2593.695 1615.225 2594.025 ;
        RECT 1610.295 2591.655 1610.625 2591.985 ;
        RECT 1616.750 2591.305 1617.050 2599.150 ;
        RECT 1621.350 2592.665 1621.650 2600.000 ;
        RECT 1622.270 2594.025 1622.570 2600.000 ;
        RECT 1625.950 2599.450 1626.250 2602.550 ;
        RECT 1627.450 2600.000 1627.750 2602.550 ;
        RECT 1628.070 2599.450 1628.370 2604.600 ;
        RECT 1625.950 2599.150 1627.170 2599.450 ;
        RECT 1626.870 2594.025 1627.170 2599.150 ;
        RECT 1627.790 2599.150 1628.370 2599.450 ;
        RECT 1633.290 2599.450 1633.590 2604.600 ;
        RECT 1633.910 2599.450 1634.210 2604.600 ;
        RECT 1639.130 2601.150 1639.430 2604.600 ;
        RECT 1638.830 2600.000 1639.430 2601.150 ;
        RECT 1633.290 2599.150 1633.610 2599.450 ;
        RECT 1633.910 2599.150 1634.530 2599.450 ;
        RECT 1622.255 2593.695 1622.585 2594.025 ;
        RECT 1626.855 2593.695 1627.185 2594.025 ;
        RECT 1621.335 2592.335 1621.665 2592.665 ;
        RECT 1616.735 2590.975 1617.065 2591.305 ;
        RECT 1569.815 2589.615 1570.145 2589.945 ;
        RECT 1592.815 2589.615 1593.145 2589.945 ;
        RECT 1604.775 2589.615 1605.105 2589.945 ;
        RECT 1627.790 2588.585 1628.090 2599.150 ;
        RECT 1633.310 2592.665 1633.610 2599.150 ;
        RECT 1633.295 2592.335 1633.625 2592.665 ;
        RECT 1634.230 2589.265 1634.530 2599.150 ;
        RECT 1638.830 2593.345 1639.130 2600.000 ;
        RECT 1638.815 2593.015 1639.145 2593.345 ;
        RECT 1634.215 2588.935 1634.545 2589.265 ;
        RECT 1639.750 2588.585 1640.050 2604.600 ;
        RECT 1644.970 2601.150 1645.270 2604.600 ;
        RECT 1644.350 2600.850 1645.270 2601.150 ;
        RECT 1644.350 2593.345 1644.650 2600.850 ;
        RECT 1644.970 2600.000 1645.270 2600.850 ;
        RECT 1645.590 2599.450 1645.890 2604.600 ;
        RECT 1650.810 2601.150 1651.110 2604.600 ;
        RECT 1645.270 2599.150 1645.890 2599.450 ;
        RECT 1650.790 2600.000 1651.110 2601.150 ;
        RECT 1651.430 2601.150 1651.730 2604.600 ;
        RECT 1656.650 2601.150 1656.950 2604.600 ;
        RECT 1651.430 2600.000 1652.010 2601.150 ;
        RECT 1644.335 2593.015 1644.665 2593.345 ;
        RECT 1645.270 2589.945 1645.570 2599.150 ;
        RECT 1650.790 2594.025 1651.090 2600.000 ;
        RECT 1650.775 2593.695 1651.105 2594.025 ;
        RECT 1645.255 2589.615 1645.585 2589.945 ;
        RECT 1563.375 2588.255 1563.705 2588.585 ;
        RECT 1627.775 2588.255 1628.105 2588.585 ;
        RECT 1639.735 2588.255 1640.065 2588.585 ;
        RECT 1651.710 2587.905 1652.010 2600.000 ;
        RECT 1656.540 2600.000 1656.950 2601.150 ;
        RECT 1656.540 2599.450 1656.840 2600.000 ;
        RECT 1657.270 2599.450 1657.570 2604.600 ;
        RECT 1662.490 2601.150 1662.790 2604.600 ;
        RECT 1656.310 2599.150 1656.840 2599.450 ;
        RECT 1657.230 2599.150 1657.570 2599.450 ;
        RECT 1661.830 2600.850 1662.790 2601.150 ;
        RECT 1656.310 2593.345 1656.610 2599.150 ;
        RECT 1656.295 2593.015 1656.625 2593.345 ;
        RECT 1657.230 2590.625 1657.530 2599.150 ;
        RECT 1661.830 2594.025 1662.130 2600.850 ;
        RECT 1662.490 2600.000 1662.790 2600.850 ;
        RECT 1663.110 2599.450 1663.410 2604.600 ;
        RECT 1668.330 2601.150 1668.630 2604.600 ;
        RECT 1667.350 2600.850 1668.630 2601.150 ;
        RECT 1663.110 2599.150 1663.970 2599.450 ;
        RECT 1661.815 2593.695 1662.145 2594.025 ;
        RECT 1657.215 2590.295 1657.545 2590.625 ;
        RECT 1663.670 2589.945 1663.970 2599.150 ;
        RECT 1667.350 2592.665 1667.650 2600.850 ;
        RECT 1668.330 2600.000 1668.630 2600.850 ;
        RECT 1668.950 2601.150 1669.250 2604.600 ;
        RECT 1674.170 2601.150 1674.470 2604.600 ;
        RECT 1668.950 2600.000 1669.490 2601.150 ;
        RECT 1667.335 2592.335 1667.665 2592.665 ;
        RECT 1663.655 2589.615 1663.985 2589.945 ;
        RECT 1669.190 2588.585 1669.490 2600.000 ;
        RECT 1671.030 2600.850 1674.470 2601.150 ;
        RECT 1671.030 2594.025 1671.330 2600.850 ;
        RECT 1674.170 2600.000 1674.470 2600.850 ;
        RECT 1674.790 2599.450 1675.090 2604.600 ;
        RECT 1680.010 2601.150 1680.310 2604.600 ;
        RECT 1674.710 2599.150 1675.090 2599.450 ;
        RECT 1679.310 2600.850 1680.310 2601.150 ;
        RECT 1671.015 2593.695 1671.345 2594.025 ;
        RECT 1674.710 2588.585 1675.010 2599.150 ;
        RECT 1679.310 2593.345 1679.610 2600.850 ;
        RECT 1680.010 2600.000 1680.310 2600.850 ;
        RECT 1680.630 2599.450 1680.930 2604.600 ;
        RECT 1685.850 2601.150 1686.150 2604.600 ;
        RECT 1680.230 2599.150 1680.930 2599.450 ;
        RECT 1685.750 2600.000 1686.150 2601.150 ;
        RECT 1686.470 2601.150 1686.770 2604.600 ;
        RECT 1691.690 2602.850 1691.990 2604.600 ;
        RECT 1690.350 2602.550 1691.990 2602.850 ;
        RECT 1686.470 2600.000 1686.970 2601.150 ;
        RECT 1679.295 2593.015 1679.625 2593.345 ;
        RECT 1680.230 2590.625 1680.530 2599.150 ;
        RECT 1685.750 2592.665 1686.050 2600.000 ;
        RECT 1685.735 2592.335 1686.065 2592.665 ;
        RECT 1680.215 2590.295 1680.545 2590.625 ;
        RECT 1686.670 2589.265 1686.970 2600.000 ;
        RECT 1690.350 2594.025 1690.650 2602.550 ;
        RECT 1691.690 2600.000 1691.990 2602.550 ;
        RECT 1692.310 2599.450 1692.610 2604.600 ;
        RECT 1697.530 2601.150 1697.830 2604.600 ;
        RECT 1692.190 2599.150 1692.610 2599.450 ;
        RECT 1696.790 2600.850 1697.830 2601.150 ;
        RECT 1690.335 2593.695 1690.665 2594.025 ;
        RECT 1692.190 2589.265 1692.490 2599.150 ;
        RECT 1696.790 2594.025 1697.090 2600.850 ;
        RECT 1697.530 2600.000 1697.830 2600.850 ;
        RECT 1698.150 2599.450 1698.450 2604.600 ;
        RECT 1703.370 2601.150 1703.670 2604.600 ;
        RECT 1697.710 2599.150 1698.450 2599.450 ;
        RECT 1702.310 2600.850 1703.670 2601.150 ;
        RECT 1696.775 2593.695 1697.105 2594.025 ;
        RECT 1686.655 2588.935 1686.985 2589.265 ;
        RECT 1692.175 2588.935 1692.505 2589.265 ;
        RECT 1697.710 2588.585 1698.010 2599.150 ;
        RECT 1702.310 2592.665 1702.610 2600.850 ;
        RECT 1703.370 2600.000 1703.670 2600.850 ;
        RECT 1703.990 2599.450 1704.290 2604.600 ;
        RECT 1709.210 2602.850 1709.510 2604.600 ;
        RECT 1703.230 2599.150 1704.290 2599.450 ;
        RECT 1707.830 2602.550 1709.510 2602.850 ;
        RECT 1702.295 2592.335 1702.625 2592.665 ;
        RECT 1669.175 2588.255 1669.505 2588.585 ;
        RECT 1674.695 2588.255 1675.025 2588.585 ;
        RECT 1697.695 2588.255 1698.025 2588.585 ;
        RECT 1703.230 2587.905 1703.530 2599.150 ;
        RECT 1707.830 2593.345 1708.130 2602.550 ;
        RECT 1709.210 2600.000 1709.510 2602.550 ;
        RECT 1709.830 2599.450 1710.130 2604.600 ;
        RECT 1709.670 2599.150 1710.130 2599.450 ;
        RECT 1715.050 2599.450 1715.350 2604.600 ;
        RECT 1715.670 2602.850 1715.970 2604.600 ;
        RECT 1715.670 2602.550 1717.330 2602.850 ;
        RECT 1715.670 2600.000 1715.970 2602.550 ;
        RECT 1715.050 2599.150 1715.490 2599.450 ;
        RECT 1707.815 2593.015 1708.145 2593.345 ;
        RECT 1709.670 2587.905 1709.970 2599.150 ;
        RECT 1715.190 2591.985 1715.490 2599.150 ;
        RECT 1715.175 2591.655 1715.505 2591.985 ;
        RECT 1717.030 2587.905 1717.330 2602.550 ;
        RECT 1720.890 2601.150 1721.190 2604.600 ;
        RECT 1718.870 2600.850 1721.190 2601.150 ;
        RECT 1718.870 2591.985 1719.170 2600.850 ;
        RECT 1720.890 2600.000 1721.190 2600.850 ;
        RECT 1721.510 2601.150 1721.810 2604.600 ;
        RECT 1726.730 2601.150 1727.030 2604.600 ;
        RECT 1721.510 2600.000 1721.930 2601.150 ;
        RECT 1718.855 2591.655 1719.185 2591.985 ;
        RECT 1721.630 2587.905 1721.930 2600.000 ;
        RECT 1725.310 2600.850 1727.030 2601.150 ;
        RECT 1725.310 2592.665 1725.610 2600.850 ;
        RECT 1726.730 2600.000 1727.030 2600.850 ;
        RECT 1727.350 2601.150 1727.650 2604.600 ;
        RECT 1727.350 2600.850 1730.210 2601.150 ;
        RECT 1727.350 2600.000 1727.650 2600.850 ;
        RECT 1725.295 2592.335 1725.625 2592.665 ;
        RECT 1729.910 2587.905 1730.210 2600.850 ;
        RECT 1732.570 2599.450 1732.870 2604.600 ;
        RECT 1733.190 2601.150 1733.490 2604.600 ;
        RECT 1738.410 2601.150 1738.710 2604.600 ;
        RECT 1733.190 2600.850 1736.650 2601.150 ;
        RECT 1733.190 2600.000 1733.490 2600.850 ;
        RECT 1732.570 2599.150 1732.970 2599.450 ;
        RECT 1732.670 2593.345 1732.970 2599.150 ;
        RECT 1732.655 2593.015 1732.985 2593.345 ;
        RECT 1736.350 2587.905 1736.650 2600.850 ;
        RECT 1738.190 2600.000 1738.710 2601.150 ;
        RECT 1739.030 2601.150 1739.330 2604.600 ;
        RECT 1739.030 2600.850 1742.170 2601.150 ;
        RECT 1739.030 2600.000 1739.330 2600.850 ;
        RECT 1738.190 2594.025 1738.490 2600.000 ;
        RECT 1738.175 2593.695 1738.505 2594.025 ;
        RECT 1741.870 2588.585 1742.170 2600.850 ;
        RECT 1744.250 2599.450 1744.550 2604.600 ;
        RECT 1743.710 2599.150 1744.550 2599.450 ;
        RECT 1743.710 2593.345 1744.010 2599.150 ;
        RECT 1744.870 2596.050 1745.170 2604.600 ;
        RECT 2134.010 2601.150 2134.310 2604.600 ;
        RECT 1744.630 2595.750 1745.170 2596.050 ;
        RECT 2132.870 2600.850 2134.310 2601.150 ;
        RECT 1743.695 2593.015 1744.025 2593.345 ;
        RECT 1741.855 2588.255 1742.185 2588.585 ;
        RECT 1744.630 2587.905 1744.930 2595.750 ;
        RECT 2132.870 2590.625 2133.170 2600.850 ;
        RECT 2134.010 2600.000 2134.310 2600.850 ;
        RECT 2139.850 2598.785 2140.150 2604.600 ;
        RECT 2145.690 2601.150 2145.990 2604.600 ;
        RECT 2151.530 2601.150 2151.830 2604.600 ;
        RECT 2157.370 2601.150 2157.670 2604.600 ;
        RECT 2145.690 2600.000 2146.050 2601.150 ;
        RECT 2139.835 2598.455 2140.165 2598.785 ;
        RECT 2145.750 2591.985 2146.050 2600.000 ;
        RECT 2148.510 2600.850 2151.830 2601.150 ;
        RECT 2148.510 2593.345 2148.810 2600.850 ;
        RECT 2151.530 2600.000 2151.830 2600.850 ;
        RECT 2154.030 2600.850 2157.670 2601.150 ;
        RECT 2148.495 2593.015 2148.825 2593.345 ;
        RECT 2154.030 2592.665 2154.330 2600.850 ;
        RECT 2157.370 2600.000 2157.670 2600.850 ;
        RECT 2163.210 2599.450 2163.510 2604.600 ;
        RECT 2163.830 2601.150 2164.130 2604.600 ;
        RECT 2169.050 2601.150 2169.350 2604.600 ;
        RECT 2163.830 2600.850 2165.370 2601.150 ;
        RECT 2163.830 2600.000 2164.130 2600.850 ;
        RECT 2163.210 2599.150 2163.530 2599.450 ;
        RECT 2154.015 2592.335 2154.345 2592.665 ;
        RECT 2145.735 2591.655 2146.065 2591.985 ;
        RECT 2132.855 2590.295 2133.185 2590.625 ;
        RECT 2163.230 2588.585 2163.530 2599.150 ;
        RECT 2165.070 2588.585 2165.370 2600.850 ;
        RECT 2168.750 2600.000 2169.350 2601.150 ;
        RECT 2168.750 2589.265 2169.050 2600.000 ;
        RECT 2168.735 2588.935 2169.065 2589.265 ;
        RECT 2169.670 2588.585 2169.970 2604.600 ;
        RECT 2174.890 2599.450 2175.190 2604.600 ;
        RECT 2175.510 2601.150 2175.810 2604.600 ;
        RECT 2180.730 2601.150 2181.030 2604.600 ;
        RECT 2175.510 2600.850 2179.170 2601.150 ;
        RECT 2175.510 2600.000 2175.810 2600.850 ;
        RECT 2174.890 2599.150 2175.490 2599.450 ;
        RECT 2175.190 2590.625 2175.490 2599.150 ;
        RECT 2175.175 2590.295 2175.505 2590.625 ;
        RECT 2178.870 2588.585 2179.170 2600.850 ;
        RECT 2180.710 2600.000 2181.030 2601.150 ;
        RECT 2181.350 2601.150 2181.650 2604.600 ;
        RECT 2181.350 2600.850 2184.690 2601.150 ;
        RECT 2181.350 2600.000 2181.650 2600.850 ;
        RECT 2180.710 2590.625 2181.010 2600.000 ;
        RECT 2180.695 2590.295 2181.025 2590.625 ;
        RECT 2184.390 2588.585 2184.690 2600.850 ;
        RECT 2186.570 2599.450 2186.870 2604.600 ;
        RECT 2187.190 2601.150 2187.490 2604.600 ;
        RECT 2192.410 2601.150 2192.710 2604.600 ;
        RECT 2187.190 2600.850 2190.210 2601.150 ;
        RECT 2187.190 2600.000 2187.490 2600.850 ;
        RECT 2186.230 2599.150 2186.870 2599.450 ;
        RECT 2186.230 2589.945 2186.530 2599.150 ;
        RECT 2186.215 2589.615 2186.545 2589.945 ;
        RECT 2189.910 2588.585 2190.210 2600.850 ;
        RECT 2191.750 2600.850 2192.710 2601.150 ;
        RECT 2163.215 2588.255 2163.545 2588.585 ;
        RECT 2165.055 2588.255 2165.385 2588.585 ;
        RECT 2169.655 2588.255 2169.985 2588.585 ;
        RECT 2178.855 2588.255 2179.185 2588.585 ;
        RECT 2184.375 2588.255 2184.705 2588.585 ;
        RECT 2189.895 2588.255 2190.225 2588.585 ;
        RECT 2191.750 2587.905 2192.050 2600.850 ;
        RECT 2192.410 2600.000 2192.710 2600.850 ;
        RECT 2193.030 2599.450 2193.330 2604.600 ;
        RECT 2198.250 2601.150 2198.550 2604.600 ;
        RECT 2198.190 2600.000 2198.550 2601.150 ;
        RECT 2198.870 2601.150 2199.170 2604.600 ;
        RECT 2198.870 2600.850 2200.330 2601.150 ;
        RECT 2198.870 2600.000 2199.170 2600.850 ;
        RECT 2193.030 2599.150 2193.890 2599.450 ;
        RECT 2193.590 2587.905 2193.890 2599.150 ;
        RECT 2198.190 2588.585 2198.490 2600.000 ;
        RECT 2198.175 2588.255 2198.505 2588.585 ;
        RECT 2200.030 2587.905 2200.330 2600.850 ;
        RECT 2204.090 2599.450 2204.390 2604.600 ;
        RECT 2204.710 2601.150 2205.010 2604.600 ;
        RECT 2209.930 2601.150 2210.230 2604.600 ;
        RECT 2204.710 2600.850 2207.690 2601.150 ;
        RECT 2204.710 2600.000 2205.010 2600.850 ;
        RECT 2203.710 2599.150 2204.390 2599.450 ;
        RECT 2203.710 2588.585 2204.010 2599.150 ;
        RECT 2203.695 2588.255 2204.025 2588.585 ;
        RECT 2207.390 2587.905 2207.690 2600.850 ;
        RECT 2209.230 2600.850 2210.230 2601.150 ;
        RECT 2209.230 2591.305 2209.530 2600.850 ;
        RECT 2209.930 2600.000 2210.230 2600.850 ;
        RECT 2210.550 2601.150 2210.850 2604.600 ;
        RECT 2215.770 2601.150 2216.070 2604.600 ;
        RECT 2210.550 2600.850 2214.130 2601.150 ;
        RECT 2210.550 2600.000 2210.850 2600.850 ;
        RECT 2209.215 2590.975 2209.545 2591.305 ;
        RECT 2213.830 2587.905 2214.130 2600.850 ;
        RECT 2215.670 2600.000 2216.070 2601.150 ;
        RECT 2216.390 2601.150 2216.690 2604.600 ;
        RECT 2221.610 2601.150 2221.910 2604.600 ;
        RECT 2216.390 2600.850 2219.650 2601.150 ;
        RECT 2216.390 2600.000 2216.690 2600.850 ;
        RECT 2215.670 2594.025 2215.970 2600.000 ;
        RECT 2215.655 2593.695 2215.985 2594.025 ;
        RECT 2219.350 2587.905 2219.650 2600.850 ;
        RECT 2220.270 2600.850 2221.910 2601.150 ;
        RECT 2220.270 2593.345 2220.570 2600.850 ;
        RECT 2221.610 2600.000 2221.910 2600.850 ;
        RECT 2222.230 2601.150 2222.530 2604.600 ;
        RECT 2227.450 2601.150 2227.750 2604.600 ;
        RECT 2222.230 2600.850 2225.170 2601.150 ;
        RECT 2222.230 2600.000 2222.530 2600.850 ;
        RECT 2220.255 2593.015 2220.585 2593.345 ;
        RECT 2224.870 2588.585 2225.170 2600.850 ;
        RECT 2226.710 2600.850 2227.750 2601.150 ;
        RECT 2226.710 2591.305 2227.010 2600.850 ;
        RECT 2227.450 2600.000 2227.750 2600.850 ;
        RECT 2228.070 2599.450 2228.370 2604.600 ;
        RECT 2233.290 2601.150 2233.590 2604.600 ;
        RECT 2227.630 2599.150 2228.370 2599.450 ;
        RECT 2233.150 2600.000 2233.590 2601.150 ;
        RECT 2233.910 2601.150 2234.210 2604.600 ;
        RECT 2233.910 2600.850 2235.290 2601.150 ;
        RECT 2233.910 2600.000 2234.210 2600.850 ;
        RECT 2226.695 2590.975 2227.025 2591.305 ;
        RECT 2224.855 2588.255 2225.185 2588.585 ;
        RECT 2227.630 2587.905 2227.930 2599.150 ;
        RECT 2233.150 2591.985 2233.450 2600.000 ;
        RECT 2233.135 2591.655 2233.465 2591.985 ;
        RECT 2234.990 2587.905 2235.290 2600.850 ;
        RECT 2239.130 2599.450 2239.430 2604.600 ;
        RECT 2239.750 2601.150 2240.050 2604.600 ;
        RECT 2244.970 2601.150 2245.270 2604.600 ;
        RECT 2239.750 2600.850 2241.730 2601.150 ;
        RECT 2239.750 2600.000 2240.050 2600.850 ;
        RECT 2238.670 2599.150 2239.430 2599.450 ;
        RECT 2238.670 2592.665 2238.970 2599.150 ;
        RECT 2238.655 2592.335 2238.985 2592.665 ;
        RECT 2241.430 2587.905 2241.730 2600.850 ;
        RECT 2244.190 2600.850 2245.270 2601.150 ;
        RECT 2244.190 2591.985 2244.490 2600.850 ;
        RECT 2244.970 2600.000 2245.270 2600.850 ;
        RECT 2245.590 2601.150 2245.890 2604.600 ;
        RECT 2250.810 2601.150 2251.110 2604.600 ;
        RECT 2245.590 2600.850 2249.090 2601.150 ;
        RECT 2245.590 2600.000 2245.890 2600.850 ;
        RECT 2244.175 2591.655 2244.505 2591.985 ;
        RECT 2248.790 2587.905 2249.090 2600.850 ;
        RECT 2249.710 2600.850 2251.110 2601.150 ;
        RECT 2249.710 2592.665 2250.010 2600.850 ;
        RECT 2250.810 2600.000 2251.110 2600.850 ;
        RECT 2251.430 2601.150 2251.730 2604.600 ;
        RECT 2251.430 2600.850 2254.610 2601.150 ;
        RECT 2251.430 2600.000 2251.730 2600.850 ;
        RECT 2249.695 2592.335 2250.025 2592.665 ;
        RECT 2254.310 2587.905 2254.610 2600.850 ;
        RECT 2256.650 2599.450 2256.950 2604.600 ;
        RECT 2257.270 2601.150 2257.570 2604.600 ;
        RECT 2257.270 2600.850 2260.130 2601.150 ;
        RECT 2257.270 2600.000 2257.570 2600.850 ;
        RECT 2256.150 2599.150 2256.950 2599.450 ;
        RECT 2256.150 2594.025 2256.450 2599.150 ;
        RECT 2256.135 2593.695 2256.465 2594.025 ;
        RECT 2259.830 2587.905 2260.130 2600.850 ;
        RECT 2262.490 2599.450 2262.790 2604.600 ;
        RECT 2263.110 2601.150 2263.410 2604.600 ;
        RECT 2268.330 2601.150 2268.630 2604.600 ;
        RECT 2263.110 2600.850 2266.570 2601.150 ;
        RECT 2263.110 2600.000 2263.410 2600.850 ;
        RECT 2262.490 2599.150 2262.890 2599.450 ;
        RECT 2262.590 2594.025 2262.890 2599.150 ;
        RECT 2262.575 2593.695 2262.905 2594.025 ;
        RECT 2266.270 2588.585 2266.570 2600.850 ;
        RECT 2268.110 2600.000 2268.630 2601.150 ;
        RECT 2268.950 2601.150 2269.250 2604.600 ;
        RECT 2268.950 2600.000 2269.330 2601.150 ;
        RECT 2268.110 2594.025 2268.410 2600.000 ;
        RECT 2268.095 2593.695 2268.425 2594.025 ;
        RECT 2266.255 2588.255 2266.585 2588.585 ;
        RECT 2269.030 2587.905 2269.330 2600.000 ;
        RECT 2274.170 2599.450 2274.470 2604.600 ;
        RECT 2274.790 2601.150 2275.090 2604.600 ;
        RECT 2274.790 2600.850 2276.690 2601.150 ;
        RECT 2274.790 2600.000 2275.090 2600.850 ;
        RECT 2273.630 2599.150 2274.470 2599.450 ;
        RECT 2273.630 2591.985 2273.930 2599.150 ;
        RECT 2273.615 2591.655 2273.945 2591.985 ;
        RECT 2276.390 2587.905 2276.690 2600.850 ;
        RECT 2280.010 2599.450 2280.310 2604.600 ;
        RECT 2280.630 2601.150 2280.930 2604.600 ;
        RECT 2285.850 2601.150 2286.150 2604.600 ;
        RECT 2280.630 2600.850 2282.210 2601.150 ;
        RECT 2280.630 2600.000 2280.930 2600.850 ;
        RECT 2280.010 2599.150 2280.370 2599.450 ;
        RECT 2280.070 2592.665 2280.370 2599.150 ;
        RECT 2280.055 2592.335 2280.385 2592.665 ;
        RECT 2281.910 2587.905 2282.210 2600.850 ;
        RECT 2285.590 2600.000 2286.150 2601.150 ;
        RECT 2286.470 2601.150 2286.770 2604.600 ;
        RECT 2286.470 2600.850 2289.570 2601.150 ;
        RECT 2286.470 2600.000 2286.770 2600.850 ;
        RECT 2285.590 2592.665 2285.890 2600.000 ;
        RECT 2285.575 2592.335 2285.905 2592.665 ;
        RECT 2289.270 2587.905 2289.570 2600.850 ;
        RECT 2291.690 2599.450 2291.990 2604.600 ;
        RECT 2292.310 2601.150 2292.610 2604.600 ;
        RECT 2292.310 2600.850 2296.010 2601.150 ;
        RECT 2292.310 2600.000 2292.610 2600.850 ;
        RECT 2291.690 2599.150 2292.330 2599.450 ;
        RECT 2292.030 2593.345 2292.330 2599.150 ;
        RECT 2292.015 2593.015 2292.345 2593.345 ;
        RECT 2295.710 2587.905 2296.010 2600.850 ;
        RECT 2297.530 2599.450 2297.830 2604.600 ;
        RECT 2298.150 2601.150 2298.450 2604.600 ;
        RECT 2303.370 2601.150 2303.670 2604.600 ;
        RECT 2298.150 2600.850 2301.530 2601.150 ;
        RECT 2298.150 2600.000 2298.450 2600.850 ;
        RECT 2297.530 2599.150 2297.850 2599.450 ;
        RECT 2297.550 2593.345 2297.850 2599.150 ;
        RECT 2297.535 2593.015 2297.865 2593.345 ;
        RECT 2301.230 2588.585 2301.530 2600.850 ;
        RECT 2302.150 2600.850 2303.670 2601.150 ;
        RECT 2302.150 2594.025 2302.450 2600.850 ;
        RECT 2303.370 2600.000 2303.670 2600.850 ;
        RECT 2302.135 2593.695 2302.465 2594.025 ;
        RECT 2301.215 2588.255 2301.545 2588.585 ;
        RECT 2303.990 2587.905 2304.290 2604.600 ;
        RECT 2309.210 2601.150 2309.510 2604.600 ;
        RECT 2305.830 2600.850 2309.510 2601.150 ;
        RECT 2305.830 2594.025 2306.130 2600.850 ;
        RECT 2309.210 2600.000 2309.510 2600.850 ;
        RECT 2309.830 2601.150 2310.130 2604.600 ;
        RECT 2315.050 2601.150 2315.350 2604.600 ;
        RECT 2309.830 2600.850 2310.730 2601.150 ;
        RECT 2309.830 2600.000 2310.130 2600.850 ;
        RECT 2305.815 2593.695 2306.145 2594.025 ;
        RECT 2310.430 2587.905 2310.730 2600.850 ;
        RECT 2312.270 2600.850 2315.350 2601.150 ;
        RECT 2312.270 2593.345 2312.570 2600.850 ;
        RECT 2315.050 2600.000 2315.350 2600.850 ;
        RECT 2315.670 2601.150 2315.970 2604.600 ;
        RECT 2320.890 2601.150 2321.190 2604.600 ;
        RECT 2315.670 2600.850 2318.090 2601.150 ;
        RECT 2315.670 2600.000 2315.970 2600.850 ;
        RECT 2312.255 2593.015 2312.585 2593.345 ;
        RECT 2317.790 2587.905 2318.090 2600.850 ;
        RECT 2319.630 2600.850 2321.190 2601.150 ;
        RECT 2319.630 2591.985 2319.930 2600.850 ;
        RECT 2320.890 2600.000 2321.190 2600.850 ;
        RECT 2321.510 2601.150 2321.810 2604.600 ;
        RECT 2326.730 2601.150 2327.030 2604.600 ;
        RECT 2321.510 2600.850 2324.530 2601.150 ;
        RECT 2321.510 2600.000 2321.810 2600.850 ;
        RECT 2319.615 2591.655 2319.945 2591.985 ;
        RECT 2324.230 2587.905 2324.530 2600.850 ;
        RECT 2326.070 2600.850 2327.030 2601.150 ;
        RECT 2326.070 2591.305 2326.370 2600.850 ;
        RECT 2326.730 2600.000 2327.030 2600.850 ;
        RECT 2327.350 2601.150 2327.650 2604.600 ;
        RECT 2332.570 2601.150 2332.870 2604.600 ;
        RECT 2327.350 2600.850 2330.970 2601.150 ;
        RECT 2327.350 2600.000 2327.650 2600.850 ;
        RECT 2326.055 2590.975 2326.385 2591.305 ;
        RECT 2330.670 2587.905 2330.970 2600.850 ;
        RECT 2332.510 2600.000 2332.870 2601.150 ;
        RECT 2333.190 2601.150 2333.490 2604.600 ;
        RECT 2338.410 2601.150 2338.710 2604.600 ;
        RECT 2333.190 2600.850 2336.490 2601.150 ;
        RECT 2333.190 2600.000 2333.490 2600.850 ;
        RECT 2332.510 2591.985 2332.810 2600.000 ;
        RECT 2332.495 2591.655 2332.825 2591.985 ;
        RECT 2336.190 2587.905 2336.490 2600.850 ;
        RECT 2337.110 2600.850 2338.710 2601.150 ;
        RECT 2337.110 2593.345 2337.410 2600.850 ;
        RECT 2338.410 2600.000 2338.710 2600.850 ;
        RECT 2339.030 2601.150 2339.330 2604.600 ;
        RECT 2344.250 2601.150 2344.550 2604.600 ;
        RECT 2339.030 2600.850 2342.010 2601.150 ;
        RECT 2339.030 2600.000 2339.330 2600.850 ;
        RECT 2337.095 2593.015 2337.425 2593.345 ;
        RECT 2341.710 2588.585 2342.010 2600.850 ;
        RECT 2342.630 2600.850 2344.550 2601.150 ;
        RECT 2342.630 2592.665 2342.930 2600.850 ;
        RECT 2344.250 2600.000 2344.550 2600.850 ;
        RECT 2344.870 2599.450 2345.170 2604.600 ;
        RECT 2344.870 2599.150 2345.690 2599.450 ;
        RECT 2342.615 2592.335 2342.945 2592.665 ;
        RECT 2341.695 2588.255 2342.025 2588.585 ;
        RECT 2345.390 2587.905 2345.690 2599.150 ;
        RECT 1536.695 2587.575 1537.025 2587.905 ;
        RECT 1543.135 2587.575 1543.465 2587.905 ;
        RECT 1548.655 2587.575 1548.985 2587.905 ;
        RECT 1558.775 2587.575 1559.105 2587.905 ;
        RECT 1651.695 2587.575 1652.025 2587.905 ;
        RECT 1703.215 2587.575 1703.545 2587.905 ;
        RECT 1709.655 2587.575 1709.985 2587.905 ;
        RECT 1717.015 2587.575 1717.345 2587.905 ;
        RECT 1721.615 2587.575 1721.945 2587.905 ;
        RECT 1729.895 2587.575 1730.225 2587.905 ;
        RECT 1736.335 2587.575 1736.665 2587.905 ;
        RECT 1744.615 2587.575 1744.945 2587.905 ;
        RECT 2191.735 2587.575 2192.065 2587.905 ;
        RECT 2193.575 2587.575 2193.905 2587.905 ;
        RECT 2200.015 2587.575 2200.345 2587.905 ;
        RECT 2207.375 2587.575 2207.705 2587.905 ;
        RECT 2213.815 2587.575 2214.145 2587.905 ;
        RECT 2219.335 2587.575 2219.665 2587.905 ;
        RECT 2227.615 2587.575 2227.945 2587.905 ;
        RECT 2234.975 2587.575 2235.305 2587.905 ;
        RECT 2241.415 2587.575 2241.745 2587.905 ;
        RECT 2248.775 2587.575 2249.105 2587.905 ;
        RECT 2254.295 2587.575 2254.625 2587.905 ;
        RECT 2259.815 2587.575 2260.145 2587.905 ;
        RECT 2269.015 2587.575 2269.345 2587.905 ;
        RECT 2276.375 2587.575 2276.705 2587.905 ;
        RECT 2281.895 2587.575 2282.225 2587.905 ;
        RECT 2289.255 2587.575 2289.585 2587.905 ;
        RECT 2295.695 2587.575 2296.025 2587.905 ;
        RECT 2303.975 2587.575 2304.305 2587.905 ;
        RECT 2310.415 2587.575 2310.745 2587.905 ;
        RECT 2317.775 2587.575 2318.105 2587.905 ;
        RECT 2324.215 2587.575 2324.545 2587.905 ;
        RECT 2330.655 2587.575 2330.985 2587.905 ;
        RECT 2336.175 2587.575 2336.505 2587.905 ;
        RECT 2345.375 2587.575 2345.705 2587.905 ;
        RECT 1498.020 2415.000 1501.020 2585.000 ;
        RECT 1678.020 2415.000 1681.020 2585.000 ;
        RECT 1858.020 2415.000 1861.020 2585.000 ;
        RECT 2218.020 2415.000 2221.020 2585.000 ;
        RECT 2398.020 2415.000 2401.020 2585.000 ;
      LAYER met4 ;
        RECT 1415.935 2389.280 2588.345 2395.945 ;
        RECT 1415.935 1210.640 1420.640 2389.280 ;
        RECT 1423.040 1210.640 1497.440 2389.280 ;
        RECT 1499.840 1210.640 2588.345 2389.280 ;
      LAYER met4 ;
        RECT 1552.020 1021.235 1555.020 1185.000 ;
        RECT 1647.095 1062.335 1647.425 1062.665 ;
        RECT 1641.575 1016.775 1641.905 1017.105 ;
        RECT 1640.655 1016.095 1640.985 1016.425 ;
        RECT 1640.670 1004.850 1640.970 1016.095 ;
        RECT 1641.590 1008.250 1641.890 1016.775 ;
        RECT 1641.590 1007.950 1642.230 1008.250 ;
        RECT 1641.310 1004.850 1641.610 1006.235 ;
        RECT 1640.670 1004.550 1641.610 1004.850 ;
        RECT 1641.310 1001.635 1641.610 1004.550 ;
        RECT 1641.930 1001.635 1642.230 1007.950 ;
        RECT 1647.110 1006.235 1647.410 1062.335 ;
        RECT 1682.055 1038.535 1682.385 1038.865 ;
        RECT 1654.455 1016.775 1654.785 1017.105 ;
        RECT 1671.015 1016.775 1671.345 1017.105 ;
        RECT 1653.535 1016.095 1653.865 1016.425 ;
        RECT 1648.015 1014.735 1648.345 1015.065 ;
        RECT 1648.030 1006.235 1648.330 1014.735 ;
        RECT 1653.550 1008.250 1653.850 1016.095 ;
        RECT 1647.110 1004.550 1647.450 1006.235 ;
        RECT 1647.150 1001.635 1647.450 1004.550 ;
        RECT 1647.770 1004.550 1648.330 1006.235 ;
        RECT 1652.990 1007.950 1653.850 1008.250 ;
        RECT 1647.770 1001.635 1648.070 1004.550 ;
        RECT 1652.990 1001.635 1653.290 1007.950 ;
        RECT 1653.610 1004.850 1653.910 1006.235 ;
        RECT 1654.470 1004.850 1654.770 1016.775 ;
        RECT 1658.135 1016.095 1658.465 1016.425 ;
        RECT 1664.575 1016.095 1664.905 1016.425 ;
        RECT 1653.610 1004.550 1654.770 1004.850 ;
        RECT 1658.150 1004.850 1658.450 1016.095 ;
        RECT 1661.815 1015.415 1662.145 1015.745 ;
        RECT 1658.830 1004.850 1659.130 1006.235 ;
        RECT 1658.150 1004.550 1659.130 1004.850 ;
        RECT 1653.610 1001.635 1653.910 1004.550 ;
        RECT 1658.830 1001.635 1659.130 1004.550 ;
        RECT 1659.450 1004.850 1659.750 1006.235 ;
        RECT 1661.830 1004.850 1662.130 1015.415 ;
        RECT 1659.450 1004.550 1662.130 1004.850 ;
        RECT 1664.590 1006.235 1664.890 1016.095 ;
        RECT 1668.255 1015.415 1668.585 1015.745 ;
        RECT 1664.590 1004.550 1664.970 1006.235 ;
        RECT 1659.450 1001.635 1659.750 1004.550 ;
        RECT 1664.670 1001.635 1664.970 1004.550 ;
        RECT 1665.290 1004.850 1665.590 1006.235 ;
        RECT 1668.270 1004.850 1668.570 1015.415 ;
        RECT 1671.030 1008.250 1671.330 1016.775 ;
        RECT 1675.615 1016.095 1675.945 1016.425 ;
        RECT 1673.775 1015.415 1674.105 1015.745 ;
        RECT 1665.290 1004.550 1668.570 1004.850 ;
        RECT 1670.510 1007.950 1671.330 1008.250 ;
        RECT 1665.290 1001.635 1665.590 1004.550 ;
        RECT 1670.510 1001.635 1670.810 1007.950 ;
        RECT 1671.130 1004.850 1671.430 1006.235 ;
        RECT 1673.790 1004.850 1674.090 1015.415 ;
        RECT 1671.130 1004.550 1674.090 1004.850 ;
        RECT 1675.630 1004.850 1675.930 1016.095 ;
        RECT 1680.215 1014.735 1680.545 1015.065 ;
        RECT 1676.350 1004.850 1676.650 1006.235 ;
        RECT 1675.630 1004.550 1676.650 1004.850 ;
        RECT 1671.130 1001.635 1671.430 1004.550 ;
        RECT 1676.350 1001.635 1676.650 1004.550 ;
        RECT 1676.970 1004.850 1677.270 1006.235 ;
        RECT 1680.230 1004.850 1680.530 1014.735 ;
        RECT 1676.970 1004.550 1680.530 1004.850 ;
        RECT 1682.070 1006.235 1682.370 1038.535 ;
        RECT 1732.020 1021.235 1735.020 1185.000 ;
        RECT 2092.020 1021.235 2095.020 1185.000 ;
        RECT 2272.020 1021.235 2275.020 1185.000 ;
        RECT 2452.020 1021.235 2455.020 1185.000 ;
        RECT 1704.135 1020.855 1704.465 1021.185 ;
        RECT 1834.775 1020.855 1835.105 1021.185 ;
        RECT 1843.975 1020.855 1844.305 1021.185 ;
        RECT 1855.015 1020.855 1855.345 1021.185 ;
        RECT 2241.415 1020.855 2241.745 1021.185 ;
        RECT 2260.735 1020.855 2261.065 1021.185 ;
        RECT 2266.255 1020.855 2266.585 1021.185 ;
        RECT 2270.855 1020.855 2271.185 1021.185 ;
        RECT 2281.895 1020.855 2282.225 1021.185 ;
        RECT 2328.815 1020.855 2329.145 1021.185 ;
        RECT 2333.415 1020.855 2333.745 1021.185 ;
        RECT 2340.775 1020.855 2341.105 1021.185 ;
        RECT 2351.815 1020.855 2352.145 1021.185 ;
        RECT 2358.255 1020.855 2358.585 1021.185 ;
        RECT 2373.895 1020.855 2374.225 1021.185 ;
        RECT 2403.335 1020.855 2403.665 1021.185 ;
        RECT 2421.735 1020.855 2422.065 1021.185 ;
        RECT 1684.815 1016.775 1685.145 1017.105 ;
        RECT 1682.975 1015.415 1683.305 1015.745 ;
        RECT 1682.990 1006.235 1683.290 1015.415 ;
        RECT 1682.070 1004.550 1682.490 1006.235 ;
        RECT 1676.970 1001.635 1677.270 1004.550 ;
        RECT 1682.190 1001.635 1682.490 1004.550 ;
        RECT 1682.810 1004.550 1683.290 1006.235 ;
        RECT 1684.830 1004.850 1685.130 1016.775 ;
        RECT 1692.175 1016.095 1692.505 1016.425 ;
        RECT 1698.615 1016.095 1698.945 1016.425 ;
        RECT 1689.415 1014.735 1689.745 1015.065 ;
        RECT 1688.030 1004.850 1688.330 1006.235 ;
        RECT 1684.830 1004.550 1688.330 1004.850 ;
        RECT 1682.810 1001.635 1683.110 1004.550 ;
        RECT 1688.030 1001.635 1688.330 1004.550 ;
        RECT 1688.650 1004.850 1688.950 1006.235 ;
        RECT 1689.430 1004.850 1689.730 1014.735 ;
        RECT 1688.650 1004.550 1689.730 1004.850 ;
        RECT 1692.190 1004.850 1692.490 1016.095 ;
        RECT 1695.855 1014.735 1696.185 1015.065 ;
        RECT 1693.870 1004.850 1694.170 1006.235 ;
        RECT 1692.190 1004.550 1694.170 1004.850 ;
        RECT 1688.650 1001.635 1688.950 1004.550 ;
        RECT 1693.870 1001.635 1694.170 1004.550 ;
        RECT 1694.490 1004.085 1694.790 1006.235 ;
        RECT 1695.870 1004.085 1696.170 1014.735 ;
        RECT 1698.630 1004.850 1698.930 1016.095 ;
        RECT 1700.455 1014.735 1700.785 1015.065 ;
        RECT 1700.470 1006.235 1700.770 1014.735 ;
        RECT 1699.710 1004.850 1700.010 1006.235 ;
        RECT 1698.630 1004.550 1700.010 1004.850 ;
        RECT 1694.490 1003.785 1696.170 1004.085 ;
        RECT 1694.490 1001.635 1694.790 1003.785 ;
        RECT 1699.710 1001.635 1700.010 1004.550 ;
        RECT 1700.330 1004.550 1700.770 1006.235 ;
        RECT 1700.330 1001.635 1700.630 1004.550 ;
        RECT 1704.150 1004.085 1704.450 1020.855 ;
        RECT 1786.935 1019.495 1787.265 1019.825 ;
        RECT 1801.655 1019.495 1801.985 1019.825 ;
        RECT 1832.015 1019.495 1832.345 1019.825 ;
        RECT 1711.495 1018.135 1711.825 1018.465 ;
        RECT 1719.775 1018.135 1720.105 1018.465 ;
        RECT 1745.535 1018.135 1745.865 1018.465 ;
        RECT 1763.935 1018.135 1764.265 1018.465 ;
        RECT 1774.055 1018.135 1774.385 1018.465 ;
        RECT 1706.895 1014.735 1707.225 1015.065 ;
        RECT 1705.550 1004.085 1705.850 1006.235 ;
        RECT 1704.150 1003.785 1705.850 1004.085 ;
        RECT 1705.550 1001.635 1705.850 1003.785 ;
        RECT 1706.170 1004.850 1706.470 1006.235 ;
        RECT 1706.910 1004.850 1707.210 1014.735 ;
        RECT 1711.510 1008.250 1711.810 1018.135 ;
        RECT 1714.255 1017.455 1714.585 1017.785 ;
        RECT 1713.335 1014.735 1713.665 1015.065 ;
        RECT 1706.170 1004.550 1707.210 1004.850 ;
        RECT 1711.390 1007.950 1711.810 1008.250 ;
        RECT 1706.170 1001.635 1706.470 1004.550 ;
        RECT 1711.390 1001.635 1711.690 1007.950 ;
        RECT 1712.010 1004.085 1712.310 1006.235 ;
        RECT 1713.350 1004.085 1713.650 1014.735 ;
        RECT 1714.270 1004.850 1714.570 1017.455 ;
        RECT 1717.935 1014.735 1718.265 1015.065 ;
        RECT 1717.950 1006.235 1718.250 1014.735 ;
        RECT 1717.230 1004.850 1717.530 1006.235 ;
        RECT 1714.270 1004.550 1717.530 1004.850 ;
        RECT 1712.010 1003.785 1713.650 1004.085 ;
        RECT 1712.010 1001.635 1712.310 1003.785 ;
        RECT 1717.230 1001.635 1717.530 1004.550 ;
        RECT 1717.850 1004.550 1718.250 1006.235 ;
        RECT 1719.790 1004.850 1720.090 1018.135 ;
        RECT 1726.215 1016.095 1726.545 1016.425 ;
        RECT 1732.655 1016.095 1732.985 1016.425 ;
        RECT 1724.375 1014.735 1724.705 1015.065 ;
        RECT 1723.070 1004.850 1723.370 1006.235 ;
        RECT 1719.790 1004.550 1723.370 1004.850 ;
        RECT 1717.850 1001.635 1718.150 1004.550 ;
        RECT 1723.070 1001.635 1723.370 1004.550 ;
        RECT 1723.690 1004.850 1723.990 1006.235 ;
        RECT 1724.390 1004.850 1724.690 1014.735 ;
        RECT 1723.690 1004.550 1724.690 1004.850 ;
        RECT 1726.230 1004.850 1726.530 1016.095 ;
        RECT 1730.815 1014.735 1731.145 1015.065 ;
        RECT 1728.910 1004.850 1729.210 1006.235 ;
        RECT 1726.230 1004.550 1729.210 1004.850 ;
        RECT 1723.690 1001.635 1723.990 1004.550 ;
        RECT 1728.910 1001.635 1729.210 1004.550 ;
        RECT 1729.530 1004.085 1729.830 1006.235 ;
        RECT 1730.830 1004.085 1731.130 1014.735 ;
        RECT 1732.670 1004.850 1732.970 1016.095 ;
        RECT 1739.095 1015.415 1739.425 1015.745 ;
        RECT 1735.415 1014.735 1735.745 1015.065 ;
        RECT 1735.430 1006.235 1735.730 1014.735 ;
        RECT 1734.750 1004.850 1735.050 1006.235 ;
        RECT 1732.670 1004.550 1735.050 1004.850 ;
        RECT 1729.530 1003.785 1731.130 1004.085 ;
        RECT 1729.530 1001.635 1729.830 1003.785 ;
        RECT 1734.750 1001.635 1735.050 1004.550 ;
        RECT 1735.370 1004.550 1735.730 1006.235 ;
        RECT 1739.110 1004.850 1739.410 1015.415 ;
        RECT 1741.855 1014.735 1742.185 1015.065 ;
        RECT 1740.590 1004.850 1740.890 1006.235 ;
        RECT 1739.110 1004.550 1740.890 1004.850 ;
        RECT 1735.370 1001.635 1735.670 1004.550 ;
        RECT 1740.590 1001.635 1740.890 1004.550 ;
        RECT 1741.210 1004.850 1741.510 1006.235 ;
        RECT 1741.870 1004.850 1742.170 1014.735 ;
        RECT 1741.210 1004.550 1742.170 1004.850 ;
        RECT 1745.550 1004.850 1745.850 1018.135 ;
        RECT 1749.215 1016.095 1749.545 1016.425 ;
        RECT 1748.295 1014.735 1748.625 1015.065 ;
        RECT 1746.430 1004.850 1746.730 1006.235 ;
        RECT 1745.550 1004.550 1746.730 1004.850 ;
        RECT 1741.210 1001.635 1741.510 1004.550 ;
        RECT 1746.430 1001.635 1746.730 1004.550 ;
        RECT 1747.050 1004.085 1747.350 1006.235 ;
        RECT 1748.310 1004.085 1748.610 1014.735 ;
        RECT 1749.230 1004.850 1749.530 1016.095 ;
        RECT 1755.655 1015.415 1755.985 1015.745 ;
        RECT 1754.735 1014.735 1755.065 1015.065 ;
        RECT 1752.270 1004.850 1752.570 1006.235 ;
        RECT 1749.230 1004.550 1752.570 1004.850 ;
        RECT 1747.050 1003.785 1748.610 1004.085 ;
        RECT 1747.050 1001.635 1747.350 1003.785 ;
        RECT 1752.270 1001.635 1752.570 1004.550 ;
        RECT 1752.890 1004.850 1753.190 1006.235 ;
        RECT 1754.750 1004.850 1755.050 1014.735 ;
        RECT 1752.890 1004.550 1755.050 1004.850 ;
        RECT 1755.670 1004.850 1755.970 1015.415 ;
        RECT 1758.415 1014.735 1758.745 1015.065 ;
        RECT 1758.430 1008.250 1758.730 1014.735 ;
        RECT 1758.430 1007.950 1759.030 1008.250 ;
        RECT 1758.110 1004.850 1758.410 1006.235 ;
        RECT 1755.670 1004.550 1758.410 1004.850 ;
        RECT 1752.890 1001.635 1753.190 1004.550 ;
        RECT 1758.110 1001.635 1758.410 1004.550 ;
        RECT 1758.730 1001.635 1759.030 1007.950 ;
        RECT 1763.950 1001.635 1764.250 1018.135 ;
        RECT 1766.695 1015.415 1767.025 1015.745 ;
        RECT 1765.775 1014.735 1766.105 1015.065 ;
        RECT 1764.570 1004.850 1764.870 1006.235 ;
        RECT 1765.790 1004.850 1766.090 1014.735 ;
        RECT 1764.570 1004.550 1766.090 1004.850 ;
        RECT 1766.710 1004.850 1767.010 1015.415 ;
        RECT 1772.215 1014.735 1772.545 1015.065 ;
        RECT 1769.790 1004.850 1770.090 1006.235 ;
        RECT 1766.710 1004.550 1770.090 1004.850 ;
        RECT 1764.570 1001.635 1764.870 1004.550 ;
        RECT 1769.790 1001.635 1770.090 1004.550 ;
        RECT 1770.410 1004.850 1770.710 1006.235 ;
        RECT 1772.230 1004.850 1772.530 1014.735 ;
        RECT 1770.410 1004.550 1772.530 1004.850 ;
        RECT 1774.070 1004.850 1774.370 1018.135 ;
        RECT 1780.495 1016.095 1780.825 1016.425 ;
        RECT 1777.735 1014.735 1778.065 1015.065 ;
        RECT 1775.630 1004.850 1775.930 1006.235 ;
        RECT 1774.070 1004.550 1775.930 1004.850 ;
        RECT 1770.410 1001.635 1770.710 1004.550 ;
        RECT 1775.630 1001.635 1775.930 1004.550 ;
        RECT 1776.250 1004.085 1776.550 1006.235 ;
        RECT 1777.750 1004.085 1778.050 1014.735 ;
        RECT 1780.510 1004.850 1780.810 1016.095 ;
        RECT 1782.335 1014.735 1782.665 1015.065 ;
        RECT 1782.350 1006.235 1782.650 1014.735 ;
        RECT 1786.950 1008.250 1787.250 1019.495 ;
        RECT 1788.775 1015.415 1789.105 1015.745 ;
        RECT 1786.950 1007.950 1787.610 1008.250 ;
        RECT 1781.470 1004.850 1781.770 1006.235 ;
        RECT 1780.510 1004.550 1781.770 1004.850 ;
        RECT 1776.250 1003.785 1778.050 1004.085 ;
        RECT 1776.250 1001.635 1776.550 1003.785 ;
        RECT 1781.470 1001.635 1781.770 1004.550 ;
        RECT 1782.090 1004.550 1782.650 1006.235 ;
        RECT 1782.090 1001.635 1782.390 1004.550 ;
        RECT 1787.310 1001.635 1787.610 1007.950 ;
        RECT 1787.930 1004.850 1788.230 1006.235 ;
        RECT 1788.790 1004.850 1789.090 1015.415 ;
        RECT 1789.695 1014.735 1790.025 1015.065 ;
        RECT 1793.375 1014.735 1793.705 1015.065 ;
        RECT 1796.135 1014.735 1796.465 1015.065 ;
        RECT 1799.815 1014.735 1800.145 1015.065 ;
        RECT 1787.930 1004.550 1789.090 1004.850 ;
        RECT 1789.710 1004.850 1790.010 1014.735 ;
        RECT 1793.390 1008.250 1793.690 1014.735 ;
        RECT 1793.390 1007.950 1794.070 1008.250 ;
        RECT 1793.150 1004.850 1793.450 1006.235 ;
        RECT 1789.710 1004.550 1793.450 1004.850 ;
        RECT 1787.930 1001.635 1788.230 1004.550 ;
        RECT 1793.150 1001.635 1793.450 1004.550 ;
        RECT 1793.770 1001.635 1794.070 1007.950 ;
        RECT 1796.150 1004.850 1796.450 1014.735 ;
        RECT 1799.830 1006.235 1800.130 1014.735 ;
        RECT 1798.990 1004.850 1799.290 1006.235 ;
        RECT 1796.150 1004.550 1799.290 1004.850 ;
        RECT 1798.990 1001.635 1799.290 1004.550 ;
        RECT 1799.610 1004.550 1800.130 1006.235 ;
        RECT 1801.670 1004.850 1801.970 1019.495 ;
        RECT 1808.095 1018.815 1808.425 1019.145 ;
        RECT 1806.255 1014.735 1806.585 1015.065 ;
        RECT 1804.830 1004.850 1805.130 1006.235 ;
        RECT 1801.670 1004.550 1805.130 1004.850 ;
        RECT 1799.610 1001.635 1799.910 1004.550 ;
        RECT 1804.830 1001.635 1805.130 1004.550 ;
        RECT 1805.450 1004.850 1805.750 1006.235 ;
        RECT 1806.270 1004.850 1806.570 1014.735 ;
        RECT 1805.450 1004.550 1806.570 1004.850 ;
        RECT 1808.110 1004.850 1808.410 1018.815 ;
        RECT 1814.535 1016.775 1814.865 1017.105 ;
        RECT 1821.895 1016.775 1822.225 1017.105 ;
        RECT 1812.695 1014.735 1813.025 1015.065 ;
        RECT 1810.670 1004.850 1810.970 1006.235 ;
        RECT 1808.110 1004.550 1810.970 1004.850 ;
        RECT 1805.450 1001.635 1805.750 1004.550 ;
        RECT 1810.670 1001.635 1810.970 1004.550 ;
        RECT 1811.290 1004.085 1811.590 1006.235 ;
        RECT 1812.710 1004.085 1813.010 1014.735 ;
        RECT 1814.550 1004.850 1814.850 1016.775 ;
        RECT 1817.295 1014.735 1817.625 1015.065 ;
        RECT 1817.310 1006.235 1817.610 1014.735 ;
        RECT 1821.910 1008.250 1822.210 1016.775 ;
        RECT 1823.735 1014.735 1824.065 1015.065 ;
        RECT 1821.910 1007.950 1822.650 1008.250 ;
        RECT 1816.510 1004.850 1816.810 1006.235 ;
        RECT 1814.550 1004.550 1816.810 1004.850 ;
        RECT 1811.290 1003.785 1813.010 1004.085 ;
        RECT 1811.290 1001.635 1811.590 1003.785 ;
        RECT 1816.510 1001.635 1816.810 1004.550 ;
        RECT 1817.130 1004.550 1817.610 1006.235 ;
        RECT 1817.130 1001.635 1817.430 1004.550 ;
        RECT 1822.350 1001.635 1822.650 1007.950 ;
        RECT 1822.970 1004.850 1823.270 1006.235 ;
        RECT 1823.750 1004.850 1824.050 1014.735 ;
        RECT 1822.970 1004.550 1824.050 1004.850 ;
        RECT 1828.810 1004.850 1829.110 1006.235 ;
        RECT 1832.030 1004.850 1832.330 1019.495 ;
        RECT 1834.790 1006.235 1835.090 1020.855 ;
        RECT 1837.535 1020.175 1837.865 1020.505 ;
        RECT 1828.810 1004.550 1832.330 1004.850 ;
        RECT 1834.650 1004.550 1835.090 1006.235 ;
        RECT 1837.550 1004.850 1837.850 1020.175 ;
        RECT 1840.490 1004.850 1840.790 1006.235 ;
        RECT 1837.550 1004.550 1840.790 1004.850 ;
        RECT 1843.990 1004.850 1844.290 1020.855 ;
        RECT 1846.330 1004.850 1846.630 1006.235 ;
        RECT 1843.990 1004.550 1846.630 1004.850 ;
        RECT 1822.970 1001.635 1823.270 1004.550 ;
        RECT 1828.810 1001.635 1829.110 1004.550 ;
        RECT 1834.650 1001.635 1834.950 1004.550 ;
        RECT 1840.490 1001.635 1840.790 1004.550 ;
        RECT 1846.330 1001.635 1846.630 1004.550 ;
        RECT 1852.170 1004.850 1852.470 1006.235 ;
        RECT 1855.030 1004.850 1855.330 1020.855 ;
        RECT 2241.430 1007.570 2241.730 1020.855 ;
        RECT 2247.855 1020.175 2248.185 1020.505 ;
        RECT 2254.295 1020.175 2254.625 1020.505 ;
        RECT 2246.935 1014.735 2247.265 1015.065 ;
        RECT 1852.170 1004.550 1855.330 1004.850 ;
        RECT 2241.310 1007.270 2241.730 1007.570 ;
        RECT 1852.170 1001.635 1852.470 1004.550 ;
        RECT 2241.310 1001.635 2241.610 1007.270 ;
        RECT 2241.915 1006.575 2242.245 1006.905 ;
        RECT 2241.930 1001.635 2242.230 1006.575 ;
        RECT 2246.950 1006.235 2247.250 1014.735 ;
        RECT 2247.870 1006.235 2248.170 1020.175 ;
        RECT 2253.375 1014.735 2253.705 1015.065 ;
        RECT 2253.390 1007.570 2253.690 1014.735 ;
        RECT 2246.950 1004.550 2247.450 1006.235 ;
        RECT 2247.150 1001.635 2247.450 1004.550 ;
        RECT 2247.770 1004.550 2248.170 1006.235 ;
        RECT 2252.990 1007.270 2253.690 1007.570 ;
        RECT 2247.770 1001.635 2248.070 1004.550 ;
        RECT 2252.990 1001.635 2253.290 1007.270 ;
        RECT 2253.610 1004.850 2253.910 1006.235 ;
        RECT 2254.310 1004.850 2254.610 1020.175 ;
        RECT 2258.895 1014.735 2259.225 1015.065 ;
        RECT 2258.910 1007.570 2259.210 1014.735 ;
        RECT 2253.610 1004.550 2254.610 1004.850 ;
        RECT 2258.830 1007.270 2259.210 1007.570 ;
        RECT 2253.610 1001.635 2253.910 1004.550 ;
        RECT 2258.830 1001.635 2259.130 1007.270 ;
        RECT 2259.450 1004.085 2259.750 1006.235 ;
        RECT 2260.750 1004.085 2261.050 1020.855 ;
        RECT 2264.415 1016.775 2264.745 1017.105 ;
        RECT 2264.430 1006.235 2264.730 1016.775 ;
        RECT 2264.430 1004.550 2264.970 1006.235 ;
        RECT 2259.450 1003.785 2261.050 1004.085 ;
        RECT 2259.450 1001.635 2259.750 1003.785 ;
        RECT 2264.670 1001.635 2264.970 1004.550 ;
        RECT 2265.290 1004.850 2265.590 1006.235 ;
        RECT 2266.270 1004.850 2266.570 1020.855 ;
        RECT 2270.870 1007.570 2271.170 1020.855 ;
        RECT 2272.695 1019.495 2273.025 1019.825 ;
        RECT 2276.375 1019.495 2276.705 1019.825 ;
        RECT 2265.290 1004.550 2266.570 1004.850 ;
        RECT 2270.510 1007.270 2271.170 1007.570 ;
        RECT 2265.290 1001.635 2265.590 1004.550 ;
        RECT 2270.510 1001.635 2270.810 1007.270 ;
        RECT 2271.130 1004.850 2271.430 1006.235 ;
        RECT 2272.710 1004.850 2273.010 1019.495 ;
        RECT 2276.390 1007.570 2276.690 1019.495 ;
        RECT 2280.055 1016.775 2280.385 1017.105 ;
        RECT 2271.130 1004.550 2273.010 1004.850 ;
        RECT 2276.350 1007.270 2276.690 1007.570 ;
        RECT 2271.130 1001.635 2271.430 1004.550 ;
        RECT 2276.350 1001.635 2276.650 1007.270 ;
        RECT 2276.970 1004.850 2277.270 1006.235 ;
        RECT 2280.070 1004.850 2280.370 1016.775 ;
        RECT 2276.970 1004.550 2280.370 1004.850 ;
        RECT 2281.910 1006.235 2282.210 1020.855 ;
        RECT 2282.815 1020.175 2283.145 1020.505 ;
        RECT 2282.830 1006.235 2283.130 1020.175 ;
        RECT 2300.295 1016.775 2300.625 1017.105 ;
        RECT 2311.335 1016.775 2311.665 1017.105 ;
        RECT 2289.255 1016.095 2289.585 1016.425 ;
        RECT 2293.855 1016.095 2294.185 1016.425 ;
        RECT 2287.415 1014.735 2287.745 1015.065 ;
        RECT 2281.910 1004.550 2282.490 1006.235 ;
        RECT 2276.970 1001.635 2277.270 1004.550 ;
        RECT 2282.190 1001.635 2282.490 1004.550 ;
        RECT 2282.810 1004.550 2283.130 1006.235 ;
        RECT 2287.430 1004.850 2287.730 1014.735 ;
        RECT 2288.030 1004.850 2288.330 1006.235 ;
        RECT 2287.430 1004.550 2288.330 1004.850 ;
        RECT 2282.810 1001.635 2283.110 1004.550 ;
        RECT 2288.030 1001.635 2288.330 1004.550 ;
        RECT 2288.650 1004.850 2288.950 1006.235 ;
        RECT 2289.270 1004.850 2289.570 1016.095 ;
        RECT 2288.650 1004.550 2289.570 1004.850 ;
        RECT 2288.650 1001.635 2288.950 1004.550 ;
        RECT 2293.870 1001.635 2294.170 1016.095 ;
        RECT 2294.775 1014.735 2295.105 1015.065 ;
        RECT 2294.790 1006.235 2295.090 1014.735 ;
        RECT 2300.310 1008.250 2300.610 1016.775 ;
        RECT 2304.895 1016.095 2305.225 1016.425 ;
        RECT 2303.055 1014.735 2303.385 1015.065 ;
        RECT 2294.490 1004.550 2295.090 1006.235 ;
        RECT 2299.710 1007.950 2300.610 1008.250 ;
        RECT 2294.490 1001.635 2294.790 1004.550 ;
        RECT 2299.710 1001.635 2300.010 1007.950 ;
        RECT 2300.330 1004.850 2300.630 1006.235 ;
        RECT 2303.070 1004.850 2303.370 1014.735 ;
        RECT 2300.330 1004.550 2303.370 1004.850 ;
        RECT 2304.910 1004.850 2305.210 1016.095 ;
        RECT 2307.655 1014.735 2307.985 1015.065 ;
        RECT 2305.550 1004.850 2305.850 1006.235 ;
        RECT 2304.910 1004.550 2305.850 1004.850 ;
        RECT 2300.330 1001.635 2300.630 1004.550 ;
        RECT 2305.550 1001.635 2305.850 1004.550 ;
        RECT 2306.170 1004.850 2306.470 1006.235 ;
        RECT 2307.670 1004.850 2307.970 1014.735 ;
        RECT 2306.170 1004.550 2307.970 1004.850 ;
        RECT 2311.350 1006.235 2311.650 1016.775 ;
        RECT 2315.935 1016.095 2316.265 1016.425 ;
        RECT 2322.375 1016.095 2322.705 1016.425 ;
        RECT 2312.255 1014.735 2312.585 1015.065 ;
        RECT 2312.270 1006.235 2312.570 1014.735 ;
        RECT 2311.350 1004.550 2311.690 1006.235 ;
        RECT 2306.170 1001.635 2306.470 1004.550 ;
        RECT 2311.390 1001.635 2311.690 1004.550 ;
        RECT 2312.010 1004.550 2312.570 1006.235 ;
        RECT 2312.010 1001.635 2312.310 1004.550 ;
        RECT 2315.950 1004.085 2316.250 1016.095 ;
        RECT 2317.775 1014.735 2318.105 1015.065 ;
        RECT 2317.790 1008.250 2318.090 1014.735 ;
        RECT 2317.790 1007.950 2318.150 1008.250 ;
        RECT 2317.230 1004.085 2317.530 1006.235 ;
        RECT 2315.950 1003.785 2317.530 1004.085 ;
        RECT 2317.230 1001.635 2317.530 1003.785 ;
        RECT 2317.850 1001.635 2318.150 1007.950 ;
        RECT 2322.390 1004.850 2322.690 1016.095 ;
        RECT 2323.295 1014.735 2323.625 1015.065 ;
        RECT 2323.310 1008.250 2323.610 1014.735 ;
        RECT 2323.310 1007.950 2323.990 1008.250 ;
        RECT 2323.070 1004.850 2323.370 1006.235 ;
        RECT 2322.390 1004.550 2323.370 1004.850 ;
        RECT 2323.070 1001.635 2323.370 1004.550 ;
        RECT 2323.690 1001.635 2323.990 1007.950 ;
        RECT 2328.830 1006.235 2329.130 1020.855 ;
        RECT 2329.735 1014.735 2330.065 1015.065 ;
        RECT 2329.750 1006.235 2330.050 1014.735 ;
        RECT 2328.830 1004.550 2329.210 1006.235 ;
        RECT 2328.910 1001.635 2329.210 1004.550 ;
        RECT 2329.530 1004.550 2330.050 1006.235 ;
        RECT 2329.530 1001.635 2329.830 1004.550 ;
        RECT 2333.430 1004.085 2333.730 1020.855 ;
        RECT 2335.255 1014.735 2335.585 1015.065 ;
        RECT 2335.270 1007.570 2335.570 1014.735 ;
        RECT 2340.790 1007.570 2341.090 1020.855 ;
        RECT 2346.295 1020.175 2346.625 1020.505 ;
        RECT 2342.615 1014.735 2342.945 1015.065 ;
        RECT 2335.270 1007.270 2335.670 1007.570 ;
        RECT 2334.750 1004.085 2335.050 1006.235 ;
        RECT 2333.430 1003.785 2335.050 1004.085 ;
        RECT 2334.750 1001.635 2335.050 1003.785 ;
        RECT 2335.370 1001.635 2335.670 1007.270 ;
        RECT 2340.590 1007.270 2341.090 1007.570 ;
        RECT 2340.590 1001.635 2340.890 1007.270 ;
        RECT 2341.210 1004.085 2341.510 1006.235 ;
        RECT 2342.630 1004.085 2342.930 1014.735 ;
        RECT 2346.310 1006.235 2346.610 1020.175 ;
        RECT 2347.215 1014.735 2347.545 1015.065 ;
        RECT 2347.230 1006.235 2347.530 1014.735 ;
        RECT 2351.830 1007.570 2352.130 1020.855 ;
        RECT 2355.495 1014.735 2355.825 1015.065 ;
        RECT 2351.830 1007.270 2352.570 1007.570 ;
        RECT 2346.310 1004.550 2346.730 1006.235 ;
        RECT 2341.210 1003.785 2342.930 1004.085 ;
        RECT 2341.210 1001.635 2341.510 1003.785 ;
        RECT 2346.430 1001.635 2346.730 1004.550 ;
        RECT 2347.050 1004.550 2347.530 1006.235 ;
        RECT 2347.050 1001.635 2347.350 1004.550 ;
        RECT 2352.270 1001.635 2352.570 1007.270 ;
        RECT 2352.890 1004.850 2353.190 1006.235 ;
        RECT 2355.510 1004.850 2355.810 1014.735 ;
        RECT 2358.270 1007.570 2358.570 1020.855 ;
        RECT 2361.015 1020.175 2361.345 1020.505 ;
        RECT 2359.175 1016.095 2359.505 1016.425 ;
        RECT 2352.890 1004.550 2355.810 1004.850 ;
        RECT 2358.110 1007.270 2358.570 1007.570 ;
        RECT 2359.190 1007.570 2359.490 1016.095 ;
        RECT 2359.190 1007.270 2360.410 1007.570 ;
        RECT 2352.890 1001.635 2353.190 1004.550 ;
        RECT 2358.110 1001.635 2358.410 1007.270 ;
        RECT 2358.730 1004.085 2359.030 1006.235 ;
        RECT 2360.110 1004.085 2360.410 1007.270 ;
        RECT 2361.030 1004.850 2361.330 1020.175 ;
        RECT 2364.695 1014.735 2365.025 1015.065 ;
        RECT 2367.455 1014.735 2367.785 1015.065 ;
        RECT 2372.975 1014.735 2373.305 1015.065 ;
        RECT 2364.710 1006.235 2365.010 1014.735 ;
        RECT 2363.950 1004.850 2364.250 1006.235 ;
        RECT 2361.030 1004.550 2364.250 1004.850 ;
        RECT 2358.730 1003.785 2360.410 1004.085 ;
        RECT 2358.730 1001.635 2359.030 1003.785 ;
        RECT 2363.950 1001.635 2364.250 1004.550 ;
        RECT 2364.570 1004.550 2365.010 1006.235 ;
        RECT 2367.470 1004.850 2367.770 1014.735 ;
        RECT 2369.790 1004.850 2370.090 1006.235 ;
        RECT 2367.470 1004.550 2370.090 1004.850 ;
        RECT 2364.570 1001.635 2364.870 1004.550 ;
        RECT 2369.790 1001.635 2370.090 1004.550 ;
        RECT 2370.410 1004.850 2370.710 1006.235 ;
        RECT 2372.990 1004.850 2373.290 1014.735 ;
        RECT 2370.410 1004.550 2373.290 1004.850 ;
        RECT 2373.910 1004.850 2374.210 1020.855 ;
        RECT 2381.255 1020.175 2381.585 1020.505 ;
        RECT 2387.695 1020.175 2388.025 1020.505 ;
        RECT 2377.575 1014.735 2377.905 1015.065 ;
        RECT 2375.630 1004.850 2375.930 1006.235 ;
        RECT 2373.910 1004.550 2375.930 1004.850 ;
        RECT 2370.410 1001.635 2370.710 1004.550 ;
        RECT 2375.630 1001.635 2375.930 1004.550 ;
        RECT 2376.250 1004.085 2376.550 1006.235 ;
        RECT 2377.590 1004.085 2377.890 1014.735 ;
        RECT 2381.270 1006.235 2381.570 1020.175 ;
        RECT 2382.175 1014.735 2382.505 1015.065 ;
        RECT 2382.190 1006.235 2382.490 1014.735 ;
        RECT 2387.710 1007.570 2388.010 1020.175 ;
        RECT 2393.215 1016.775 2393.545 1017.105 ;
        RECT 2395.975 1016.775 2396.305 1017.105 ;
        RECT 2390.455 1016.095 2390.785 1016.425 ;
        RECT 2388.615 1014.735 2388.945 1015.065 ;
        RECT 2381.270 1004.550 2381.770 1006.235 ;
        RECT 2376.250 1003.785 2377.890 1004.085 ;
        RECT 2376.250 1001.635 2376.550 1003.785 ;
        RECT 2381.470 1001.635 2381.770 1004.550 ;
        RECT 2382.090 1004.550 2382.490 1006.235 ;
        RECT 2387.310 1007.270 2388.010 1007.570 ;
        RECT 2382.090 1001.635 2382.390 1004.550 ;
        RECT 2387.310 1001.635 2387.610 1007.270 ;
        RECT 2387.930 1004.850 2388.230 1006.235 ;
        RECT 2388.630 1004.850 2388.930 1014.735 ;
        RECT 2387.930 1004.550 2388.930 1004.850 ;
        RECT 2390.470 1004.850 2390.770 1016.095 ;
        RECT 2393.230 1007.570 2393.530 1016.775 ;
        RECT 2393.230 1007.270 2394.070 1007.570 ;
        RECT 2393.150 1004.850 2393.450 1006.235 ;
        RECT 2390.470 1004.550 2393.450 1004.850 ;
        RECT 2387.930 1001.635 2388.230 1004.550 ;
        RECT 2393.150 1001.635 2393.450 1004.550 ;
        RECT 2393.770 1001.635 2394.070 1007.270 ;
        RECT 2395.990 1004.850 2396.290 1016.775 ;
        RECT 2399.655 1014.735 2399.985 1015.065 ;
        RECT 2399.670 1006.235 2399.970 1014.735 ;
        RECT 2398.990 1004.850 2399.290 1006.235 ;
        RECT 2395.990 1004.550 2399.290 1004.850 ;
        RECT 2398.990 1001.635 2399.290 1004.550 ;
        RECT 2399.610 1004.550 2399.970 1006.235 ;
        RECT 2403.350 1004.850 2403.650 1020.855 ;
        RECT 2408.855 1018.135 2409.185 1018.465 ;
        RECT 2406.095 1014.735 2406.425 1015.065 ;
        RECT 2404.830 1004.850 2405.130 1006.235 ;
        RECT 2403.350 1004.550 2405.130 1004.850 ;
        RECT 2399.610 1001.635 2399.910 1004.550 ;
        RECT 2404.830 1001.635 2405.130 1004.550 ;
        RECT 2405.450 1004.850 2405.750 1006.235 ;
        RECT 2406.110 1004.850 2406.410 1014.735 ;
        RECT 2405.450 1004.550 2406.410 1004.850 ;
        RECT 2408.870 1004.850 2409.170 1018.135 ;
        RECT 2410.695 1017.455 2411.025 1017.785 ;
        RECT 2410.710 1008.250 2411.010 1017.455 ;
        RECT 2415.295 1016.775 2415.625 1017.105 ;
        RECT 2410.710 1007.950 2411.590 1008.250 ;
        RECT 2410.670 1004.850 2410.970 1006.235 ;
        RECT 2408.870 1004.550 2410.970 1004.850 ;
        RECT 2405.450 1001.635 2405.750 1004.550 ;
        RECT 2410.670 1001.635 2410.970 1004.550 ;
        RECT 2411.290 1001.635 2411.590 1007.950 ;
        RECT 2415.310 1004.850 2415.610 1016.775 ;
        RECT 2417.135 1014.735 2417.465 1015.065 ;
        RECT 2417.150 1006.235 2417.450 1014.735 ;
        RECT 2416.510 1004.850 2416.810 1006.235 ;
        RECT 2415.310 1004.550 2416.810 1004.850 ;
        RECT 2416.510 1001.635 2416.810 1004.550 ;
        RECT 2417.130 1004.550 2417.450 1006.235 ;
        RECT 2421.750 1004.850 2422.050 1020.855 ;
        RECT 2451.175 1020.175 2451.505 1020.505 ;
        RECT 2429.095 1018.815 2429.425 1019.145 ;
        RECT 2423.575 1016.775 2423.905 1017.105 ;
        RECT 2422.350 1004.850 2422.650 1006.235 ;
        RECT 2421.750 1004.550 2422.650 1004.850 ;
        RECT 2417.130 1001.635 2417.430 1004.550 ;
        RECT 2422.350 1001.635 2422.650 1004.550 ;
        RECT 2422.970 1004.850 2423.270 1006.235 ;
        RECT 2423.590 1004.850 2423.890 1016.775 ;
        RECT 2429.110 1006.235 2429.410 1018.815 ;
        RECT 2431.855 1018.135 2432.185 1018.465 ;
        RECT 2422.970 1004.550 2423.890 1004.850 ;
        RECT 2428.810 1004.550 2429.410 1006.235 ;
        RECT 2431.870 1004.850 2432.170 1018.135 ;
        RECT 2437.375 1017.455 2437.705 1017.785 ;
        RECT 2434.650 1004.850 2434.950 1006.235 ;
        RECT 2431.870 1004.550 2434.950 1004.850 ;
        RECT 2437.390 1004.850 2437.690 1017.455 ;
        RECT 2442.895 1016.095 2443.225 1016.425 ;
        RECT 2440.490 1004.850 2440.790 1006.235 ;
        RECT 2437.390 1004.550 2440.790 1004.850 ;
        RECT 2442.910 1004.850 2443.210 1016.095 ;
        RECT 2446.330 1004.850 2446.630 1006.235 ;
        RECT 2442.910 1004.550 2446.630 1004.850 ;
        RECT 2451.190 1004.850 2451.490 1020.175 ;
        RECT 2452.170 1004.850 2452.470 1006.235 ;
        RECT 2451.190 1004.550 2452.470 1004.850 ;
        RECT 2422.970 1001.635 2423.270 1004.550 ;
        RECT 2428.810 1001.635 2429.110 1004.550 ;
        RECT 2434.650 1001.635 2434.950 1004.550 ;
        RECT 2440.490 1001.635 2440.790 1004.550 ;
        RECT 2446.330 1001.635 2446.630 1004.550 ;
        RECT 2452.170 1001.635 2452.470 1004.550 ;
      LAYER met4 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met4 ;
        RECT 1598.715 550.000 1599.015 554.600 ;
        RECT 1604.955 550.000 1605.255 554.600 ;
        RECT 1611.195 550.000 1611.495 554.600 ;
        RECT 1617.435 550.000 1617.735 554.600 ;
        RECT 1623.675 550.000 1623.975 554.600 ;
        RECT 1629.915 550.000 1630.215 554.600 ;
        RECT 1636.155 550.000 1636.455 554.600 ;
        RECT 1642.395 550.000 1642.695 554.600 ;
        RECT 1648.635 550.000 1648.935 554.600 ;
        RECT 1654.875 550.000 1655.175 554.600 ;
        RECT 1661.115 550.000 1661.415 554.600 ;
        RECT 1667.355 550.000 1667.655 554.600 ;
        RECT 1673.595 550.000 1673.895 554.600 ;
        RECT 1679.835 550.000 1680.135 554.600 ;
        RECT 1686.075 550.000 1686.375 554.600 ;
        RECT 1692.315 550.000 1692.615 554.600 ;
        RECT 1698.555 550.000 1698.855 554.600 ;
        RECT 1704.795 550.000 1705.095 554.600 ;
        RECT 1711.035 550.000 1711.335 554.600 ;
        RECT 1717.275 550.000 1717.575 554.600 ;
        RECT 1723.515 550.000 1723.815 554.600 ;
        RECT 1729.755 550.000 1730.055 554.600 ;
        RECT 1735.995 550.000 1736.295 554.600 ;
        RECT 1742.235 550.000 1742.535 554.600 ;
        RECT 1748.475 550.000 1748.775 554.600 ;
        RECT 1754.715 550.000 1755.015 554.600 ;
        RECT 1760.955 550.000 1761.255 554.600 ;
        RECT 1767.195 550.000 1767.495 554.600 ;
        RECT 1773.435 550.000 1773.735 554.600 ;
        RECT 1779.675 550.000 1779.975 554.600 ;
        RECT 1785.915 550.000 1786.215 554.600 ;
        RECT 1792.155 550.000 1792.455 554.600 ;
        RECT 2198.715 550.000 2199.015 554.600 ;
        RECT 2204.955 550.000 2205.255 554.600 ;
        RECT 2211.195 550.000 2211.495 554.600 ;
        RECT 2217.435 550.000 2217.735 554.600 ;
        RECT 2223.675 550.000 2223.975 554.600 ;
        RECT 2229.915 550.000 2230.215 554.600 ;
        RECT 2236.155 550.000 2236.455 554.600 ;
        RECT 2242.395 550.000 2242.695 554.600 ;
        RECT 2248.635 550.000 2248.935 554.600 ;
        RECT 2254.875 550.000 2255.175 554.600 ;
        RECT 2261.115 550.000 2261.415 554.600 ;
        RECT 2267.355 550.000 2267.655 554.600 ;
        RECT 2273.595 550.000 2273.895 554.600 ;
        RECT 2279.835 550.000 2280.135 554.600 ;
        RECT 2286.075 550.000 2286.375 554.600 ;
        RECT 2292.315 550.000 2292.615 554.600 ;
        RECT 2298.555 550.000 2298.855 554.600 ;
        RECT 2304.795 550.000 2305.095 554.600 ;
        RECT 2311.035 550.000 2311.335 554.600 ;
        RECT 2317.275 550.000 2317.575 554.600 ;
        RECT 2323.515 550.000 2323.815 554.600 ;
        RECT 2329.755 550.000 2330.055 554.600 ;
        RECT 2335.995 550.000 2336.295 554.600 ;
        RECT 2342.235 550.000 2342.535 554.600 ;
        RECT 2348.475 550.000 2348.775 554.600 ;
        RECT 2354.715 550.000 2355.015 554.600 ;
        RECT 2360.955 550.000 2361.255 554.600 ;
        RECT 2367.195 550.000 2367.495 554.600 ;
        RECT 2373.435 550.000 2373.735 554.600 ;
        RECT 2379.675 550.000 2379.975 554.600 ;
        RECT 2385.915 550.000 2386.215 554.600 ;
        RECT 2392.155 550.000 2392.455 554.600 ;
  END
END user_project_wrapper
END LIBRARY

